* NGSPICE file created from core0.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_12 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

.subckt core0 dbg_pc[0] dbg_pc[10] dbg_pc[11] dbg_pc[12] dbg_pc[13] dbg_pc[14] dbg_pc[15]
+ dbg_pc[1] dbg_pc[2] dbg_pc[3] dbg_pc[4] dbg_pc[5] dbg_pc[6] dbg_pc[7] dbg_pc[8]
+ dbg_pc[9] dbg_r0[0] dbg_r0[10] dbg_r0[11] dbg_r0[12] dbg_r0[13] dbg_r0[14] dbg_r0[15]
+ dbg_r0[1] dbg_r0[2] dbg_r0[3] dbg_r0[4] dbg_r0[5] dbg_r0[6] dbg_r0[7] dbg_r0[8]
+ dbg_r0[9] i_clk i_core_int_sreg[0] i_core_int_sreg[10] i_core_int_sreg[11] i_core_int_sreg[12]
+ i_core_int_sreg[13] i_core_int_sreg[14] i_core_int_sreg[15] i_core_int_sreg[1] i_core_int_sreg[2]
+ i_core_int_sreg[3] i_core_int_sreg[4] i_core_int_sreg[5] i_core_int_sreg[6] i_core_int_sreg[7]
+ i_core_int_sreg[8] i_core_int_sreg[9] i_disable i_irq i_mc_core_int i_mem_ack i_mem_data[0]
+ i_mem_data[10] i_mem_data[11] i_mem_data[12] i_mem_data[13] i_mem_data[14] i_mem_data[15]
+ i_mem_data[1] i_mem_data[2] i_mem_data[3] i_mem_data[4] i_mem_data[5] i_mem_data[6]
+ i_mem_data[7] i_mem_data[8] i_mem_data[9] i_mem_exception i_req_data[0] i_req_data[10]
+ i_req_data[11] i_req_data[12] i_req_data[13] i_req_data[14] i_req_data[15] i_req_data[16]
+ i_req_data[17] i_req_data[18] i_req_data[19] i_req_data[1] i_req_data[20] i_req_data[21]
+ i_req_data[22] i_req_data[23] i_req_data[24] i_req_data[25] i_req_data[26] i_req_data[27]
+ i_req_data[28] i_req_data[29] i_req_data[2] i_req_data[30] i_req_data[31] i_req_data[3]
+ i_req_data[4] i_req_data[5] i_req_data[6] i_req_data[7] i_req_data[8] i_req_data[9]
+ i_req_data_valid i_rst o_c_data_page o_c_instr_long o_c_instr_page o_icache_flush
+ o_instr_long_addr[0] o_instr_long_addr[1] o_instr_long_addr[2] o_instr_long_addr[3]
+ o_instr_long_addr[4] o_instr_long_addr[5] o_instr_long_addr[6] o_instr_long_addr[7]
+ o_mem_addr[0] o_mem_addr[10] o_mem_addr[11] o_mem_addr[12] o_mem_addr[13] o_mem_addr[14]
+ o_mem_addr[15] o_mem_addr[1] o_mem_addr[2] o_mem_addr[3] o_mem_addr[4] o_mem_addr[5]
+ o_mem_addr[6] o_mem_addr[7] o_mem_addr[8] o_mem_addr[9] o_mem_addr_high[0] o_mem_addr_high[1]
+ o_mem_addr_high[2] o_mem_addr_high[3] o_mem_addr_high[4] o_mem_addr_high[5] o_mem_addr_high[6]
+ o_mem_data[0] o_mem_data[10] o_mem_data[11] o_mem_data[12] o_mem_data[13] o_mem_data[14]
+ o_mem_data[15] o_mem_data[1] o_mem_data[2] o_mem_data[3] o_mem_data[4] o_mem_data[5]
+ o_mem_data[6] o_mem_data[7] o_mem_data[8] o_mem_data[9] o_mem_long o_mem_req o_mem_sel[0]
+ o_mem_sel[1] o_mem_we o_req_active o_req_addr[0] o_req_addr[10] o_req_addr[11] o_req_addr[12]
+ o_req_addr[13] o_req_addr[14] o_req_addr[15] o_req_addr[1] o_req_addr[2] o_req_addr[3]
+ o_req_addr[4] o_req_addr[5] o_req_addr[6] o_req_addr[7] o_req_addr[8] o_req_addr[9]
+ o_req_ppl_submit sr_bus_addr[0] sr_bus_addr[10] sr_bus_addr[11] sr_bus_addr[12]
+ sr_bus_addr[13] sr_bus_addr[14] sr_bus_addr[15] sr_bus_addr[1] sr_bus_addr[2] sr_bus_addr[3]
+ sr_bus_addr[4] sr_bus_addr[5] sr_bus_addr[6] sr_bus_addr[7] sr_bus_addr[8] sr_bus_addr[9]
+ sr_bus_data_o[0] sr_bus_data_o[10] sr_bus_data_o[11] sr_bus_data_o[12] sr_bus_data_o[13]
+ sr_bus_data_o[14] sr_bus_data_o[15] sr_bus_data_o[1] sr_bus_data_o[2] sr_bus_data_o[3]
+ sr_bus_data_o[4] sr_bus_data_o[5] sr_bus_data_o[6] sr_bus_data_o[7] sr_bus_data_o[8]
+ sr_bus_data_o[9] sr_bus_we vccd1 vssd1 o_mem_addr_high[7]
XFILLER_0_185_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__A2 _1833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7963_ core_0.execute.rf.reg_outputs\[5\]\[5\] _3679_ _3677_ _3681_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5968__A1 _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8126__B _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6914_ _2510_ _2845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7894_ _3451_ _3628_ _3640_ _0387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7709__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_2418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7965__B _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ _1405_ net227 _2683_ _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_9633_ _0643_ clknet_leaf_96_i_clk net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_175_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9564_ _0574_ clknet_leaf_81_i_clk core_0.execute.sreg_irq_pc.o_d\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_190_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6776_ _2708_ _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6393__A1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8515_ net85 _4040_ _4101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5727_ _1714_ _1722_ _0138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4943__A2 _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9495_ _0505_ clknet_leaf_18_i_clk net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_134_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8134__A2 _3758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8446_ _2136_ _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_72_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ _1628_ _1665_ _1666_ _0125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8796__B _4324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_211_3040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7893__A1 core_0.execute.rf.reg_outputs\[7\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4609_ _0794_ _0799_ _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_170_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8377_ _3802_ _3989_ _3990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5589_ _1465_ core_0.fetch.submitable _1625_ _0097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7328_ _1338_ _1988_ _1285_ _3249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_102_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_217_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6448__A2 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7645__A1 core_0.ew_reg_ie\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_2703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7259_ _2564_ _2844_ _3181_ _3182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_217_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_183_2714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7948__A2 _3394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5959__A1 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_222_3180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8036__B _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4631__A1 core_0.execute.rf.reg_outputs\[12\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4631__B2 core_0.execute.rf.reg_outputs\[13\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7875__B _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_103_1749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8373__A2 _3886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_194_2843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5187__A2 _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4934__A2 _1060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8125__A2 _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xrebuffer7 _1831_ net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_106_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6687__A2 net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7884__A1 core_0.execute.rf.reg_outputs\[7\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4698__A1 core_0.execute.rf.reg_outputs\[5\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8428__A3 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7636__A1 _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7487__I1 core_0.ew_reg_ie\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_225_3209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_120_i_clk clknet_4_7__leaf_i_clk clknet_leaf_120_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5111__A2 core_0.decode.i_instr_l\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4870__A1 _1016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7939__A2 _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8061__A1 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_135_i_clk clknet_4_3__leaf_i_clk clknet_leaf_135_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4960_ _1070_ _1139_ _1140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_35_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_148_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4891_ net59 core_0.fetch.out_buffer_data_instr\[2\] _0894_ _1072_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_175_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_236_3349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6630_ _2070_ _2041_ _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5178__A2 _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6561_ _1869_ _1873_ _1877_ _1811_ _2503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__8116__A2 _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8300_ _3914_ _1812_ _3917_ _1536_ _3918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_144_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5512_ net53 _1556_ _1583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_154_2359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9280_ _0290_ clknet_leaf_32_i_clk core_0.execute.rf.reg_outputs\[13\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6127__A1 _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7009__C _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9305__CLK clknet_leaf_3_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6492_ _1749_ net218 _2434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_125_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8231_ _2090_ _2102_ _2115_ _1812_ core_0.execute.alu_mul_div.cbit\[0\] core_0.execute.alu_mul_div.cbit\[1\]
+ _3854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_125_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6678__A2 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ core_0.execute.alu_mul_div.cbit\[2\] _1538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7875__A1 core_0.execute.rf.reg_outputs\[7\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4689__A1 core_0.execute.rf.reg_outputs\[7\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6848__C core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4689__B2 core_0.execute.rf.reg_outputs\[13\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8162_ _3456_ _3781_ _3794_ _0501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_196_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5374_ _1464_ _1483_ _0023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5350__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7113_ core_0.execute.alu_mul_div.div_cur\[7\] _1317_ _3037_ _3039_ _3040_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_8093_ _3465_ _3738_ _3754_ _0472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_238_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _1326_ _2970_ _2971_ _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_129_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5102__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6864__B _2795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6356__S _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5653__A3 net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_2488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8052__A1 _3459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8995_ _0022_ clknet_leaf_140_i_clk core_0.dec_rf_ie\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7946_ core_0.execute.rf.reg_outputs\[6\]\[15\] _3650_ _3663_ _3670_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4613__A1 core_0.execute.rf.reg_outputs\[5\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5810__B1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7877_ core_0.execute.rf.reg_outputs\[7\]\[1\] _3629_ _3621_ _3631_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8355__A2 _3915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9616_ _0626_ clknet_leaf_109_i_clk core_0.dec_sreg_irt vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_42_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6828_ _2745_ _2754_ _2760_ _2761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5169__A2 _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4916__A2 _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9547_ _0557_ clknet_leaf_134_i_clk core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6759_ _1690_ net177 _1405_ _1421_ _2693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_162_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8107__A2 _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9478_ _0488_ clknet_leaf_145_i_clk core_0.execute.rf.reg_outputs\[1\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6669__A2 _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7866__A1 core_0.execute.rf.reg_outputs\[8\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8429_ _4013_ _4029_ core_0.execute.alu_mul_div.div_res\[8\] _4030_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7618__A1 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5234__I _1362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8291__A1 _3901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5644__A3 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6841__A2 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_52_i_clk clknet_4_10__leaf_i_clk clknet_leaf_52_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8043__A1 _3446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4604__A1 core_0.execute.rf.reg_outputs\[1\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_67_i_clk clknet_4_12__leaf_i_clk clknet_leaf_67_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Left_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_200_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4907__A2 _1023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7306__B1 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5580__A2 _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_231_3279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9478__CLK clknet_leaf_145_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5332__A2 _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__B1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_74_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8282__A1 _3893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5090_ _1246_ _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5096__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8034__A1 _3420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6045__B1 _1801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7800_ core_0.execute.rf.reg_outputs\[9\]\[0\] _3586_ _3580_ _3587_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8780_ _0713_ _4295_ _4314_ _4307_ _0599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_188_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5992_ core_0.execute.rf.reg_outputs\[5\]\[13\] _1785_ _1802_ core_0.execute.rf.reg_outputs\[14\]\[13\]
+ _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7731_ core_0.execute.rf.reg_outputs\[11\]\[3\] _3543_ _3539_ _3547_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4943_ core_0.fetch.prev_request_pc\[8\] _1046_ _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8337__A2 _2366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6703__I _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7662_ core_0.execute.rf.reg_outputs\[13\]\[6\] _3504_ _3500_ _3507_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4874_ core_0.fetch.out_buffer_data_instr\[27\] _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9401_ _0411_ clknet_leaf_25_i_clk core_0.execute.rf.reg_outputs\[5\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6613_ _2423_ _2482_ _2554_ _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7593_ core_0.execute.rf.reg_outputs\[15\]\[12\] _3429_ _3422_ _3464_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5020__A1 net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9332_ _0342_ clknet_leaf_6_i_clk core_0.execute.rf.reg_outputs\[10\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6544_ _2060_ _2061_ _2062_ _2067_ _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_104_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9263_ _0273_ clknet_leaf_33_i_clk core_0.execute.rf.reg_outputs\[14\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7848__A1 _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6475_ _0891_ _1420_ _2418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__7534__I _3414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8214_ _3838_ _3839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5426_ _1321_ _1322_ _1340_ _1507_ _1523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_9194_ _0205_ clknet_leaf_54_i_clk core_0.ew_data\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5323__A2 core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6520__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_2517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8145_ _0891_ _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5357_ _1471_ _1437_ _1461_ _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XPHY_EDGE_ROW_206_Left_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_239_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8076_ core_0.execute.rf.reg_outputs\[2\]\[5\] _3743_ _3745_ _3746_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5288_ net188 net187 net190 net189 _1409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA_input36_I i_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5087__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7027_ core_0.execute.sreg_irq_pc.o_d\[5\] _2774_ _2775_ core_0.execute.pc_high_out\[5\]
+ _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_226_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__A1 _1011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8978_ core_0.dec_rf_ie\[0\] _1482_ _1470_ _1462_ _4457_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_242_17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7929_ core_0.execute.rf.reg_outputs\[6\]\[7\] _3657_ _3648_ _3661_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_178_2646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_215_Left_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_210_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6339__A1 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_191_2802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7000__A2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5011__A1 core_0.fetch.prev_request_pc\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9620__CLK clknet_leaf_133_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_137_Right_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5562__A2 _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6511__A1 _1745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_224_Left_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_189_2775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_2786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9000__CLK clknet_leaf_133_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__A2 _2115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8016__A1 _3462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_2956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_233_Left_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4589__B1 _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7619__I _3475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_233_3308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5139__I core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_104_Right_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5553__A2 _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _0778_ _0779_ _0780_ _0781_ _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_142_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6750__A1 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_2329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__I _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5583__B _1622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6260_ _2215_ _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6502__A1 _2008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5305__A2 _1418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5211_ core_0.ew_data\[1\] net156 _1351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4513__B1 _0710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6191_ core_0.execute.alu_mul_div.div_cur\[3\] _2075_ _2180_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_244_3437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5142_ _1232_ _1241_ _1280_ _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_209_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_236_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6805__A2 _2492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5073_ _0891_ _1229_ _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_208_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8901_ _1231_ _1528_ _4412_ _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7022__C _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_2458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_239_Right_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_8832_ core_0.execute.pc_high_buff_out\[4\] _4335_ _4357_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7230__A2 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5975_ _1963_ _1964_ _1965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8763_ core_0.execute.sreg_scratch.o_d\[8\] _4300_ _4305_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8134__B _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ core_0.fetch.prev_request_pc\[6\] _1106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7714_ _3463_ _3521_ _3536_ _0311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8694_ net72 _1740_ _1721_ _4256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_192_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5792__A2 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clone29_I _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7973__B _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4857_ net51 core_0.fetch.out_buffer_data_instr\[22\] _0893_ _1038_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7645_ core_0.ew_reg_ie\[13\] _3395_ _3496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_7_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8730__A2 _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7576_ _3450_ _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_15_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5544__A2 _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4788_ _0962_ _0968_ _0969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6527_ net240 _1988_ _2469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9315_ _0325_ clknet_leaf_10_i_clk core_0.execute.rf.reg_outputs\[11\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9246_ _0256_ clknet_leaf_37_i_clk core_0.execute.rf.reg_outputs\[15\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6458_ _2411_ _2386_ _2412_ _0179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5409_ _0958_ _1486_ _1511_ _1501_ _0030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_9177_ _0188_ clknet_leaf_41_i_clk core_0.execute.sreg_irq_flags.i_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6389_ _1544_ _2362_ _2363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_208_3012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8128_ core_0.execute.rf.reg_outputs\[1\]\[12\] _3765_ _3771_ _3775_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_50_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8059_ core_0.execute.rf.reg_outputs\[3\]\[15\] _3714_ _3730_ _3735_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4807__A1 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9173__CLK clknet_leaf_42_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_126_2022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_82_Left_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_230_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_206_Right_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7221__A2 _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8044__B _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_22_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_219_3141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6980__A1 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5783__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8721__A2 _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6732__A1 core_0.execute.rf.reg_outputs\[1\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_91_Left_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6732__B2 core_0.execute.rf.reg_outputs\[3\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8485__A1 _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6011__C _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5299__A1 _0995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8237__A1 _2349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5422__I _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_148_2291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_233_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8733__I _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__A1 core_0.ew_data\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _1519_ net185 _1750_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8889__B _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_174_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5774__A2 _1760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4711_ _0892_ _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_29_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7793__B _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5691_ _1420_ _1695_ _1696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_29_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7430_ _2130_ _2419_ _3348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4642_ _0826_ _0827_ _0828_ _0829_ _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_154_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5526__A2 _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6723__A1 core_0.execute.rf.reg_outputs\[7\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6723__B2 core_0.execute.rf.reg_outputs\[5\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4734__B1 _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7361_ _2554_ _3280_ _1326_ _3281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4573_ core_0.execute.rf.reg_outputs\[10\]\[10\] net221 net220 core_0.execute.rf.reg_outputs\[9\]\[10\]
+ _0766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_130_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6312_ _2291_ _2292_ _0153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9100_ _0125_ clknet_leaf_97_i_clk core_0.decode.i_jmp_pred_pass vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8476__A1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8476__B2 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7292_ _1338_ _3212_ _2471_ _1885_ _3213_ _3214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_9031_ _0058_ clknet_leaf_88_i_clk core_0.fetch.out_buffer_data_instr\[19\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6243_ core_0.execute.alu_mul_div.div_cur\[1\] _1930_ _2231_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8228__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6174_ _2161_ _2162_ _2163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_139_Left_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5125_ core_0.decode.i_instr_l\[3\] core_0.decode.i_instr_l\[2\] _1280_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_209_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7451__A2 _3155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ core_0.fetch.prev_request_pc\[1\] core_0.fetch.prev_request_pc\[0\] _1222_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_137_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_224_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5462__A1 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__A2 _3126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8815_ core_0.execute.pc_high_out\[2\] core_0.execute.pc_high_out\[1\] core_0.execute.pc_high_out\[0\]
+ _4342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_39_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8400__A1 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_220_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8951__A2 _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_148_Left_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8746_ core_0.execute.sreg_scratch.o_d\[0\] _4295_ _4296_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_2616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5958_ core_0.execute.rf.reg_outputs\[6\]\[11\] _1799_ _1819_ core_0.execute.rf.reg_outputs\[12\]\[11\]
+ _1788_ core_0.execute.rf.reg_outputs\[3\]\[11\] _1948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5765__A2 net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4909_ core_0.fetch.prev_request_pc\[13\] _1026_ _1089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8677_ net84 _1699_ _1715_ _4205_ _4242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5889_ _1292_ _1326_ _1876_ _1877_ _1879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_35_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8703__A2 _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7506__A3 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5517__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7628_ _3447_ _3476_ _3487_ _0274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6714__A1 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_214_3082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7559_ _3397_ _3435_ _3436_ _0256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6190__A2 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_160_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9229_ _0240_ clknet_leaf_142_i_clk core_0.ew_reg_ie\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_132_2092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_2745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8219__A1 _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7690__A2 _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7442__A2 _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5453__A1 _1001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_201_2926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8942__A2 _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_197_2874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6953__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6705__A1 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__A2 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_5 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7130__A1 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7681__A2 _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5692__A1 _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7788__B _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7433__A2 _2766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer17 net208 net245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_179_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer28 net254 net256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6930_ _2076_ _2733_ _2860_ _1898_ _2861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_178_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer39 net319 net320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5995__A2 _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7300__C _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7197__A1 core_0.execute.sreg_priv_control.o_d\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6861_ _1896_ _2505_ _2506_ _2793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7197__B2 net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8600_ core_0.execute.alu_flag_reg.o_d\[2\] _4167_ _3797_ _4176_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5812_ _1801_ _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_201_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6792_ _1898_ _2723_ _2724_ _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_9580_ _0590_ clknet_leaf_21_i_clk core_0.execute.sreg_scratch.o_d\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5747__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6944__A1 core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6944__B2 core_0.execute.sreg_scratch.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8531_ _4039_ _4114_ _4115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5743_ _1714_ _1733_ _0143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8462_ net79 _4053_ _4054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5674_ _1538_ _1670_ _1680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_199_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4970__A3 _1149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7413_ _1743_ _3330_ _3331_ _0996_ _3332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4625_ core_0.execute.rf.reg_outputs\[10\]\[6\] net221 net220 core_0.execute.rf.reg_outputs\[9\]\[6\]
+ _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_154_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8393_ _2140_ _3954_ _4003_ _4004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6172__A2 _1835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_2557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7344_ core_0.execute.sreg_irq_pc.o_d\[13\] _3042_ _3044_ core_0.execute.sreg_scratch.o_d\[13\]
+ _3265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4556_ core_0.execute.rf.reg_outputs\[6\]\[12\] _0670_ _0710_ core_0.execute.rf.reg_outputs\[8\]\[12\]
+ _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_96_1662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7275_ _1684_ _3196_ _3197_ _3198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7121__A1 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7542__I _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4487_ _0668_ net300 net292 _0685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_9014_ _0041_ clknet_leaf_102_i_clk core_0.fetch.out_buffer_data_instr\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6226_ _2206_ _2214_ _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_0_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_216_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__A2 _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ _2145_ _1852_ _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XTAP_TAPCELL_ROW_5_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _1263_ _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__8621__A1 net243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6088_ core_0.execute.rf.reg_outputs\[9\]\[3\] net224 _2078_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_240_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5039_ _1158_ _1149_ _1208_ _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_181_2686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5986__A2 _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_156_Left_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output105_I net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6935__A1 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__A2 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_216_3100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8729_ _1396_ _4283_ _4284_ _1431_ _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_192_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8688__A1 _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6699__B1 _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6163__A2 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_165_Left_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5910__A2 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7112__A1 _3038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7663__A2 _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput75 net75 dbg_pc[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_227_3240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput86 net86 dbg_pc[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput97 net97 dbg_r0[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8612__A1 _3079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7415__A2 _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_199_2903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_174_Left_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5700__I _1417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5977__A2 _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7179__A1 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8915__A2 _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6926__A1 _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5729__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5856__B _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8679__A1 _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_1938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_183_Left_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_30_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_156_2390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5390_ _1249_ _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_124_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5591__B _1626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8458__I _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7103__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_144_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7060_ _2587_ net272 _2987_ _2759_ _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__8851__A1 net288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7654__A2 _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_226_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6011_ _1874_ _1988_ _2000_ _1897_ _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5665__A1 _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4468__A2 _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8603__A1 _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5417__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7962_ _3427_ _3672_ _3680_ _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_178_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6090__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6913_ _2843_ _2586_ _2844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7893_ core_0.execute.rf.reg_outputs\[7\]\[8\] _3634_ _3636_ _3640_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__A2 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_2419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9632_ _0642_ clknet_leaf_101_i_clk net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6844_ _1405_ _1689_ _1691_ _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_92_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4928__B1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_69_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9563_ _0573_ clknet_leaf_71_i_clk core_0.execute.sreg_irq_pc.o_d\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6775_ core_0.dec_mem_access _2708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__6393__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7590__A1 _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_147_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8514_ _2401_ _4099_ _4100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5726_ core_0.execute.sreg_priv_control.o_d\[10\] _1701_ _1721_ _1698_ _1722_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9494_ _0504_ clknet_leaf_18_i_clk net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_162_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8445_ _2230_ _4038_ _0540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7342__A1 _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5657_ core_0.decode.i_jmp_pred_pass _1368_ _1666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7473__S _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_211_3041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4608_ _0795_ _0796_ _0797_ _0798_ _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__5353__B1 _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7893__A2 _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8376_ _3979_ _3974_ _3987_ _3989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_4_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5588_ _1137_ _1369_ _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_input66_I i_req_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4539_ _0731_ _0732_ _0733_ _0734_ _0735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7327_ net240 _2371_ _3248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__8842__A1 _4324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7645__A2 _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7258_ _2568_ _3179_ _3180_ _2563_ _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_183_2704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__A1 _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6209_ core_0.execute.alu_mul_div.div_cur\[10\] _1833_ _2198_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7189_ _2524_ _3112_ _3113_ _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_245_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5408__A1 core_0.decode.i_instr_l\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7221__B _3073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5408__B2 core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8070__A2 _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_222_3181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4631__A2 _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4919__B1 _1026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_194_2844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5395__C _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7891__B _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer8 net235 net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7884__A2 _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4698__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8428__A4 _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8833__A1 _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7636__A2 _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5647__A1 _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_208_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9257__CLK clknet_leaf_3_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4755__B _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8061__A2 _3394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A1 core_0.execute.rf.reg_outputs\[10\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_204_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4890_ net63 core_0.fetch.out_buffer_data_instr\[4\] _0893_ _1071_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_70_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_236_3339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7572__A1 core_0.execute.rf.reg_outputs\[15\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6375__A2 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6560_ _2501_ _2493_ _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_82_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5511_ _1027_ _1552_ _1582_ _0062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6491_ _1745_ _2039_ _2433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_202_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7324__A1 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8230_ _3847_ _3851_ _3852_ _3853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5442_ _1536_ _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7875__A2 _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4689__A2 net296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5886__A1 _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5373_ core_0.dec_rf_ie\[13\] _1482_ _1441_ _1472_ _1483_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8161_ net88 _3787_ _3785_ _3794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7112_ _3038_ _1314_ _2128_ _3039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8824__A1 core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8092_ core_0.execute.rf.reg_outputs\[2\]\[13\] _3743_ _3745_ _3754_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7627__A2 _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5638__A1 core_0.decode.i_imm_pass\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7043_ _2491_ _2499_ _2969_ _2971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_38_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5653__A4 core_0.ew_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_2489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6436__I net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8052__A2 _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8994_ _0021_ clknet_leaf_141_i_clk core_0.dec_rf_ie\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_210_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7945_ _3470_ _3652_ _3669_ _0409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_210_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_118_Right_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4613__A2 net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7876_ _3402_ _3628_ _3630_ _0379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9615_ _0625_ clknet_leaf_132_i_clk core_0.dec_sys vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_148_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6827_ _2341_ _2755_ _2758_ _2759_ _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5169__A3 _1289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9546_ _0556_ clknet_leaf_131_i_clk core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6758_ net186 _1688_ _1423_ _1424_ _2692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_190_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5709_ _1608_ _1710_ _0132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9477_ _0487_ clknet_leaf_145_i_clk core_0.execute.rf.reg_outputs\[1\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6118__A2 _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6689_ core_0.execute.rf.reg_outputs\[1\]\[2\] _2608_ _2609_ core_0.execute.rf.reg_outputs\[3\]\[2\]
+ _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_72_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8600__B _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8428_ _1537_ _2140_ _2354_ _3878_ _4029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_103_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7866__A2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5877__A1 _1768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output172_I net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8359_ core_0.execute.alu_mul_div.mul_res\[12\] _3972_ _3973_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_103_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7618__A2 _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5629__A1 _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_245_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_129_2064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8043__A2 _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6054__A1 core_0.execute.rf.reg_outputs\[8\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4604__A2 net308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5801__A1 _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7306__A1 core_0.execute.sreg_priv_control.o_d\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6109__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6949__C _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7857__A2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4540__A1 core_0.execute.rf.reg_outputs\[14\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__B2 core_0.execute.rf.reg_outputs\[12\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_102_Left_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8736__I _4288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6293__A1 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8034__A2 _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__A1 core_0.execute.rf.reg_outputs\[5\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5991_ core_0.execute.rf.reg_outputs\[1\]\[13\] _1779_ _1804_ core_0.execute.rf.reg_outputs\[11\]\[13\]
+ _1981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7793__A1 core_0.execute.rf.reg_outputs\[10\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7730_ _3415_ _3542_ _3546_ _0317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4942_ _1121_ _1096_ _1122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_111_Left_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7661_ _3435_ _3497_ _3506_ _0288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7545__A1 net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4873_ _1017_ net44 _1053_ _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_7_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9400_ _0410_ clknet_leaf_145_i_clk core_0.execute.rf.reg_outputs\[6\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6612_ _2550_ _2553_ _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7592_ _3462_ _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_55_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5020__A2 _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9331_ _0341_ clknet_leaf_8_i_clk core_0.execute.rf.reg_outputs\[10\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_171_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6543_ _1772_ _2056_ _2057_ _2058_ _2485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7815__I _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9262_ _0272_ clknet_leaf_26_i_clk core_0.execute.rf.reg_outputs\[14\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7848__A2 _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6474_ _2417_ _0189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5859__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8213_ _1679_ core_0.execute.alu_mul_div.mul_res\[1\] _3837_ _3838_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_42_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Right_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5425_ _1492_ _1520_ _1521_ _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_140_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9193_ _0204_ clknet_leaf_55_i_clk core_0.ew_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_113_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5323__A3 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6520__A2 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_120_Left_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5356_ core_0.decode.i_instr_l\[10\] _1471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8144_ _3414_ _3780_ _3784_ _0493_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_167_2518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9572__CLK clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6875__B _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8075_ _3647_ _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5287_ net186 net191 _1406_ _1407_ _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__7550__I _3396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5087__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7026_ core_0.execute.sreg_priv_control.o_d\[5\] _1692_ _2780_ net12 _2955_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_214_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input29_I i_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6166__I _1833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5070__I _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7233__B1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5003__C _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8576__A3 _3220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_195_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8977_ _1734_ _1438_ _1530_ _4307_ _0654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_195_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7928_ _3441_ _3651_ _3660_ _0401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_2647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6115__B _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7536__A1 _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7859_ core_0.execute.rf.reg_outputs\[8\]\[10\] _3613_ _3609_ _3620_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_100_1709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_191_2803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5547__B1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9529_ _0539_ clknet_leaf_120_i_clk core_0.execute.alu_mul_div.div_res\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_162_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output97_I net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_134_i_clk clknet_4_6__leaf_i_clk clknet_leaf_134_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6511__A2 _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4522__A1 net293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_2776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6277__S _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_149_i_clk clknet_4_0__leaf_i_clk clknet_leaf_149_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4825__A2 _0995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8016__A2 _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6027__A1 core_0.execute.rf.reg_outputs\[1\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_204_2957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7775__A1 _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4589__A1 core_0.execute.rf.reg_outputs\[7\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4589__B2 core_0.execute.rf.reg_outputs\[3\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9445__CLK clknet_leaf_145_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_122_1978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_233_3309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5002__A2 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6750__A2 _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_2319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6502__A2 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5210_ _1350_ net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4513__B2 core_0.execute.rf.reg_outputs\[8\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6190_ core_0.execute.alu_mul_div.div_cur\[4\] _1749_ _2179_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5141_ _1260_ _1261_ _1294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_244_3438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6266__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5072_ _1007_ _1228_ _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_224_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8900_ _4224_ _1286_ _4412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8007__A2 _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_162_2459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6018__A1 net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8831_ core_0.execute.pc_high_out\[4\] _4349_ _4356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_88_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8762_ _0813_ _4294_ _4304_ _4287_ _0591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_177_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5974_ core_0.execute.rf.reg_outputs\[13\]\[14\] _1792_ _1815_ core_0.execute.rf.reg_outputs\[9\]\[14\]
+ _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_177_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7713_ core_0.execute.rf.reg_outputs\[12\]\[12\] _3526_ _3528_ _3536_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4925_ core_0.fetch.prev_request_pc\[5\] _1105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_192_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8693_ _4219_ _4114_ _4255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7644_ _3473_ _3477_ _3495_ _0282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_157_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4856_ _0893_ net55 _1036_ _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_16_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8191__A1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7575_ _3387_ core_0.ew_data\[8\] _3449_ net35 _3450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4787_ _0965_ _0967_ _0968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_173_2588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9314_ _0324_ clknet_leaf_27_i_clk core_0.execute.rf.reg_outputs\[11\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_51_i_clk clknet_4_11__leaf_i_clk clknet_leaf_51_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6526_ _2424_ _2426_ _2467_ _2468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_42_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4752__A1 core_0.ew_reg_ie\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9245_ _0255_ clknet_leaf_33_i_clk core_0.execute.rf.reg_outputs\[15\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5065__I _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6457_ core_0.execute.mem_stage_pc\[15\] _1433_ _2404_ _2412_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7481__S _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ core_0.decode.i_instr_l\[11\] _1509_ _1510_ core_0.decode.i_instr_l\[7\] _1495_
+ _1511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_9176_ _0187_ clknet_leaf_42_i_clk core_0.execute.prev_pc_high\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6388_ _1542_ _1925_ _2361_ _2362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_208_3013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8127_ _3459_ _3760_ _3774_ _0486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_66_i_clk clknet_4_12__leaf_i_clk clknet_leaf_66_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_227_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5339_ _1257_ _1320_ _1324_ _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_50_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6257__A1 core_0.execute.alu_mul_div.div_cur\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8058_ _3469_ _3716_ _3734_ _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_242_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_242_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__A2 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7009_ _2009_ _2726_ _2937_ _2075_ _2938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_214_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_214_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6009__A1 net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_170_Right_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_214_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7757__A1 core_0.execute.rf.reg_outputs\[11\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_219_3142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7509__A1 core_0.ew_reg_ie\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__A3 _0960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4991__A1 _1163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8182__A1 _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6732__A2 _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_19_i_clk clknet_4_3__leaf_i_clk clknet_leaf_19_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_80_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6496__A1 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8237__A2 _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6799__A2 _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7996__A1 _3420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_148_2292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8235__B _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7748__A1 _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__A2 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4710_ core_0.fetch.out_buffer_valid _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_17_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5690_ _1403_ _1694_ _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8173__A1 _3472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ core_0.execute.rf.reg_outputs\[2\]\[5\] net250 _0716_ _0829_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6723__A2 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7360_ _3278_ _2483_ _3280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4572_ _0765_ net195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_142_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5931__B1 _1787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6311_ core_0.execute.alu_mul_div.div_cur\[9\] _2219_ _0999_ _2292_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8476__A2 _4048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7291_ _3071_ net236 _1999_ _3072_ _3073_ _3213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_13_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6487__A1 _2428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9030_ _0057_ clknet_leaf_91_i_clk core_0.fetch.out_buffer_data_instr\[18\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6242_ _2219_ _2226_ _2227_ _2230_ _0145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4498__B1 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8228__A2 core_0.execute.alu_mul_div.cbit\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6173_ core_0.execute.alu_mul_div.div_cur\[11\] _1835_ _2162_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_237_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6239__A1 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5124_ core_0.decode.i_instr_l\[1\] _1233_ _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_224_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5055_ _1086_ _1220_ _1221_ _1162_ net168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__5462__A2 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7739__A1 _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4670__B1 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8814_ _4316_ _4341_ _0606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_204_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8400__A2 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clone41_I net337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_rebuffer69_I _0682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_139_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7984__B _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8745_ _4293_ _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5957_ _1945_ _1946_ _1947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_175_2617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4973__A1 core_0.fetch.prev_request_pc\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4908_ core_0.fetch.prev_request_pc\[14\] _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8676_ core_0.execute.sreg_irq_pc.o_d\[7\] _4209_ _4241_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5888_ _1876_ _1877_ _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8164__A1 _3459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7506__A4 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7627_ core_0.execute.rf.reg_outputs\[14\]\[7\] _3482_ _3486_ _3487_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4839_ _0893_ net57 _1019_ _1020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__7911__A1 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7558_ core_0.execute.rf.reg_outputs\[15\]\[5\] _3429_ _3422_ _3436_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_214_3083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6509_ _1759_ _2349_ _2444_ _2449_ _2450_ _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_31_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7489_ core_0.dec_rf_ie\[13\] core_0.ew_reg_ie\[13\] _2421_ _3378_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9228_ _0239_ clknet_leaf_144_i_clk core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_219_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_2746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5150__A1 _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9159_ _0170_ clknet_leaf_75_i_clk core_0.execute.mem_stage_pc\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8219__A2 _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7978__A1 _3462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9290__CLK clknet_leaf_155_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6782__C _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5453__A2 _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8055__B _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_2927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5398__C _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6402__A1 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_197_2875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6953__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4964__A1 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8155__A1 net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7902__A1 _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6303__B _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4716__A1 net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_6 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7418__B1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5692__A2 _1696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7969__A1 core_0.execute.rf.reg_outputs\[5\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_206_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5589__B _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer18 net208 net246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_178_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer29 _1798_ net317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__4652__B1 _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6860_ _2450_ _2791_ _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_202_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7197__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8394__A1 _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_140_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5811_ _0954_ _0955_ _1790_ _1801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_202_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9013__CLK clknet_leaf_92_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6791_ _1899_ _1999_ _2724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6944__A2 _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8530_ net72 _4113_ _4114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_8_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5742_ core_0.execute.sreg_priv_control.o_d\[15\] _1700_ _1732_ _1697_ _1733_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8146__A1 net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8461_ _4052_ _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8697__A2 _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5673_ _1535_ _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_115_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7412_ _2124_ core_0.execute.alu_mul_div.mul_res\[15\] _3331_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4707__A1 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4512__I _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Right_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4624_ _0813_ net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_44_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8392_ _1540_ _4002_ _4003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_170_2547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_2558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7343_ net75 _2995_ _3264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5380__A1 _1289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4555_ core_0.execute.rf.reg_outputs\[7\]\[12\] _0683_ _0703_ core_0.execute.rf.reg_outputs\[15\]\[12\]
+ _0750_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xmax_cap220 _0704_ net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_96_1663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8449__A2 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7274_ _1684_ core_0.execute.sreg_irq_pc.o_d\[11\] _3197_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4486_ _0660_ _0662_ _0684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_9013_ _0040_ clknet_leaf_92_i_clk core_0.fetch.out_buffer_data_instr\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6439__I net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5132__A1 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6225_ _2165_ _2175_ _2189_ _2213_ _2214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_110_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6156_ _1519_ _0713_ _2145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5107_ _1230_ _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_225_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ core_0.execute.rf.reg_outputs\[7\]\[3\] _1773_ _2077_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5038_ core_0.fetch.prev_request_pc\[4\] _1207_ core_0.fetch.prev_request_pc\[5\]
+ _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_181_2687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I i_core_int_sreg[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_196_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4643__B1 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6989_ core_0.execute.alu_mul_div.i_mul core_0.execute.alu_mul_div.mul_res\[4\] _2919_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_216_3101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8728_ _4204_ _4283_ _4284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9506__CLK clknet_leaf_122_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8659_ _1658_ _4223_ _4227_ _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_192_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6699__A1 core_0.execute.rf.reg_outputs\[1\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6699__B2 core_0.execute.rf.reg_outputs\[3\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5371__A1 _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7733__I _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7112__A2 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5123__A1 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8860__A2 _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput76 net76 dbg_pc[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput87 net87 dbg_r0[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_227_3241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5674__A2 _1670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput98 net98 dbg_r0[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7889__B _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6285__S _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6623__A1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5426__A2 _1322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_243_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_199_2904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7908__I _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_238_3370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8128__A1 core_0.execute.rf.reg_outputs\[1\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_59_Right_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_1939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6968__B _2896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5362__A1 _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8300__B2 _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5163__I core_0.execute.alu_mul_div.i_div vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8851__A2 _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6010_ _1874_ _1999_ _2000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5665__A2 _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I i_core_int_sreg[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_68_Right_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8603__A2 _2556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6614__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__A2 _1297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7961_ core_0.execute.rf.reg_outputs\[5\]\[4\] _3679_ _3677_ _3680_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4625__B1 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6912_ _2571_ _2841_ _2842_ _2843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4507__I net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7892_ _3447_ _3628_ _3639_ _0386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_178_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8367__A1 _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9631_ _0641_ clknet_leaf_100_i_clk net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6843_ core_0.execute.sreg_irq_pc.o_d\[1\] _2774_ _2775_ core_0.execute.pc_high_out\[1\]
+ _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9562_ _0572_ clknet_leaf_73_i_clk core_0.execute.sreg_irq_pc.o_d\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4928__A1 core_0.fetch.prev_request_pc\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5766__C _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6774_ _2422_ _2706_ _2707_ _0200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8119__A1 core_0.execute.rf.reg_outputs\[1\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4928__B2 core_0.fetch.prev_request_pc\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Right_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7590__A2 _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8513_ _2399_ _4091_ _4099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_73_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5725_ _0777_ _1699_ _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_9493_ _0503_ clknet_leaf_22_i_clk net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_134_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8444_ _1680_ _4031_ core_0.execute.alu_mul_div.div_res\[15\] _4038_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5656_ _1591_ core_0.fetch.out_buffer_data_pred _1664_ _1665_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7342__A2 core_0.execute.sreg_irq_pc.o_d\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4607_ core_0.execute.rf.reg_outputs\[2\]\[8\] net312 _0715_ _0798_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8649__I core_0.dec_wfi vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_211_3042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8375_ _3979_ _3974_ _3987_ _3988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5587_ _1440_ core_0.fetch.submitable _1624_ _0096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7326_ _3060_ _2934_ _3246_ _3063_ _3247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4538_ core_0.execute.rf.reg_outputs\[5\]\[13\] _0677_ _0720_ core_0.execute.rf.reg_outputs\[4\]\[13\]
+ _0734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input59_I i_req_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5105__A1 core_0.decode.i_instr_l\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7257_ _2567_ _3031_ _3180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4469_ _0666_ _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_86_Right_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_183_2705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6208_ core_0.execute.alu_mul_div.div_cur\[9\] net234 _2197_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7188_ _2524_ _3112_ _1326_ _3113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9059__CLK clknet_leaf_92_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6139_ _2128_ core_0.execute.alu_mul_div.div_cur\[0\] _2129_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_222_3171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_222_3182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_95_Right_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7030__A1 net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7030__B2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4919__A1 core_0.fetch.prev_request_pc\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4919__B2 core_0.fetch.prev_request_pc\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_194_2845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7581__A2 _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8530__A1 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer9 net235 net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_58_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5344__A1 core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Left_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_210_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5647__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__A1 _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__C1 net336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6072__A2 net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_24_Left_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8349__A1 _2366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8349__B2 _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4771__B _0951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7021__A1 _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_13_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6542__I net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7572__A2 _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5510_ net52 _1554_ _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6490_ _2429_ _2430_ _2431_ _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_81_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5441_ _1535_ _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_14_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5886__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8160_ _3453_ _3780_ _3793_ _0500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5372_ _1437_ _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_93_1633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7088__A1 _2439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7111_ core_0.execute.alu_mul_div.div_res\[7\] _3038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_140_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8091_ _3462_ _3738_ _3753_ _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_238_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6835__A1 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7042_ _2499_ _2969_ _2491_ _2970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__B _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8993_ _0020_ clknet_leaf_141_i_clk core_0.dec_rf_ie\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_222_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7260__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7944_ core_0.execute.rf.reg_outputs\[6\]\[14\] _3650_ _3663_ _3669_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5810__A2 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7875_ core_0.execute.rf.reg_outputs\[7\]\[0\] _3629_ _3621_ _3630_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_194_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8153__B _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7012__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ _1768_ _2563_ _2759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_9614_ _0624_ clknet_leaf_132_i_clk core_0.dec_mem_width vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_rebuffer51_I net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7563__A2 core_0.ew_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8760__A1 _0825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9545_ _0555_ clknet_leaf_103_i_clk net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6757_ net1 _2691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__5574__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5068__I _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ core_0.execute.sreg_priv_control.o_d\[4\] _1701_ _1709_ _1698_ _1710_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_33_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9476_ _0486_ clknet_leaf_13_i_clk core_0.execute.rf.reg_outputs\[1\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6688_ net210 _2621_ _2622_ _2627_ _2628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8427_ _3038_ _4028_ _2258_ _0532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5639_ _1026_ _1628_ _1655_ _0117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5877__A2 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8358_ _3970_ _3971_ _3972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7079__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5017__B core_0.fetch.prev_request_pc\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7309_ _1684_ _3230_ _3231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output165_I net165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8815__A2 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8289_ _1535_ _3907_ _3908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5629__A2 _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6826__A1 _1768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_217_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone78_B _1847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8579__A1 _3150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A2 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_wire214_I _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8751__A1 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5565__A1 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7306__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_116_1909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_153_2350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6311__B _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8806__A2 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__A2 _0686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_184_Right_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6817__A1 _2480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_246_3480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7142__B _2795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5441__I _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7242__A1 _2708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6045__A2 net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5990_ core_0.execute.rf.reg_outputs\[6\]\[13\] net322 _1819_ core_0.execute.rf.reg_outputs\[12\]\[13\]
+ _1788_ core_0.execute.rf.reg_outputs\[3\]\[13\] _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__7793__A2 _3562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5597__B _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4941_ _1095_ _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_4_0__f_i_clk_I clknet_3_0_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_176_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6272__I _2229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7660_ core_0.execute.rf.reg_outputs\[13\]\[5\] _3504_ _3500_ _3506_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4872_ _0892_ _1052_ _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_191_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6611_ _2551_ _2552_ _2547_ _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_46_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5556__A1 _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7591_ _3387_ core_0.ew_data\[12\] _3449_ net24 _3462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__8701__B _4249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer1_I _0713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9330_ _0340_ clknet_leaf_8_i_clk core_0.execute.rf.reg_outputs\[10\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_171_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6542_ net99 _2484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9261_ _0271_ clknet_leaf_26_i_clk core_0.execute.rf.reg_outputs\[14\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6473_ core_0.dec_sys _0199_ _2417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_70_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8212_ _3835_ _3836_ core_0.execute.alu_mul_div.cbit\[2\] core_0.execute.alu_mul_div.cbit\[1\]
+ _3837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__5859__A2 _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5424_ _1232_ _1267_ _1280_ _1521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput200 net200 sr_bus_data_o[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9192_ _0203_ clknet_leaf_54_i_clk core_0.ew_data\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_100_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8143_ net95 _3781_ _3771_ _3784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5355_ core_0.decode.i_instr_l\[9\] core_0.decode.i_instr_l\[8\] core_0.decode.i_instr_l\[7\]
+ _1470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_2_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_2519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_151_Right_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6808__A1 _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8074_ _3427_ _3737_ _3744_ _0463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5286_ net192 net179 net178 net181 _1407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_10_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5087__A3 _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7025_ _2951_ _2952_ _2953_ _2954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_226_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_rebuffer99_I net345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7479__S _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7233__A1 core_0.execute.sreg_priv_control.o_d\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6036__A2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7233__B2 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8576__A4 _3256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8976_ _4455_ _4456_ _0653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_222_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8981__A1 _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7784__A2 _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7927_ core_0.execute.rf.reg_outputs\[6\]\[6\] _3657_ _3648_ _3660_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_178_2648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7858_ _3454_ _3606_ _3619_ _0372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7536__A2 _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5547__A1 core_0.fetch.prev_request_pc\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_191_2804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6809_ _1896_ _2738_ _2741_ _2742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5547__B2 net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7789_ _3463_ _3564_ _3579_ _0343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9528_ _0538_ clknet_leaf_120_i_clk core_0.execute.alu_mul_div.div_res\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9459_ _0469_ clknet_leaf_14_i_clk core_0.execute.rf.reg_outputs\[2\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4770__A2 core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_230_3270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4522__A2 _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_2777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7897__B _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__A1 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6027__A2 _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__B2 core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_204_2958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7775__A2 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4589__A2 net297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A1 _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8521__B _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6750__A3 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8948__S _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5710__A1 net251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4513__A2 _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5140_ _1263_ _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_244_3439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6266__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5071_ core_0.decode.input_valid core_0.decode.i_submit _0924_ _1228_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_236_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__A2 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8830_ _4316_ _4355_ _0608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_189_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7766__A2 _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5777__A1 _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8761_ core_0.execute.sreg_scratch.o_d\[7\] _4300_ _4304_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5973_ core_0.execute.rf.reg_outputs\[8\]\[14\] _1794_ _1776_ core_0.execute.rf.reg_outputs\[4\]\[14\]
+ _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_177_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7712_ _3460_ _3521_ _3535_ _0310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4924_ core_0.fetch.prev_request_pc\[7\] _1029_ _1039_ core_0.fetch.prev_request_pc\[6\]
+ _1104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8692_ _4210_ _4253_ _4254_ _0571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7518__A2 core_0.ew_data\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7643_ core_0.execute.rf.reg_outputs\[14\]\[15\] _3475_ _3486_ _3495_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4855_ _1017_ _1035_ _1036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8191__A2 _1835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_220_Right_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7574_ _3387_ core_0.ew_mem_width _3449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4786_ core_0.ew_reg_ie\[3\] _0966_ _0948_ core_0.ew_reg_ie\[0\] _0967_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_133_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9313_ _0323_ clknet_leaf_29_i_clk core_0.execute.rf.reg_outputs\[11\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_173_2589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6525_ _2459_ _2463_ _2466_ _2467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_145_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9244_ _0254_ clknet_leaf_10_i_clk core_0.execute.rf.reg_outputs\[15\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6456_ net77 _2411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_rebuffer14_I net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5407_ _1304_ _1491_ _1510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_9175_ _0186_ clknet_leaf_42_i_clk core_0.execute.prev_pc_high\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5701__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6387_ _1542_ _2360_ _2361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_135_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_208_3003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8126_ core_0.execute.rf.reg_outputs\[1\]\[11\] _3765_ _3771_ _3774_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_208_3014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5338_ _1278_ _1306_ _1454_ _1455_ _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA_input41_I i_req_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6257__A2 _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8057_ core_0.execute.rf.reg_outputs\[3\]\[14\] _3714_ _3730_ _3734_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5269_ core_0.execute.alu_flag_reg.o_d\[1\] core_0.execute.alu_flag_reg.o_d\[0\]
+ _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5081__I core_0.decode.i_instr_l\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7008_ _2009_ _1898_ _2735_ _2937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_126_2024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6009__A2 _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7206__A1 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7757__A2 _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5768__A1 _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8959_ _4447_ _0645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_219_3143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8706__A1 net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7509__A2 core_0.ew_reg_ie\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6980__A3 _2074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4991__A2 _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8182__A2 _2428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6193__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6496__A2 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7693__A1 core_0.execute.rf.reg_outputs\[12\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7404__C _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7445__A1 _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6248__A2 _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7996__A2 _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_214_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7748__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7646__I _3496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8173__A2 _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6550__I net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4640_ core_0.execute.rf.reg_outputs\[9\]\[5\] _0705_ net284 core_0.execute.rf.reg_outputs\[13\]\[5\]
+ _0828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_154_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5231__I0 core_0.ew_data\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7920__A2 _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Left_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4734__A2 _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4571_ net89 _0666_ _0764_ _0765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__5931__B2 core_0.execute.rf.reg_outputs\[3\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6310_ core_0.execute.alu_mul_div.div_cur\[8\] _2220_ _2256_ _2290_ _2291_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_188_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7290_ _2470_ _3212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_4_14__f_i_clk clknet_3_7_0_i_clk clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_229_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7684__A1 core_0.ew_reg_ie\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6487__A2 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6241_ _2229_ _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_40_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4498__A1 core_0.execute.rf.reg_outputs\[1\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4498__B2 core_0.execute.rf.reg_outputs\[10\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6172_ core_0.execute.alu_mul_div.div_cur\[11\] _1835_ _2161_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7436__A1 net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6239__A2 _0998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ _1240_ _1274_ _1278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_243_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ net79 _1085_ _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5998__A1 _0730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8936__A1 core_0.decode.i_imm_pass\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7739__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4670__B2 core_0.execute.rf.reg_outputs\[10\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8813_ core_0.execute.pc_high_out\[1\] _4327_ _4340_ _4341_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6947__B1 _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_133_i_clk clknet_4_6__leaf_i_clk clknet_leaf_133_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5956_ core_0.execute.rf.reg_outputs\[13\]\[11\] _1792_ _1815_ core_0.execute.rf.reg_outputs\[9\]\[11\]
+ _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8744_ _4293_ _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_clone34_I _0685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_2607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6962__A3 _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_2618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ core_0.fetch.prev_request_pc\[15\] _1023_ _1087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_61_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8675_ _1658_ _4236_ _4240_ _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_192_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5887_ core_0.execute.alu_flag_reg.o_d\[1\] core_0.dec_alu_carry_en _1877_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__8161__B _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8164__A2 _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4838_ _1017_ _1018_ _1019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7626_ _1430_ _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_173_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_148_i_clk clknet_4_0__leaf_i_clk clknet_leaf_148_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7911__A2 _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7557_ _3434_ _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5922__A1 _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4769_ core_0.dec_l_reg_sel\[1\] core_0.dec_l_reg_sel\[0\] _0950_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_105_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_214_3084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6508_ _2008_ _2102_ _2450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5009__C _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7488_ _3377_ _0244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_160_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7675__A1 _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6439_ net85 _2401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9227_ _0238_ clknet_leaf_142_i_clk core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_2094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9158_ _0169_ clknet_leaf_56_i_clk core_0.execute.mem_stage_pc\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_186_2747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7427__A1 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8109_ _3420_ _3759_ _3764_ _0478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9089_ _0114_ clknet_leaf_94_i_clk core_0.decode.i_imm_pass\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_243_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7978__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_242_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6650__A2 _2591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8927__A1 _1494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4661__A1 net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9585__CLK clknet_leaf_108_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_201_2928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_195_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_197_2876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4964__A2 _1143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7466__I _2418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8155__A2 _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7902__A2 _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4716__A2 net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5913__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_7 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7666__A1 core_0.execute.rf.reg_outputs\[13\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7418__B2 net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_241_3409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7969__A2 _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8091__A1 _3462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer19 _1833_ net247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_221_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8918__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_50_i_clk clknet_4_11__leaf_i_clk clknet_leaf_50_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__B2 core_0.execute.rf.reg_outputs\[13\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_85_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ core_0.execute.rf.reg_outputs\[2\]\[0\] _1797_ _1799_ core_0.execute.rf.reg_outputs\[6\]\[0\]
+ _1800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_159_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6790_ _1875_ _1956_ _2723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5741_ net229 _1704_ _1732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_225_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8146__A2 _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8460_ _4040_ _2136_ _4052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_84_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5672_ _1672_ _1676_ _1677_ _1678_ _0127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_44_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7411_ _1829_ _1888_ _3311_ _1292_ _3329_ _3330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_115_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4623_ net100 net324 _0812_ _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_8391_ _1674_ _1829_ _2372_ _1973_ _3982_ _1545_ _4002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_60_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4707__A2 _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_2548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7342_ _1684_ core_0.execute.sreg_irq_pc.o_d\[13\] _3263_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4554_ core_0.execute.rf.reg_outputs\[2\]\[12\] _0673_ _0693_ core_0.execute.rf.reg_outputs\[1\]\[12\]
+ _0749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmax_cap221 _0694_ net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_96_1664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7273_ net73 _2995_ _3195_ _2893_ _3196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4485_ net297 _0683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
X_9012_ _0039_ clknet_leaf_97_i_clk core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6224_ _2210_ _2211_ _2212_ _2213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_111_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5132__A2 _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7409__A1 _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6155_ _2142_ _2143_ _2144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_225_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5106_ _1260_ _1261_ _1262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_32_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6086_ _1930_ _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5037_ _1147_ _1148_ _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_212_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_18_i_clk clknet_4_3__leaf_i_clk clknet_leaf_18_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_181_2688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_rebuffer81_I _0685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4643__A1 core_0.execute.rf.reg_outputs\[7\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4643__B2 core_0.execute.rf.reg_outputs\[10\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7995__B _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7487__S _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8385__A2 _3995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6988_ _2759_ _2901_ _2917_ _2918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_105_1771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_216_3102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8727_ _4282_ _4283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5939_ net314 net200 _1928_ _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_35_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6148__A1 _2130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7345__B1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8658_ _4212_ core_0.execute.mem_stage_pc\[3\] _4202_ _4226_ _4227_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_91_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output195_I net304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6699__A2 _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7896__A1 _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7609_ _3475_ _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_63_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8589_ _4166_ _4165_ _1371_ _4167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_105_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7499__I1 core_0.ew_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_79_Left_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output72_I net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_227_3231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput77 net77 dbg_pc[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_227_3242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput88 net88 dbg_r0[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput99 net99 dbg_r0[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__5470__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4882__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8066__B _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4594__B _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_145_2252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6623__A2 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7820__A1 core_0.execute.rf.reg_outputs\[9\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_199_2905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6387__A1 _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_88_Left_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_224_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_238_3371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8128__A2 _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6139__A1 _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7887__A1 core_0.execute.rf.reg_outputs\[7\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_2381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7639__A1 core_0.execute.rf.reg_outputs\[14\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8956__S _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_97_Left_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_239_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8300__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6311__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4873__A1 _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6075__B1 _1818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6614__A2 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7960_ _3671_ _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_221_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4625__A1 core_0.execute.rf.reg_outputs\[10\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__B2 core_0.execute.rf.reg_outputs\[9\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6911_ _1864_ _2571_ _2756_ _2842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7891_ core_0.execute.rf.reg_outputs\[7\]\[7\] _3634_ _3636_ _3639_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8704__B _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8367__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9630_ _0640_ clknet_leaf_97_i_clk net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6378__A1 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6842_ _1686_ _1410_ _2687_ _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_0_187_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6773_ core_0.ew_data\[0\] _2642_ _2707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4928__A2 _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9561_ _0571_ clknet_leaf_68_i_clk core_0.execute.sreg_irq_pc.o_d\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5050__A1 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8119__A2 _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__I _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4523__I _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8512_ _4095_ _4098_ _4051_ _0547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5724_ _1714_ _1720_ _0137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9492_ _0502_ clknet_leaf_17_i_clk net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_162_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7878__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_198_Right_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5655_ _0895_ _1345_ _1664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8443_ _2230_ _4037_ _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4606_ core_0.execute.rf.reg_outputs\[6\]\[8\] net223 _0699_ core_0.execute.rf.reg_outputs\[12\]\[8\]
+ _0797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8374_ core_0.execute.alu_mul_div.mul_res\[13\] _3986_ _3987_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5353__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5586_ _1134_ _1369_ _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_211_3043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7325_ _2568_ _3104_ _3245_ _3060_ _3246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4537_ core_0.execute.rf.reg_outputs\[11\]\[13\] _0680_ _0716_ _0733_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4561__B1 _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7256_ _2588_ _3177_ _3178_ _3179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_111_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5105__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6302__A1 _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4468_ _0661_ _0663_ _0665_ _0666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_217_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_183_2706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6207_ core_0.execute.alu_mul_div.div_cur\[9\] net234 _2196_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7187_ _2529_ _3066_ _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4864__A1 _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8055__A1 core_0.execute.rf.reg_outputs\[3\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6138_ core_0.execute.alu_mul_div.i_mod _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_213_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6605__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7802__A1 core_0.execute.rf.reg_outputs\[9\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6069_ _1770_ _2056_ _2057_ _2058_ _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_107_1800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_222_3172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output208_I net245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7030__A2 _2829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_140_2193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4919__A2 _1020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_194_2835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5041__A1 _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_194_2846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7869__A1 _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_165_Right_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5465__S _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7744__I _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5344__A2 _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__A2 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6844__A2 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4855__A1 _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8046__A1 core_0.execute.rf.reg_outputs\[3\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6057__B1 net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_204_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8349__A2 _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7021__A2 _2949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_158_2410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5032__A1 _1106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5583__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5883__B net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_132_Right_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5440_ core_0.execute.alu_mul_div.cbit\[3\] _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_2_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4543__B1 _0710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_2__f_i_clk clknet_3_1_0_i_clk clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5371_ _1464_ _1481_ _0022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_93_1623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_1634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7110_ _1290_ _3035_ _3036_ _1742_ _3037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_112_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8285__A1 _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8090_ core_0.execute.rf.reg_outputs\[2\]\[12\] _3743_ _3745_ _3753_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_196_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5099__A1 core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7041_ _2502_ _2907_ _2969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6835__A2 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8037__A1 _3427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8992_ _0019_ clknet_leaf_127_i_clk core_0.dec_rf_ie\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__A2 _2366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7943_ _3466_ _3652_ _3668_ _0408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7874_ _3627_ _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7012__A2 _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9613_ _0623_ clknet_leaf_19_i_clk core_0.dec_mem_long vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6825_ _2587_ _2757_ _2758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_65_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_1741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8760__A2 _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9544_ _0554_ clknet_leaf_103_i_clk net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__5574__A2 _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6756_ core_0.execute.pc_high_out\[0\] _1686_ _1410_ _2687_ _2690_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_46_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5707_ _0848_ _1704_ _1709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6687_ _2146_ net210 _2627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_190_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9475_ _0485_ clknet_leaf_16_i_clk core_0.execute.rf.reg_outputs\[1\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7564__I _3440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8426_ _1537_ _1680_ _4013_ _4028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5638_ core_0.decode.i_imm_pass\[13\] _1645_ _1655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5569_ _1345_ _1551_ _1614_ _0088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8357_ _1536_ _3868_ _3971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7079__A2 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7308_ net74 _2995_ _3229_ _2893_ _3230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8276__A1 _3893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8815__A3 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8288_ _1538_ _3905_ _3906_ _3907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_229_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6908__I _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6826__A2 _2563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7239_ _3156_ _3161_ _3127_ _3163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5812__I _1801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_224_3201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9176__CLK clknet_leaf_42_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6039__B1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_234_Right_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5801__A3 _1790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_240_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8200__A1 core_0.execute.alu_mul_div.mul_res\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5014__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5259__I core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8751__A2 _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_235_3330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__B1 _0686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8519__B _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8806__A3 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_246_3470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8019__A1 core_0.execute.rf.reg_outputs\[4\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_164_2480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7242__A2 net307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_201_Right_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4940_ _1104_ _1119_ _1120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_188_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ core_0.fetch.out_buffer_data_instr\[16\] _1052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_157_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ _2470_ _2471_ _2543_ _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_129_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7590_ _3403_ _3460_ _3461_ _0262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6753__A1 _1687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6541_ _2423_ _2482_ _2483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_6_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6472_ _2416_ _0188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9260_ _0270_ clknet_leaf_10_i_clk core_0.execute.rf.reg_outputs\[14\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8211_ net94 _1813_ _2109_ _2114_ _1668_ _3836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_5423_ _1278_ _1282_ _1301_ _1306_ _1520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_9191_ _0202_ clknet_leaf_57_i_clk core_0.ew_data\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xoutput201 net201 sr_bus_data_o[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_112_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8258__A1 _3835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5354_ _1464_ _1469_ _0017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8142_ _3408_ _3780_ _3783_ _0492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7333__B _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8073_ core_0.execute.rf.reg_outputs\[2\]\[4\] _3743_ _3730_ _3744_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5285_ net180 net183 net182 _1406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4819__A1 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7024_ core_0.execute.alu_mul_div.div_cur\[5\] _2128_ _2953_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_199_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7233__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8430__A1 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8975_ core_0.decode.i_instr_l\[10\] _1293_ _1271_ _4456_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5244__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7926_ _3435_ _3651_ _3659_ _0400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6992__A1 _2921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_131_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_2649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7857_ core_0.execute.rf.reg_outputs\[8\]\[9\] _3613_ _3609_ _3619_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_182_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6808_ _1896_ _2739_ _2740_ _2741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_163_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5547__A2 _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_191_2805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6744__A1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7788_ core_0.execute.rf.reg_outputs\[10\]\[12\] _3570_ _3568_ _3579_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9527_ _0537_ clknet_leaf_119_i_clk core_0.execute.alu_mul_div.div_res\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6739_ core_0.dec_sreg_jal_over _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_135_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5807__I _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__I _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8497__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9458_ _0468_ clknet_leaf_24_i_clk core_0.execute.rf.reg_outputs\[2\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8409_ _4015_ _4016_ _4017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_230_3271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9389_ _0399_ clknet_leaf_23_i_clk core_0.execute.rf.reg_outputs\[6\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_2778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_56_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A3 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_204_2959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8972__A2 _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6373__I net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_17_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6983__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8724__A2 _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__A1 _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7160__A1 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5710__A2 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8964__S _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5452__I _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ _0911_ net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6992__B core_0.execute.alu_mul_div.i_mod vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6671__B1 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_231_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8760_ _0825_ _4294_ _4303_ _4287_ _0590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5777__A2 _1766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5972_ _1961_ _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_75_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7711_ core_0.execute.rf.reg_outputs\[12\]\[11\] _3526_ _3528_ _3535_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4923_ _1090_ _1100_ _1102_ _1103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_176_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8691_ core_0.execute.sreg_irq_pc.o_d\[9\] _4210_ _3797_ _4254_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7642_ _3470_ _3477_ _3494_ _0281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4854_ core_0.fetch.out_buffer_data_instr\[26\] _1035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7328__B _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7573_ _3397_ _3447_ _3448_ _0258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4785_ _0954_ _0955_ _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_133_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9312_ _0322_ clknet_leaf_26_i_clk core_0.execute.rf.reg_outputs\[11\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6524_ _2464_ _2465_ _2466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_1695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9243_ _0253_ clknet_leaf_2_i_clk core_0.execute.rf.reg_outputs\[15\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _1163_ _2386_ _2410_ _0178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6886__C _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5406_ _1444_ _1453_ _1506_ _1508_ _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_2
X_9174_ _0185_ clknet_leaf_42_i_clk core_0.execute.prev_pc_high\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6386_ _2358_ _1962_ _2359_ _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__8159__B _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5701__A2 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_208_3004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8125_ _3456_ _3760_ _3773_ _0485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5337_ _1239_ _1261_ _1280_ _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_239_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7998__B _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8056_ _3465_ _3716_ _3733_ _0456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5268_ core_0.execute.alu_flag_reg.o_d\[4\] _1387_ _1388_ _1375_ core_0.dec_jump_cond_code\[2\]
+ _1389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__8651__A1 _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input34_I i_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7007_ _2502_ _2935_ _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_199_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5199_ _1342_ _0005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_242_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7206__A2 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8403__A1 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5217__A1 core_0.ew_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6965__A1 _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__A2 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8958_ net179 core_0.decode.i_imm_pass\[11\] _1263_ _4447_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_195_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__C _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7909_ core_0.execute.rf.reg_outputs\[7\]\[15\] _3627_ _3648_ _3649_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8889_ core_0.execute.pc_high_buff_out\[5\] _4385_ _1430_ _4405_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8706__A2 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7509__A3 core_0.ew_reg_ie\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_219_3144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9364__CLK clknet_leaf_7_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8341__C _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_232_3300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4728__B1 _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7390__A1 core_0.ew_data\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6193__A2 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_150_2310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7142__A1 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8890__A1 _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Left_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7693__A2 _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4597__B _0788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7445__A2 _3040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8642__A1 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5456__A1 _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7701__B _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_2450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6956__A1 core_0.ew_data\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_201_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8532__B _3156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7381__A1 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6184__A2 _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5231__I1 core_0.ew_data\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7381__B2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4570_ _0758_ _0763_ _0764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5392__B1 _1494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5931__A2 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6240_ _2228_ _2229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8881__A1 core_0.execute.pc_high_buff_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7684__A2 _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4498__A2 _0693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5695__A1 _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6892__B1 _2768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6171_ core_0.execute.alu_mul_div.div_cur\[9\] net234 _2160_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_110_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _1272_ _1276_ _1277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_237_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7436__A2 _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8707__B _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5053_ _1219_ _1063_ _1145_ _1220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7611__B _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5998__A2 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_108_Left_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8936__A2 _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4670__A2 _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8812_ net215 _4328_ _4326_ _4339_ _4340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6947__A1 core_0.execute.alu_flag_reg.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9387__CLK clknet_leaf_2_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8743_ _1419_ _1420_ _3044_ _4293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_153_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5955_ core_0.execute.rf.reg_outputs\[8\]\[11\] _1794_ _1776_ core_0.execute.rf.reg_outputs\[4\]\[11\]
+ _1945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_175_2608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5470__I1 net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4906_ _1085_ _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__8244__S0 core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8674_ _1662_ core_0.execute.mem_stage_pc\[6\] _4238_ _4239_ _4201_ _4240_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_47_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5886_ _1875_ _1812_ _1876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_192_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7625_ _3441_ _3476_ _3485_ _0273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4837_ core_0.fetch.out_buffer_data_instr\[28\] _1018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7372__A1 _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_117_Left_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_117_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7556_ _3382_ core_0.ew_data\[5\] _3433_ _3434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_160_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5922__A2 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4768_ _0947_ _0948_ _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_214_3085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6507_ _2445_ _2447_ _2448_ _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_31_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7487_ core_0.dec_rf_ie\[12\] core_0.ew_reg_ie\[12\] _2421_ _3377_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4699_ core_0.execute.rf.reg_outputs\[7\]\[0\] net296 net284 core_0.execute.rf.reg_outputs\[13\]\[0\]
+ _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_31_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9226_ _0237_ clknet_leaf_138_i_clk core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_101_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ _2399_ _2385_ _2400_ _0171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8872__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7675__A2 _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5686__A1 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6883__B1 _2759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5092__I net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9157_ _0168_ clknet_leaf_70_i_clk core_0.execute.mem_stage_pc\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_186_2748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6369_ _1541_ _1669_ _1812_ _2343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_87_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8108_ core_0.execute.rf.reg_outputs\[1\]\[3\] _3760_ _3756_ _3764_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5025__C _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9088_ _0113_ clknet_leaf_91_i_clk core_0.decode.i_imm_pass\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5438__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7521__B _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_126_Left_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_8039_ _3434_ _3715_ _3724_ _0448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_215_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6137__B _2126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A2 net324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_2929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_197_2877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_rebuffer102_I _2528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_135_Left_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_213_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7363__A1 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8578__I _3188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_8 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8863__A1 _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7666__A2 _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_144_Left_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7418__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6477__I0 core_0.dec_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8091__A2 _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__A2 _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6929__A1 _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_179_Right_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7657__I _3496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5601__A1 _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _1714_ _1731_ _0142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7354__A1 core_0.ew_data\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5671_ _1540_ _1534_ _1678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5177__I core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6157__A2 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7410_ _2795_ _3314_ _3321_ _3328_ _3329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_154_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4622_ _0806_ _0811_ _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_170_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8390_ core_0.execute.alu_mul_div.mul_res\[14\] _2375_ _4001_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_170_2549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7341_ _2703_ _3261_ _3262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4553_ core_0.execute.rf.reg_outputs\[14\]\[12\] _0686_ _0700_ core_0.execute.rf.reg_outputs\[12\]\[12\]
+ _0748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7606__B _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5905__I _1753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap222 _0676_ net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_96_1665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7272_ _3193_ _3194_ _3195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4484_ net293 _0663_ _0678_ _0682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__5668__A1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9011_ _0038_ clknet_leaf_100_i_clk core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6223_ _2176_ _2179_ _2183_ _2212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_12_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6154_ _1855_ _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_209_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5105_ core_0.decode.i_instr_l\[1\] _1241_ _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6085_ _2074_ _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__8082__A2 _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5036_ net82 _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__7060__C _2759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_181_2689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4643__A2 _0683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5840__A1 _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_rebuffer74_I core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_146_Right_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8172__B _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6987_ _2905_ _2908_ _2916_ _2917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_105_1772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8726_ net209 _2778_ _4282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5938_ net314 _1690_ _1928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_216_3103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8657_ _4224_ _4063_ _4225_ _1662_ _4226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6148__A2 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7345__A1 core_0.execute.sreg_priv_control.o_d\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5869_ _1838_ _1844_ _1849_ _1859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_90_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7345__B2 net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7608_ core_0.ew_reg_ie\[14\] _3395_ _3475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_118_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7896__A2 _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8588_ core_0.dec_alu_flags_ie _4166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_161_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4954__I0 net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output188_I net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7539_ _3381_ _3417_ _3418_ _3419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5815__I core_0.execute.rf.reg_outputs\[12\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8845__A1 _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7648__A2 _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5659__A1 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9209_ _0220_ clknet_leaf_52_i_clk net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput78 net78 dbg_pc[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_227_3232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput89 net89 dbg_r0[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_101_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_228_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4882__A2 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7251__B core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8073__A2 _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7820__A2 _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_2906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__A2 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Right_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8082__B _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8781__B1 _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6381__I net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_238_3372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7336__A1 core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7887__A2 _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5898__A1 _1766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8101__I _3758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8836__A1 core_0.execute.pc_high_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7639__A2 _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_132_i_clk clknet_4_6__leaf_i_clk clknet_leaf_132_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6311__A2 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4873__A2 net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8064__A2 _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_206_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6075__A1 core_0.execute.rf.reg_outputs\[9\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6075__B2 core_0.execute.rf.reg_outputs\[12\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7811__A2 _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4625__A2 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6910_ net267 _2840_ _2841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_222_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7890_ _3441_ _3628_ _3638_ _0385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6841_ _1686_ _1689_ _2676_ _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_193_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7575__B2 net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9560_ _0570_ clknet_leaf_73_i_clk core_0.execute.sreg_irq_pc.o_d\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_202_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _2672_ net193 _2705_ _2706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8511_ _4047_ _4097_ _4098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_44_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5723_ core_0.execute.sreg_priv_control.o_d\[9\] _1701_ _1719_ _1698_ _1720_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7327__A1 net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9491_ _0501_ clknet_leaf_17_i_clk net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__8524__B1 _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8442_ _4026_ _4031_ core_0.execute.alu_mul_div.div_res\[14\] _4037_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5654_ _1003_ _1663_ _1435_ _0124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7878__A2 _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5889__A1 _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4605_ core_0.execute.rf.reg_outputs\[14\]\[8\] net309 net286 core_0.execute.rf.reg_outputs\[13\]\[8\]
+ _0796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8373_ _1536_ _3886_ _3985_ _3986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5585_ _1623_ _0095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_211_3044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8827__A1 _4324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7324_ _2571_ _3177_ _3244_ _2568_ _3245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4561__A1 core_0.execute.rf.reg_outputs\[5\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4536_ core_0.execute.rf.reg_outputs\[3\]\[13\] _0698_ _0708_ core_0.execute.rf.reg_outputs\[13\]\[13\]
+ _0732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _2588_ _3102_ _3178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4467_ net273 net301 _0665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_clone94_I _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ core_0.execute.alu_mul_div.div_cur\[15\] net238 _2195_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_183_2707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7186_ _2728_ _3069_ _3107_ _3110_ _3111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_55_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_215_Right_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8055__A2 _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6137_ core_0.execute.alu_mul_div.div_res\[0\] _1742_ _2126_ _2127_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_225_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6066__A1 core_0.execute.rf.reg_outputs\[7\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7802__A2 _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6068_ core_0.execute.rf.reg_outputs\[13\]\[6\] _1791_ net331 core_0.execute.rf.reg_outputs\[4\]\[6\]
+ _2058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_107_1801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5813__A1 _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _1192_ _1049_ _1158_ _1193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_222_3173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__A1 _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output103_I net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4714__I net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5041__A2 _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_194_2836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8709_ _4212_ core_0.execute.mem_stage_pc\[12\] _4201_ _4268_ _4269_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_181_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7318__A1 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7869__A2 _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8818__A1 _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7760__I _3562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_64_i_clk clknet_4_9__leaf_i_clk clknet_leaf_64_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8046__A2 _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_216_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6057__A1 core_0.execute.rf.reg_outputs\[5\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6309__C _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6057__B2 core_0.execute.rf.reg_outputs\[10\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__A2 net312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_69_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_79_i_clk clknet_4_14__leaf_i_clk clknet_leaf_79_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_231_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_2411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5032__A2 _1149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7309__A1 _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4791__A1 core_0.ew_reg_ie\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7156__B core_0.execute.alu_mul_div.i_div vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6532__A2 _2371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_17_i_clk clknet_4_3__leaf_i_clk clknet_leaf_17_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8809__A1 core_0.execute.pc_high_buff_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A1 core_0.execute.rf.reg_outputs\[6\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ core_0.dec_rf_ie\[12\] _1438_ _1472_ _1480_ _1481_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4543__B2 core_0.execute.rf.reg_outputs\[8\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8766__I _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_2540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7040_ _2968_ _0205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_239_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8037__A2 _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8991_ _0018_ clknet_leaf_141_i_clk core_0.dec_rf_ie\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7796__A1 _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7942_ core_0.execute.rf.reg_outputs\[6\]\[13\] _3657_ _3663_ _3668_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7873_ _3627_ _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_194_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4534__I net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9612_ _0622_ clknet_leaf_109_i_clk core_0.dec_wfi vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6824_ net270 _2588_ _2756_ _2757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_187_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_102_1731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9543_ _0553_ clknet_4_14__leaf_i_clk net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_161_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6755_ _1405_ _1689_ _2676_ _2689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_18_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4782__A1 _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5706_ _1608_ _1708_ _0131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_73_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9474_ _0484_ clknet_leaf_16_i_clk core_0.execute.rf.reg_outputs\[1\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6686_ _2626_ _0192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer37_I net264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8425_ _2230_ _4027_ _0531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5637_ _1020_ _1628_ _1654_ _0116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8356_ _1539_ _3968_ _3969_ _1679_ _3970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_131_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5731__B1 _1700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ core_0.fetch.out_buffer_data_pred _1556_ _1614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input64_I i_req_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7307_ _3227_ _3228_ _3229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4519_ _0715_ _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__7580__I _3453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8287_ _1538_ _3854_ _3906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5499_ _1041_ _1551_ _1576_ _0056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6287__A1 _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7238_ _3127_ _3156_ _3161_ _3162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_111_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_113_1871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4709__I net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7169_ _2703_ _3085_ _3092_ _3094_ _3095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_129_2056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7787__A1 _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8984__B1 _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_201_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_206_2990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7539__A1 _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6211__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_235_3331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5476__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6762__A2 _2689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_153_2352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6514__A2 _1925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7711__A1 core_0.execute.rf.reg_outputs\[12\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__B2 core_0.execute.rf.reg_outputs\[14\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_246_3460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_224_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7778__A1 core_0.execute.rf.reg_outputs\[10\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_2481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4870_ _1016_ _1030_ _1040_ _1050_ _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_87_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6753__A2 net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6540_ net241 _1988_ _2482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_40_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5961__B1 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6471_ core_0.execute.trap_flag _0199_ _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_113_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7702__A1 _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8210_ net87 _1813_ _1783_ _1810_ core_0.execute.alu_mul_div.cbit\[0\] _3835_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_125_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5422_ _1518_ _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_9190_ _0201_ clknet_leaf_51_i_clk core_0.ew_data\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5713__B1 _1700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput202 net202 sr_bus_data_o[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_113_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8141_ net94 _3781_ _3771_ _3783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8258__A2 _3836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5353_ core_0.dec_rf_ie\[7\] _1438_ _1462_ _1468_ _1469_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6269__A1 _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8072_ _3736_ _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6808__A3 _2740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5284_ _1404_ _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4819__A2 core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7023_ core_0.execute.alu_mul_div.div_res\[5\] _1742_ _0997_ _2952_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_4_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5492__A2 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7769__A1 core_0.execute.rf.reg_outputs\[10\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8974_ core_0.dec_jump_cond_code\[3\] _1251_ _4455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7925_ core_0.execute.rf.reg_outputs\[6\]\[5\] _3657_ _3648_ _3659_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6992__A2 core_0.execute.alu_mul_div.i_div vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7856_ _3451_ _3606_ _3618_ _0371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8194__A1 _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_6_0_i_clk clknet_0_i_clk clknet_3_6_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6807_ _1875_ _2102_ _2740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_147_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_191_2806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7787_ _3460_ _3564_ _3578_ _0342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4999_ _1020_ _1176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7941__A1 _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6744__A2 _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4755__A1 core_0.ew_reg_ie\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9526_ _0536_ clknet_leaf_119_i_clk core_0.execute.alu_mul_div.div_res\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6738_ core_0.dec_mem_access _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_190_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9457_ _0467_ clknet_leaf_62_i_clk core_0.execute.rf.reg_outputs\[2\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6669_ _0947_ _0954_ _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_45_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8408_ _2140_ _1543_ _3878_ _4016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_103_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9388_ _0398_ clknet_4_3__leaf_i_clk core_0.execute.rf.reg_outputs\[6\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_230_3272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output170_I net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8339_ _3878_ _3929_ _3953_ _3954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5823__I _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_2779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_245_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6680__A1 _2614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5698__C _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6027__A4 _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A2 _2492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4994__A1 _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8802__C _4324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8090__B _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6735__A2 _2668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7932__A1 _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7418__C _2689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__A2 _4076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5171__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5733__I net197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_166_2510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7999__A1 _3427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6120__B1 _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8660__A2 _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6671__A1 core_0.execute.rf.reg_outputs\[7\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6671__B2 core_0.execute.rf.reg_outputs\[5\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4793__B _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__B1 net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_232_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5971_ _0950_ _0951_ _1961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_150_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7710_ _3457_ _3521_ _3534_ _0309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4922_ _1088_ _1016_ _1101_ _1102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8690_ _4249_ core_0.execute.mem_stage_pc\[9\] _4252_ _4253_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8176__A1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8712__C _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7641_ core_0.execute.rf.reg_outputs\[14\]\[14\] _3475_ _3486_ _3494_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4853_ _1033_ _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_145_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5908__I _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7572_ core_0.execute.rf.reg_outputs\[15\]\[7\] _3429_ _3422_ _3448_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4784_ core_0.ew_reg_ie\[1\] _0963_ _0964_ core_0.ew_reg_ie\[2\] _0965_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_144_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9311_ _0321_ clknet_4_8__leaf_i_clk core_0.execute.rf.reg_outputs\[11\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6523_ _2425_ _2424_ _2465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_42_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9242_ _0252_ clknet_leaf_2_i_clk core_0.execute.rf.reg_outputs\[15\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6454_ core_0.execute.mem_stage_pc\[14\] _1433_ _2404_ _2410_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7151__A2 _3069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _1313_ _1502_ _1507_ _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_9173_ _0184_ clknet_leaf_42_i_clk core_0.execute.prev_pc_high\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6739__I core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6385_ _2046_ _2053_ _2359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8124_ core_0.execute.rf.reg_outputs\[1\]\[10\] _3765_ _3771_ _3773_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7063__C _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5336_ _1240_ _1443_ _1454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_208_3005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_110_1830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8055_ core_0.execute.rf.reg_outputs\[3\]\[13\] _3722_ _3730_ _3733_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5267_ _1376_ core_0.execute.alu_flag_reg.o_d\[1\] _1388_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6662__A1 core_0.decode.oc_alu_mode\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7006_ _2497_ _2907_ _2935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_215_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5198_ _1338_ _1251_ _1293_ _1341_ _1342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_126_2026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input27_I i_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8403__A2 _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5217__A2 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8957_ _4446_ _0644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_167_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7908_ _3647_ _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8888_ net204 _4387_ _4403_ _4404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_219_3145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7509__A4 core_0.ew_reg_ie\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7839_ _3512_ _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_65_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_1970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8962__I0 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_232_3301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7390__A2 _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9509_ _0519_ clknet_leaf_124_i_clk core_0.execute.alu_mul_div.mul_res\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_199_Left_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_150_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_150_2311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output95_I net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8642__A2 _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_243_3430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6653__A1 _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4664__B1 net302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6384__I net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_161_2440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6405__A1 _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6317__C _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6956__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8158__A1 _3450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7148__C _3073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5916__B1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7381__A2 _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5392__A1 core_0.decode.i_imm_pass\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5392__B2 core_0.decode.i_instr_l\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_2580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8330__A1 core_0.execute.alu_mul_div.mul_res\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7164__B _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__A1 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8881__A2 _4385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6892__A1 net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5695__A2 _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6892__B2 core_0.execute.sreg_scratch.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6170_ _2157_ _2158_ _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_198_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5121_ _1244_ _1274_ _1275_ _1267_ _1276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_236_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6644__A1 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5052_ core_0.fetch.prev_request_pc\[2\] _1218_ _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_127_Right_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4655__B1 _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8811_ _4328_ _4338_ _4339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_204_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8723__B _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_212_Left_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_153_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6947__A2 _2770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4958__A1 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8742_ _4291_ _4292_ _1435_ _0583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5954_ net89 _1772_ _1944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8149__A1 net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4905_ core_0.fetch.pc_flush_override core_0.decode.i_flush _1085_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_175_2609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8673_ _4224_ _4085_ _1662_ _4239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_47_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ _1874_ _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__8244__S1 core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8944__I0 net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7624_ core_0.execute.rf.reg_outputs\[14\]\[6\] _3482_ _3467_ _3485_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4836_ core_0.fetch.out_buffer_valid _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_35_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_99_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7555_ _3381_ _3431_ _3432_ _3433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5383__A1 _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4767_ core_0.dec_l_reg_sel\[1\] core_0.dec_l_reg_sel\[0\] _0948_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_132_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_3075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _1895_ _2341_ _2448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_214_3086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7486_ _3376_ _0243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_160_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8321__A1 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4698_ core_0.execute.rf.reg_outputs\[5\]\[0\] _0677_ net347 core_0.execute.rf.reg_outputs\[15\]\[0\]
+ _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XPHY_EDGE_ROW_221_Left_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9225_ _0236_ clknet_leaf_137_i_clk core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_160_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6437_ core_0.execute.mem_stage_pc\[7\] _2395_ _2387_ _2400_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8872__A2 _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6883__A1 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5686__A2 net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6883__B2 net282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9156_ _0167_ clknet_leaf_67_i_clk core_0.execute.mem_stage_pc\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6368_ _2337_ _2341_ _1541_ _2342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_2749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8107_ _3414_ _3759_ _3763_ _0477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7802__B _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5319_ _1436_ _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9087_ _0112_ clknet_leaf_93_i_clk core_0.decode.i_imm_pass\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_227_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6299_ _1547_ _2280_ _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_227_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6635__A1 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5438__A2 net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8038_ core_0.execute.rf.reg_outputs\[3\]\[5\] _3722_ _3718_ _3724_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_243_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__B _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4646__B1 net321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_230_Left_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9331__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5041__C _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6399__B1 _2371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_201_2919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6938__A2 core_0.execute.alu_mul_div.mul_res\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_195_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5610__A2 _1640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_197_2878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9481__CLK clknet_leaf_16_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8560__A1 _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7363__A2 _2370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5374__A1 _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_229_Right_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8312__A1 _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_9 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5283__I net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8863__A2 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6874__A1 _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8379__A1 core_0.execute.alu_mul_div.mul_res\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A2 net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5458__I _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5670_ _1671_ _1675_ _1677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7354__A2 _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8551__A1 _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4621_ _0807_ _0808_ _0809_ _0810_ _0811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__5365__A1 _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7673__I _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7340_ _1317_ _3259_ _3260_ _3261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_13_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ _0743_ _0744_ _0745_ _0746_ _0747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__8303__A1 _3901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xmax_cap223 _0669_ net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7271_ core_0.execute.sreg_irq_pc.o_d\[11\] _3042_ _3044_ core_0.execute.sreg_scratch.o_d\[11\]
+ _3194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4483_ core_0.execute.rf.reg_outputs\[5\]\[15\] _0677_ _0680_ core_0.execute.rf.reg_outputs\[11\]\[15\]
+ _0681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_12_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9010_ _0037_ clknet_leaf_109_i_clk core_0.dec_pc_inc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5668__A2 _1674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6865__A1 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _2182_ _2190_ _2211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8718__B _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7622__B _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6153_ core_0.execute.alu_mul_div.div_cur\[14\] _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_209_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6617__A1 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5104_ _1242_ core_0.decode.i_instr_l\[2\] _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6084_ _1687_ net217 _1519_ _2074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XANTENNA__4628__B1 _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5035_ _1202_ _1165_ _1204_ _1205_ _1080_ net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_224_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_2679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__A2 net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _2912_ _2915_ _2916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_rebuffer67_I net294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8790__A1 _4249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7593__A2 _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5937_ _1898_ _1912_ _1926_ _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_105_1773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8725_ _4280_ _4281_ _0577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_193_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_216_3104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8656_ net80 _1740_ _1707_ _4205_ _4225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5868_ _1857_ _1761_ _1328_ _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__7345__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8542__A1 net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6002__C1 _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7607_ _3403_ _3473_ _3474_ _0266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4819_ core_0.decode.o_submit core_0.execute.alu_mul_div.i_mul _1000_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_173_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8587_ _4159_ _4165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_32_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5799_ core_0.execute.rf.reg_outputs\[5\]\[0\] _1785_ net340 core_0.execute.rf.reg_outputs\[9\]\[0\]
+ _1788_ core_0.execute.rf.reg_outputs\[3\]\[0\] _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_16_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7538_ net30 _1348_ _3418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7469_ core_0.dec_rf_ie\[3\] core_0.ew_reg_ie\[3\] _3366_ _3368_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6856__A1 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5659__A2 _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9208_ _0219_ clknet_leaf_52_i_clk net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9139_ _0151_ clknet_leaf_115_i_clk core_0.execute.alu_mul_div.div_cur\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xoutput79 net79 dbg_pc[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_227_3233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5831__I _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6608__A1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4619__B1 net308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7281__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4890__I0 net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_19_Right_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8781__A1 core_0.execute.irq_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8781__B2 core_0.execute.sreg_irq_flags.o_d\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_211_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_122_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5595__A1 core_0.decode.i_instr_l\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_3373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8533__A1 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7336__A2 core_0.execute.alu_mul_div.mul_res\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7707__B _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_2383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8836__A2 _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Right_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A1 _2692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_47_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6075__A2 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_234_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_37_Right_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7024__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6840_ _2769_ _2772_ _2773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_159_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6771_ _2702_ _2704_ core_0.dec_mem_access _2705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5586__A1 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8510_ net277 _4048_ _3040_ _2133_ _4096_ _4097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_186_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5722_ _0789_ _1699_ _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4794__C1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9490_ _0500_ clknet_leaf_21_i_clk net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_17_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7327__A2 _2371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8524__B2 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8441_ _2230_ _4036_ _0538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7617__B _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5653_ _1662_ _1002_ net20 core_0.ew_submit _1663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_5_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9535__D _0545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ core_0.execute.rf.reg_outputs\[1\]\[8\] net308 _0702_ core_0.execute.rf.reg_outputs\[15\]\[8\]
+ _0795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5889__A2 _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8372_ _1539_ _3930_ _3984_ _1536_ _3985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_46_Right_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5584_ _1068_ core_0.decode.i_instr_l\[6\] _1368_ _1623_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_170_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_211_3045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7323_ net270 _3243_ _2571_ _3244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4535_ core_0.execute.rf.reg_outputs\[10\]\[13\] _0695_ _0705_ core_0.execute.rf.reg_outputs\[9\]\[13\]
+ _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_229_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6838__A1 _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7254_ _1769_ _3176_ _1864_ _3177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4466_ core_0.dec_r_reg_sel\[0\] _0664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_111_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7352__B core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6205_ core_0.execute.alu_mul_div.div_cur\[14\] _2143_ _2194_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5651__I net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_2708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7185_ _1885_ _2462_ _2457_ _1880_ _3109_ _3110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_55_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6136_ _1743_ _2123_ _2125_ _0996_ _2126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_225_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7263__A1 _2859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6066__A2 _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7263__B2 _1768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6067_ core_0.execute.rf.reg_outputs\[8\]\[6\] net346 _2057_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_55_Right_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_107_1802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5018_ _1151_ _1191_ _1192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_212_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5813__A2 _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_222_3174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7015__A1 core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__A2 _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A3 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8763__A1 core_0.execute.sreg_scratch.o_d\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5098__I core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6969_ _2699_ _2898_ _2899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_140_2195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_2837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8708_ _4203_ _4127_ _4266_ _4267_ _1661_ _4268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_48_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8515__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5329__A1 _1239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8639_ _4209_ _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_36_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Right_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4552__A2 _0744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_73_Right_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_219_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6057__A2 net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_i_clk i_clk clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_231_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_204_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_2412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8313__S _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8506__A1 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Right_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6368__I0 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__A2 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4543__A2 _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5740__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8809__A2 _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8268__B _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_169_2541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6296__A2 _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Right_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_226_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I i_core_int_sreg[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8990_ _0017_ clknet_leaf_127_i_clk core_0.dec_rf_ie\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7796__A2 _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7941_ _3463_ _3652_ _3667_ _0407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7398__I _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4815__I core_0.execute.alu_mul_div.i_div vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7872_ core_0.ew_reg_ie\[7\] _3395_ _3627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_210_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7548__A2 core_0.ew_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9611_ _0621_ clknet_leaf_106_i_clk core_0.decode.input_valid vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5559__A1 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6823_ _1329_ _2446_ _2739_ _2756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_202_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_1732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9542_ _0552_ clknet_leaf_82_i_clk net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6754_ core_0.execute.pc_high_buff_out\[0\] net185 _2680_ _2687_ _2688_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_163_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7347__B _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5705_ core_0.execute.sreg_long_ptr_en _1701_ _1707_ _1698_ _1708_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_163_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6685_ _2625_ net131 _2419_ _2626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9473_ _0483_ clknet_leaf_37_i_clk core_0.execute.rf.reg_outputs\[1\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4782__A2 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5636_ core_0.decode.i_imm_pass\[12\] _1645_ _1654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8424_ _4015_ _4026_ core_0.execute.alu_mul_div.div_res\[6\] _4027_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_162_Left_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7720__A2 _3519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8355_ _1539_ _3915_ _3969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5567_ _1608_ _1613_ _0087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_170_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5731__A1 net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5731__B2 core_0.execute.sreg_priv_control.o_d\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7861__I _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7306_ core_0.execute.sreg_priv_control.o_d\[12\] _1693_ _3042_ core_0.execute.sreg_irq_pc.o_d\[12\]
+ _3228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_229_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4518_ net326 _0671_ _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_8286_ _3878_ _3884_ _3904_ _3905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5498_ net45 _1554_ _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input57_I i_req_data[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7237_ _1684_ _3160_ _3161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_245_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2_0_i_clk clknet_0_i_clk clknet_3_2_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_113_1872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7168_ _2703_ _3093_ _3094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7236__A1 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6039__A2 _1791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7236__B2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6119_ _2105_ _2106_ _2107_ _2108_ _2109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_171_Left_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7099_ core_0.decode.oc_alu_mode\[6\] _2439_ _3023_ _3025_ _3026_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_241_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7787__A2 _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8984__B2 _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_206_2980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A3 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_131_i_clk clknet_4_6__leaf_i_clk clknet_leaf_131_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6211__A2 _1833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4758__C1 _0930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_235_3332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_193_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_180_Left_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5970__A1 _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_146_i_clk clknet_4_1__leaf_i_clk clknet_leaf_146_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7711__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_2353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4525__A2 net296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5722__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7771__I _3562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8088__B _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_246_3461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7227__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7720__B _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9415__CLK clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7778__A2 _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8975__A1 core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_2482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_189_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6450__A2 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8270__C _3830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6470_ _2415_ _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_82_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7163__B1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7702__A2 _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5421_ _1517_ _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_70_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__A1 net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__B2 core_0.execute.sreg_priv_control.o_d\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput203 net203 sr_bus_data_o[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8140_ _3401_ _3780_ _3782_ _0491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5352_ _1439_ _1465_ _1440_ _1468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_23_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6269__A2 _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8071_ _3420_ _3737_ _3742_ _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5283_ net185 _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_239_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7022_ _1290_ core_0.execute.alu_mul_div.mul_res\[5\] _2950_ _1314_ _2951_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_52_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7218__A1 _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7769__A2 _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8973_ _1439_ _1230_ _1272_ _4454_ _0652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_223_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6441__A2 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7924_ _3428_ _3651_ _3658_ _0399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8718__A1 _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7855_ core_0.execute.rf.reg_outputs\[8\]\[8\] _3613_ _3609_ _3618_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6760__I core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6806_ _1899_ _2115_ _2739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_175_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4998_ net74 _1175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__8180__C _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7786_ core_0.execute.rf.reg_outputs\[10\]\[11\] _3570_ _3568_ _3578_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_2807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7941__A2 _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6744__A3 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9525_ _0535_ clknet_leaf_115_i_clk core_0.execute.alu_mul_div.div_res\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6737_ _2616_ _2669_ _2670_ _2671_ _0198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4755__A2 _0928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_63_i_clk clknet_4_9__leaf_i_clk clknet_leaf_63_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6668_ core_0.execute.rf.reg_outputs\[1\]\[0\] _2608_ _2609_ core_0.execute.rf.reg_outputs\[3\]\[0\]
+ _2610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9456_ _0466_ clknet_leaf_24_i_clk core_0.execute.rf.reg_outputs\[2\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5619_ _1368_ _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_8407_ _1679_ _2215_ _2216_ _4015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__5704__A1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6599_ _2465_ _2535_ _2540_ _2541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9387_ _0397_ clknet_leaf_2_i_clk core_0.execute.rf.reg_outputs\[6\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_230_3273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_78_i_clk clknet_4_14__leaf_i_clk clknet_leaf_78_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8338_ _3878_ _3952_ _3953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output163_I net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8269_ _3877_ _3888_ _3889_ _3890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8636__B _4201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7209__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6432__A2 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_16_i_clk clknet_4_3__leaf_i_clk clknet_leaf_16_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_241_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8709__A1 _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7932__A2 _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7715__B _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7207__S _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_108_Right_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5171__A2 _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_2500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7999__A2 _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6120__A1 core_0.execute.rf.reg_outputs\[9\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6120__B2 core_0.execute.rf.reg_outputs\[10\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6671__A2 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_205_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6959__B1 _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7620__A1 core_0.execute.rf.reg_outputs\[14\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5970_ _1896_ _1927_ _1959_ _1960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7471__I1 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ core_0.fetch.prev_request_pc\[15\] _1023_ _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4985__A2 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8176__A2 _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4852_ net50 core_0.fetch.out_buffer_data_instr\[21\] _1017_ _1033_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_177_2640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7640_ _3466_ _3477_ _3493_ _0280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6187__A1 core_0.execute.alu_mul_div.div_cur\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7923__A2 _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7571_ _3446_ _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_27_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4737__A2 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4783_ _0957_ _0958_ _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_129_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5934__A1 _1916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6522_ net247 _1941_ _2464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_55_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9310_ _0320_ clknet_leaf_26_i_clk core_0.execute.rf.reg_outputs\[11\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7687__A1 core_0.execute.rf.reg_outputs\[12\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6453_ _1170_ _2386_ _2409_ _0177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9241_ _0251_ clknet_leaf_2_i_clk core_0.execute.rf.reg_outputs\[15\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5698__B1 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ _1240_ _1458_ _1507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9172_ _0183_ clknet_leaf_42_i_clk core_0.execute.prev_pc_high\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6384_ net100 _2358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_140_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7439__A1 _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8123_ _3453_ _3759_ _3772_ _0484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5335_ _1300_ _1452_ _1453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_11_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_208_3006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8054_ _3462_ _3716_ _3732_ _0455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5266_ core_0.dec_jump_cond_code\[1\] _1374_ _1387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_110_1831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7005_ _2568_ _2757_ _2933_ _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA_clkbuf_leaf_95_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5197_ _1256_ _1295_ _1340_ _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8939__A1 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4673__A1 net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer97_I _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7462__I1 core_0.ew_reg_ie\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8956_ net178 core_0.decode.i_imm_pass\[10\] _1263_ _4446_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_203_2950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8903__C _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7907_ _0891_ _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_195_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8887_ _0917_ _4383_ _4403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_219_3135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6178__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_219_3146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7838_ _3402_ _3606_ _3608_ _0363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5225__I0 core_0.ew_data\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7914__A2 _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_1960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8962__I1 core_0.decode.i_imm_pass\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__A2 _0904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5925__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_232_3302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7769_ core_0.execute.rf.reg_outputs\[10\]\[3\] _3564_ _3568_ _3569_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9508_ _0518_ clknet_leaf_124_i_clk core_0.execute.alu_mul_div.mul_res\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_22_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7535__B _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9439_ _0449_ clknet_leaf_46_i_clk core_0.execute.rf.reg_outputs\[3\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__9260__CLK clknet_leaf_10_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_2312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6350__A1 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output88_I net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__A1 core_0.execute.rf.reg_outputs\[12\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_243_3431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__A2 _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7850__A1 _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4664__B2 core_0.execute.rf.reg_outputs\[1\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_2441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6405__A2 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7496__I _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8158__A2 _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7905__A2 _3627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5916__A1 core_0.execute.rf.reg_outputs\[3\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__B1 _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5392__A2 _1488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7669__A1 _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_172_2581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6892__A2 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_117_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5120_ core_0.decode.i_instr_l\[3\] core_0.decode.i_instr_l\[2\] _1234_ _1275_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_20_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8276__B _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5051_ core_0.fetch.prev_request_pc\[1\] core_0.fetch.prev_request_pc\[0\] _1218_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7841__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4655__A1 core_0.execute.rf.reg_outputs\[1\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4655__B2 core_0.execute.rf.reg_outputs\[15\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8810_ _4335_ _4336_ _4337_ _4338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_189_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8741_ core_0.execute.sreg_jtr_buff.o_d\[2\] _4217_ _1415_ _4292_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4958__A2 _1135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5953_ _1874_ _1942_ _1943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8149__A2 _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _1084_ net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_192_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8672_ _1202_ _4217_ _4237_ _4219_ _4238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_62_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5884_ _1869_ _1873_ _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_75_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7623_ _3435_ _3476_ _3484_ _0272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4835_ net60 core_0.fetch.out_buffer_data_instr\[30\] _0892_ _1016_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__9283__CLK clknet_leaf_7_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7554_ net32 _1348_ _3432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4766_ core_0.dec_l_reg_sel\[2\] _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XANTENNA__5383__A2 _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6505_ _1884_ _1877_ _2446_ _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__4591__B1 _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_3076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7485_ core_0.dec_rf_ie\[11\] core_0.ew_reg_ie\[11\] _3366_ _3376_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4697_ net215 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XANTENNA__8321__A2 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9224_ _0235_ clknet_leaf_137_i_clk core_0.ew_reg_ie\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6436_ net84 _2399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_rebuffer12_I _1837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_219_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6367_ _2338_ _1962_ _2339_ _2340_ _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_9155_ _0166_ clknet_leaf_68_i_clk core_0.execute.mem_stage_pc\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_132_2097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_2739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8106_ core_0.execute.rf.reg_outputs\[1\]\[2\] _3760_ _3756_ _3763_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5318_ _1007_ _1228_ _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8085__A1 _3453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9086_ _0111_ clknet_leaf_93_i_clk core_0.decode.i_imm_pass\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6298_ _2159_ _2279_ _2280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_228_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7832__A1 core_0.execute.rf.reg_outputs\[9\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5249_ _1370_ net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8037_ _3427_ _3715_ _3723_ _0447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_215_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4646__A1 core_0.execute.rf.reg_outputs\[1\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4646__B2 core_0.execute.rf.reg_outputs\[12\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Left_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6399__A1 _1674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8939_ _1690_ _0038_ _4437_ _0635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6434__B _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5829__I _1818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_197_2879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_210_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_193_Right_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_49_Left_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8312__A2 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7823__A1 _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5834__B1 _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6328__C _2229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8379__A2 _3830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8543__C _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6344__B _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5062__A1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_43_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4620_ core_0.execute.rf.reg_outputs\[15\]\[7\] _0702_ _0715_ _0810_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4551_ core_0.execute.rf.reg_outputs\[5\]\[12\] _0677_ _0720_ core_0.execute.rf.reg_outputs\[4\]\[12\]
+ _0746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4573__B1 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_160_Right_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7270_ core_0.execute.sreg_priv_control.o_d\[11\] _1693_ _2996_ net3 _3193_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap224 _1786_ net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_96_1667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4482_ _0679_ _0680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_110_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6221_ _2209_ _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7903__B _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6865__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4876__A1 _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8067__A1 _3408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6152_ _1679_ _2140_ _1667_ _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_20_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_225_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5103_ _1243_ _1258_ _1259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6617__A2 _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7814__A1 _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6083_ _1895_ _2042_ _2072_ _1898_ _2073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4628__A1 core_0.execute.rf.reg_outputs\[7\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4628__B2 core_0.execute.rf.reg_outputs\[3\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5034_ _1038_ _1146_ _1164_ _1205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_212_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6985_ _1254_ _2495_ _2913_ _1749_ _2914_ _2915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5649__I _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_24_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8025__I _3714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8724_ core_0.execute.sreg_irq_pc.o_d\[15\] _4210_ _2387_ _4281_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7069__C _2689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5936_ _1874_ _1925_ _1926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_216_3105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8655_ _4205_ _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5867_ _1838_ _1844_ _1849_ _1856_ _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__6002__B1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8542__A2 _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6002__C2 core_0.execute.rf.reg_outputs\[3\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7606_ core_0.execute.rf.reg_outputs\[15\]\[15\] _3396_ _3467_ _3474_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6553__A1 _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ core_0.decode.o_submit _0998_ _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_145_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8586_ _4155_ _4157_ _4158_ _4163_ _4164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_133_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5798_ _1787_ _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_32_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_134_2115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7085__B core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7537_ net23 _1347_ _3417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4749_ net274 _0675_ _0930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_160_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7468_ _3367_ _0234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9207_ _0218_ clknet_leaf_52_i_clk net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7813__B _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6856__A2 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6419_ _2384_ _2385_ _2388_ _0164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4867__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7399_ _3317_ _1974_ _3071_ _3318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8058__A1 _3469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9138_ _0150_ clknet_leaf_115_i_clk core_0.execute.alu_mul_div.div_cur\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_227_3234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7805__A1 _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__B _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9069_ _0094_ clknet_leaf_111_i_clk core_0.decode.i_instr_l\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_243_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4619__B2 core_0.execute.rf.reg_outputs\[1\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7281__A2 _3192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5292__A1 _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5044__A1 _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8781__A2 net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4463__I _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6792__A1 _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5595__A2 _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_238_3363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_3374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8533__A2 _3155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_57_Left_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4555__B1 _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_2384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8049__A1 _3456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_66_Left_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_246_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7949__I _3671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8221__A1 _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7024__A2 _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A1 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5469__I _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6770_ _2130_ _2703_ _2704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_186_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6783__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5586__A2 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_75_Left_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5721_ _1714_ _1718_ _0136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4794__C2 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8524__A2 _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8440_ _4024_ _4031_ core_0.execute.alu_mul_div.div_res\[13\] _4036_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5652_ _1661_ _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6535__A1 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ _0790_ _0791_ _0792_ _0793_ _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8371_ _1544_ _3952_ _3983_ _1539_ _3984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5583_ _1268_ core_0.fetch.submitable _1622_ _0094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_211_3046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4534_ net91 _0730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7322_ _2714_ _2724_ _1329_ _3243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9321__CLK clknet_leaf_3_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7633__B _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7253_ _2721_ _2723_ _3176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4465_ net271 _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_13_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4849__A1 _1020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6204_ _2165_ _2192_ _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7184_ net213 _3072_ _3108_ net233 _3073_ _3109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XPHY_EDGE_ROW_84_Left_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5510__A2 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_2709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _2124_ core_0.execute.alu_mul_div.mul_res\[0\] _2125_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8460__A1 _4040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7263__A2 _3069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6066_ core_0.execute.rf.reg_outputs\[7\]\[6\] _1773_ _2056_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_225_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5274__A1 core_0.de_jmp_pred vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5017_ core_0.fetch.prev_request_pc\[8\] _1150_ core_0.fetch.prev_request_pc\[9\]
+ _1191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_213_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5813__A3 _0960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_222_3175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8183__C _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8212__A1 _3835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7015__A2 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5026__A1 core_0.fetch.prev_request_pc\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5379__I _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8763__A2 _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_93_Left_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6774__A1 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6968_ _2833_ _2881_ _2896_ _2898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5577__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8707_ net74 _1740_ _4205_ _4267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_194_2838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5919_ _1905_ _1906_ _1907_ _1908_ _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6899_ _1401_ _2822_ _2828_ _2830_ _2831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__8515__A2 _4040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8638_ _0900_ _4200_ _4209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_180_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5329__A2 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5328__B _1289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output193_I net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8569_ net230 _4048_ _3340_ _4046_ _4148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_51_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_1932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7543__B _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6829__A2 _2761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5501__A2 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8451__A1 _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_235_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8203__A1 _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5017__A1 core_0.fetch.prev_request_pc\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6765__A1 core_0.dec_sreg_load vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5568__A2 _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_2413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8506__A2 _4040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6368__I1 _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4528__B1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7190__A1 _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5752__I _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_2542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8690__A1 _4249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4700__B1 net321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7245__A2 _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7940_ core_0.execute.rf.reg_outputs\[6\]\[12\] _3657_ _3663_ _3667_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7871_ _3473_ _3607_ _3626_ _0378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9610_ _0620_ clknet_leaf_57_i_clk core_0.execute.pc_high_buff_out\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6822_ core_0.decode.oc_alu_mode\[3\] _1888_ _2755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_159_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6756__A1 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8731__C _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9541_ _0551_ clknet_leaf_71_i_clk net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_102_1733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6753_ _1687_ net191 _1406_ _1407_ _2687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_147_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5704_ net217 _1704_ _1707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9472_ _0482_ clknet_leaf_37_i_clk core_0.execute.rf.reg_outputs\[1\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_174_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6508__A1 _2008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6684_ _2623_ _2624_ _2625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8423_ _1540_ _2354_ _1545_ _4026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_116_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5635_ _1057_ _1628_ _1653_ _0115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8354_ _2357_ _2368_ _3878_ _3968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5566_ core_0.fetch.prev_request_pc\[15\] _1082_ _1083_ net166 _1613_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5731__A2 _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8459__B _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7305_ net4 _2996_ _3044_ core_0.execute.sreg_scratch.o_d\[12\] _3227_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4517_ net92 _0714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_130_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5497_ _1052_ _1551_ _1575_ _0055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8285_ _3878_ _3903_ _3904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7236_ net72 _2995_ _3159_ _2893_ _3160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_113_1873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7167_ _3086_ _3091_ _3051_ _3093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_226_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7236__A2 _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6118_ core_0.execute.rf.reg_outputs\[15\]\[1\] _0945_ _1797_ core_0.execute.rf.reg_outputs\[2\]\[1\]
+ _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_129_2058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ _2054_ _1889_ _3024_ net287 _3025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_241_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8984__A2 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6049_ _2027_ _2038_ _2039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_198_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_206_2981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output206_I net268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6747__A1 core_0.execute.sreg_irq_flags.o_d\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4758__B1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4758__C2 core_0.ew_reg_ie\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_235_3333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_2343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_2354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4897__B _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5722__A2 _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8672__A1 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_246_3462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7227__A2 core_0.execute.alu_mul_div.mul_res\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8975__A2 _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_2483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6986__A1 _2912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4852__S _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8551__C _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5410__A1 core_0.decode.i_instr_l\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5410__B2 core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5961__A2 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7163__A1 core_0.execute.sreg_priv_control.o_d\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7163__B2 net15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5420_ core_0.dec_r_bus_imm _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__5713__A2 _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7183__B _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput204 net204 sr_bus_data_o[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5351_ _1464_ _1467_ _0016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6578__I net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8663__A1 _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5415__C _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8070_ core_0.execute.rf.reg_outputs\[2\]\[3\] _3738_ _3730_ _3742_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5282_ _1402_ _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_121_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8793__I _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7021_ _2124_ _2949_ _2950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8972_ core_0.dec_jump_cond_code\[2\] _1250_ _4454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7923_ core_0.execute.rf.reg_outputs\[6\]\[4\] _3657_ _3648_ _3658_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_210_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8742__B _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6729__A1 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7854_ _3447_ _3606_ _3617_ _0370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_194_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6805_ _1883_ _2492_ _2737_ _2738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7785_ _3457_ _3564_ _3577_ _0341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _1170_ _1165_ _1172_ _1174_ _1080_ net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_46_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_2808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9524_ _0534_ clknet_leaf_115_i_clk core_0.execute.alu_mul_div.div_res\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6744__A4 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6736_ net137 _2419_ _2671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_91_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer42_I _0666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9455_ _0465_ clknet_leaf_24_i_clk core_0.execute.rf.reg_outputs\[2\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6667_ _0943_ _0954_ _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XPHY_EDGE_ROW_12_Left_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_8406_ _2258_ _4014_ _0525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5618_ _1060_ _1615_ _1644_ _0107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9386_ _0396_ clknet_leaf_1_i_clk core_0.execute.rf.reg_outputs\[6\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5704__A2 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6598_ _2464_ _2533_ _2540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_230_3274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8337_ _1542_ _2366_ _3951_ _3952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5549_ core_0.fetch.prev_request_pc\[7\] _1595_ _1084_ net173 _1604_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_103_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8268_ _3877_ _3888_ _3828_ _3889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output156_I net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7219_ net248 _1942_ _3143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8199_ _3823_ _3824_ _3825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8406__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6437__B _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5341__B _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_21_Left_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8371__C _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Left_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7696__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5171__A3 _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7448__A2 _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8645__A1 _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5459__A1 net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_2501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7731__B _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__A2 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_236_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4682__A2 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6959__A1 core_0.execute.pc_high_buff_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6959__B2 core_0.execute.pc_high_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7620__A2 _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7957__I _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5631__A1 _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5482__I1 net39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4920_ _1091_ _1098_ _1099_ _1100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_113_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4851_ _1031_ _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_157_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_2641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6187__A2 _2008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7570_ _3382_ core_0.ew_data\[7\] _3445_ _3446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_51_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4782_ _0957_ _0955_ _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__5934__A2 _1923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _2460_ _2461_ _2462_ _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_7_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9240_ _0250_ clknet_leaf_45_i_clk net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8884__A1 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6452_ core_0.execute.mem_stage_pc\[13\] _2395_ _2404_ _2409_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7687__A2 _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5698__A1 net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5698__B2 core_0.execute.sreg_priv_control.o_d\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _1325_ _1445_ _1459_ _1505_ _1506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_9171_ _0182_ clknet_leaf_43_i_clk core_0.execute.prev_pc_high\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6383_ _2354_ _2355_ _2356_ _2357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_140_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8122_ core_0.execute.rf.reg_outputs\[1\]\[9\] _3765_ _3771_ _3772_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7439__A2 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5334_ _1247_ _1319_ _1450_ _1451_ _1452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__8636__A1 _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_208_3007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_2770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7641__B _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8053_ core_0.execute.rf.reg_outputs\[3\]\[12\] _3722_ _3730_ _3732_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5940__I _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5265_ core_0.execute.alu_flag_reg.o_d\[3\] _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_130_i_clk clknet_4_6__leaf_i_clk clknet_leaf_130_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_227_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7004_ _2567_ _2932_ _2933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5196_ _1240_ _1302_ _1339_ _1340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_214_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5870__A1 _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8939__A2 _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4673__A2 _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8028__I _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_145_i_clk clknet_4_1__leaf_i_clk clknet_leaf_145_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7611__A2 _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8955_ _4445_ _0643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_195_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_203_2951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7906_ _3470_ _3629_ _3646_ _0393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_211_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8886_ _4386_ _4401_ _4402_ _0617_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8191__C _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_174_Right_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7088__B _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_219_3136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7837_ core_0.execute.rf.reg_outputs\[8\]\[0\] _3607_ _3595_ _3608_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7375__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6178__A2 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_121_1961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7768_ _3512_ _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_18_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9507_ _0517_ clknet_leaf_122_i_clk core_0.execute.alu_mul_div.mul_res\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_80_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ _2654_ _2655_ _2656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7816__B _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7127__A1 _2708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7699_ core_0.execute.rf.reg_outputs\[12\]\[5\] _3526_ _3528_ _3529_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9438_ _0448_ clknet_leaf_44_i_clk core_0.execute.rf.reg_outputs\[3\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__8875__A1 _0904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7678__A2 _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_2313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5689__A1 core_0.dec_sreg_store vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9369_ _0379_ clknet_leaf_4_i_clk core_0.execute.rf.reg_outputs\[7\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_131_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5055__C _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9555__CLK clknet_leaf_64_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7551__B _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__A2 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_243_3432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7850__A2 _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__A2 net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_2442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7602__A2 _3396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5613__A1 core_0.decode.i_imm_pass\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_201_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_141_Right_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7366__A1 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6169__A2 net306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8563__B1 net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7366__B2 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5916__A2 _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__A1 core_0.execute.pc_high_buff_out\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__B2 core_0.execute.sreg_scratch.o_d\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7669__A2 _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_172_2571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_2582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5144__A3 _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8618__A1 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_237_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5050_ _1086_ _1216_ _1217_ _1162_ net169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__7841__A2 _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4655__A2 _0693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5852__A1 _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_62_i_clk clknet_4_9__leaf_i_clk clknet_leaf_62_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_205_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6805__B _2737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5604__A1 _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8740_ _0901_ _1418_ _4291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5952_ _1941_ _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4958__A3 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_77_i_clk clknet_4_14__leaf_i_clk clknet_leaf_77_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_62_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5080__A2 _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4903_ _1083_ _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8671_ net279 _0900_ _4237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5883_ _1870_ _1871_ net314 _1872_ _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_192_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7622_ core_0.execute.rf.reg_outputs\[14\]\[5\] _3482_ _3467_ _3484_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4834_ _1011_ _1014_ _1015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7553_ net25 _1347_ _3431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7109__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4765_ core_0.dec_mem_long core_0.execute.sreg_long_ptr_en _0946_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_28_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6580__A2 _2521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _1755_ net344 _1812_ _2446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_214_3077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7484_ _3375_ _0242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4696_ net94 _0667_ _0875_ _0879_ _0880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_132_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9223_ _0234_ clknet_leaf_139_i_clk core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6435_ _1202_ _2385_ _2398_ _0170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_141_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_i_clk clknet_4_3__leaf_i_clk clknet_leaf_15_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8609__A1 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9154_ _0165_ clknet_leaf_67_i_clk core_0.execute.mem_stage_pc\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6366_ _2110_ _2111_ _2112_ _2113_ _2340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_60_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_228_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8105_ _3408_ _3759_ _3762_ _0476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5317_ _1253_ _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_228_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9085_ _0110_ clknet_leaf_93_i_clk core_0.decode.i_imm_pass\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8085__A2 _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6297_ _2166_ _2274_ _2168_ _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6096__A1 core_0.execute.rf.reg_outputs\[13\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__B1 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8036_ core_0.execute.rf.reg_outputs\[3\]\[4\] _3722_ _3718_ _3723_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_243_Right_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_243_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5248_ net154 core_0.ew_addr_high\[0\] _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7832__A2 _3584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input32_I i_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4646__A2 net302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5843__A1 net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5179_ _1231_ _1325_ _1327_ _0001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6399__A2 _2370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7597__I _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output119_I net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8938_ core_0.decode.i_imm_pass\[1\] _1293_ _4437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8869_ core_0.execute.pc_high_buff_out\[0\] _4386_ _3797_ _4390_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clone39_C _1862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7899__A2 _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4957__I0 net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6450__B _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_104_Left_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8076__A2 _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6087__A1 core_0.execute.rf.reg_outputs\[7\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7823__A2 _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_210_Right_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__B2 core_0.execute.rf.reg_outputs\[10\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_113_Left_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_221_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7587__B2 net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5062__A2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8387__I0 core_0.execute.alu_mul_div.mul_res\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_2600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8000__A2 _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6011__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6562__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4550_ core_0.execute.rf.reg_outputs\[11\]\[12\] _0680_ _0716_ _0745_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4481_ _0661_ net298 _0678_ _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xmax_cap225 _1784_ net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7511__A1 _3386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ _2207_ _2208_ _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_5__f_i_clk clknet_3_2_0_i_clk clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4876__A2 net56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6151_ _2139_ _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_21_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8067__A2 _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5102_ _1257_ _1241_ _1258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6617__A3 _2556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6082_ _1895_ _2071_ _2072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7814__A2 _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4628__A2 net297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5033_ _1146_ _1203_ _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_225_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7027__B1 _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8734__C _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7578__A1 _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6984_ _2492_ _2755_ _2452_ core_0.decode.oc_alu_mode\[9\] _2914_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_200_2910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6250__A1 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8723_ _4212_ core_0.execute.mem_stage_pc\[15\] _4202_ _4279_ _4280_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_24_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5935_ net101 _1772_ _1924_ _1925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_48_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_216_3106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8654_ core_0.execute.sreg_irq_pc.o_d\[3\] _4210_ _4223_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5866_ _1851_ net212 _1855_ _1856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_0_63_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6002__A1 core_0.execute.rf.reg_outputs\[6\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6002__B2 core_0.execute.rf.reg_outputs\[12\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7605_ _3472_ _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4817_ _0996_ _0997_ _0998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_146_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8585_ _2989_ _3035_ _4162_ _4163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_146_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7750__A1 _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6553__A2 _2492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ _0960_ _0951_ _1787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_16_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7536_ _3397_ _3415_ _3416_ _0253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4748_ core_0.ew_reg_ie\[6\] _0928_ _0663_ _0929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7467_ core_0.dec_rf_ie\[2\] core_0.ew_reg_ie\[2\] _3366_ _3367_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7502__A1 _0946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4679_ _0860_ _0861_ _0862_ _0863_ _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_98_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Right_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_9206_ _0217_ clknet_leaf_52_i_clk net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6418_ core_0.execute.mem_stage_pc\[0\] _2386_ _2387_ _2388_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7398_ _1338_ _3317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8058__A2 _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9137_ _0149_ clknet_leaf_115_i_clk core_0.execute.alu_mul_div.div_cur\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6349_ _2144_ _2324_ _2325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_227_3235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6069__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7805__A2 _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9068_ _0093_ clknet_leaf_100_i_clk core_0.decode.i_instr_l\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5816__A1 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8019_ core_0.execute.rf.reg_outputs\[4\]\[14\] _3693_ _3704_ _3712_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_216_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8644__C _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7569__A1 _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_3364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_7_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7741__A1 _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7790__I _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8049__A2 _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8835__B _4326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_180_2670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5035__A2 _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6783__A2 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7980__A1 core_0.execute.rf.reg_outputs\[5\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5720_ core_0.execute.sreg_priv_control.o_d\[8\] _1701_ _1717_ _1698_ _1718_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_174_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4794__A1 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__B1 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4794__B2 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7186__B _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5651_ net37 _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_150_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_216_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6535__A2 _2370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7732__A1 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4602_ core_0.execute.rf.reg_outputs\[7\]\[8\] net297 _0697_ core_0.execute.rf.reg_outputs\[3\]\[8\]
+ _0793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_182_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8370_ _1544_ _3982_ _3983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5582_ _1069_ core_0.fetch.submitable _1622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_72_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7321_ _2549_ _3241_ _3242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_53_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4533_ _0729_ net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_53_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7914__B _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_211_3047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6299__A1 _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8729__C _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7252_ _2536_ _3173_ _3174_ _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_229_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4464_ core_0.dec_r_reg_sel\[2\] _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_123_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6838__A3 _2692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4849__A2 _1023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_229_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5434__B _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6203_ _2169_ _2191_ _2192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7183_ _1337_ _2355_ _1285_ _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_55_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ core_0.execute.alu_mul_div.i_mul _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_225_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_209_Left_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_225_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8460__A2 _2136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6065_ _1757_ _2054_ _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_213_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6471__A1 core_0.execute.trap_flag vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5274__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5016_ _1185_ _1165_ _1187_ _1190_ _1080_ net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_23_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_1_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_222_3176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_178_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8212__A2 _3836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer72_I _0664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5026__A2 _1149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6967_ _2833_ _2881_ _2896_ _2897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6774__A2 _2706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7971__A1 core_0.execute.rf.reg_outputs\[5\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8706_ net196 _0900_ _4266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4785__A1 _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5918_ core_0.execute.rf.reg_outputs\[4\]\[9\] _1776_ _1804_ core_0.execute.rf.reg_outputs\[11\]\[9\]
+ _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_194_2839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6898_ net79 _2829_ _1401_ _2830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_218_Left_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8637_ _2675_ _4202_ _4208_ _1501_ _0562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5609__B _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5849_ net190 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_29_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8568_ _4080_ _3335_ _4147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_210_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7519_ _3401_ _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7824__B _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output186_I net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8499_ _4041_ _4085_ _4086_ _4087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7115__I _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_227_Left_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_219_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5063__C _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_86_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8451__A2 _4042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6462__A1 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8203__A2 _3821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7411__B1 _3311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6765__A2 _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7962__A1 _3427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_2403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_236_Left_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_2414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5973__B1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7714__A1 _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4528__B2 core_0.execute.rf.reg_outputs\[12\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7734__B _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_1627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_245_Left_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4649__I net251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_2543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__B2 core_0.execute.rf.reg_outputs\[12\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8978__B1 _1470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_219_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8442__A2 _4031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7870_ core_0.execute.rf.reg_outputs\[8\]\[15\] _3605_ _3621_ _3626_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5008__A2 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6821_ _1326_ _2747_ _2750_ _2753_ _2754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_77_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7909__B _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7953__A1 core_0.execute.rf.reg_outputs\[5\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7695__I _3519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6756__A2 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9540_ _0550_ clknet_leaf_81_i_clk net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_202_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4767__A1 core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ _2681_ _2682_ _2684_ _2685_ _2686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_174_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5703_ _1608_ _1706_ _0130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9471_ _0481_ clknet_leaf_48_i_clk core_0.execute.rf.reg_outputs\[1\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6683_ _2146_ _2614_ net210 _2624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_174_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6508__A2 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8422_ _2230_ _4025_ _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5634_ core_0.decode.i_imm_pass\[11\] _1645_ _1653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8353_ _3945_ _3947_ _3959_ _3961_ _3967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_60_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5192__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5565_ _1608_ _1612_ _0086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_170_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7304_ _2703_ _3225_ _3226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4516_ _0713_ net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_8284_ _1668_ _2054_ _3902_ _3903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5496_ net44 _1554_ _1575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8130__A1 core_0.execute.rf.reg_outputs\[1\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7235_ _3157_ _3158_ _3159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4559__I _0753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8681__A2 _4209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_108_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5495__A2 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7166_ _3051_ _3086_ _3091_ _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_224_3205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6117_ core_0.execute.rf.reg_outputs\[7\]\[1\] _1821_ _1799_ core_0.execute.rf.reg_outputs\[6\]\[1\]
+ _2107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_95_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8433__A2 _4032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _1337_ _2360_ core_0.decode.oc_alu_mode\[7\] _3024_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_225_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6048_ _2030_ _2032_ _2037_ _2038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_142_2215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_206_2982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8197__A1 _1670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7944__A1 core_0.execute.rf.reg_outputs\[6\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7999_ _3427_ _3694_ _3701_ _0431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6747__A2 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output101_I net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4758__A1 core_0.ew_reg_ie\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4758__B2 core_0.ew_reg_ie\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5955__B1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_235_3334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4930__A1 core_0.fetch.prev_request_pc\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4469__I _0666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8672__A2 _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6683__A1 _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5486__A2 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8385__B _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4694__B1 net341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_244_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_188_Right_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6435__A1 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8975__A3 _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_2484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8188__A1 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9311__CLK clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7729__B _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7935__A1 _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__B1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6352__C _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7163__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4921__A1 core_0.fetch.prev_request_pc\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5350_ core_0.dec_rf_ie\[6\] _1438_ _1462_ _1466_ _1467_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xoutput205 net279 sr_bus_data_o[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8112__A1 _3427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_239_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6123__B1 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5281_ _1401_ _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_227_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7020_ _2759_ _2934_ _2945_ _2948_ _2949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_52_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_155_Right_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_156_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5431__C _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8971_ _1465_ _1230_ _1272_ _4453_ _0651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4988__A1 _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7922_ _3650_ _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_172_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8179__A1 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7639__B _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7853_ core_0.execute.rf.reg_outputs\[8\]\[7\] _3613_ _3609_ _3617_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7926__A1 _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6804_ _1899_ _2090_ _2737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_148_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7784_ core_0.execute.rf.reg_outputs\[10\]\[10\] _3570_ _3568_ _3577_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4996_ _1165_ _1173_ _1174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_46_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5159__B _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6735_ _2662_ _2668_ _2665_ _2670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_191_2809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9523_ _0533_ clknet_leaf_117_i_clk core_0.execute.alu_mul_div.div_res\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_190_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9454_ _0464_ clknet_leaf_23_i_clk core_0.execute.rf.reg_outputs\[2\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6666_ _0943_ _0957_ _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_190_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8351__A1 _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7154__A2 _3079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer35_I _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__I _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8405_ _2221_ _4013_ core_0.execute.alu_mul_div.div_res\[0\] _4014_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5165__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ core_0.decode.i_imm_pass\[3\] _1616_ _1644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9385_ _0395_ clknet_4_3__leaf_i_clk core_0.execute.rf.reg_outputs\[6\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5673__I _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6597_ _2465_ _2535_ _2539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6901__A2 _2785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8189__C _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_230_3275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4912__A1 core_0.fetch.prev_request_pc\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8336_ _1542_ _1942_ _3951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5548_ _1597_ _1603_ _0078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8103__A1 _3401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_3_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input62_I i_req_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8267_ _3875_ _3887_ _3888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5479_ _1564_ _0048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8654__A2 _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7218_ _2564_ _2814_ _3141_ _3142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_8198_ _1535_ core_0.execute.alu_mul_div.cbit\[2\] _3824_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4676__B1 _0683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7149_ _1337_ _2461_ _3070_ _1885_ _3074_ _3075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_214_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9334__CLK clknet_leaf_155_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_122_Right_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_232_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_214_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_225_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6968__A2 _2881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7090__A1 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__A1 _1023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8652__C _4201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7917__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5928__B1 _1778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7268__C core_0.execute.alu_mul_div.i_mod vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8590__A1 _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4600__B1 _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8342__A1 _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8893__A2 _4385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6105__B1 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5459__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6656__A1 _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_2502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_217_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6408__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7456__I0 net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8843__B _4326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6959__A2 _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7081__A1 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5631__A2 _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8956__I0 net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4662__I _0848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4850_ net49 core_0.fetch.out_buffer_data_instr\[20\] _1017_ _1031_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_2631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7384__A2 _3303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_2642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8581__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6041__C1 _1787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A1 _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4781_ core_0.dec_l_reg_sel\[3\] _0943_ _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_142_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6520_ _1846_ net213 _2462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_27_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7136__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8333__B2 _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7194__B core_0.execute.alu_mul_div.i_mod vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6451_ _1175_ _2386_ _2408_ _0176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5147__A1 _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8884__A2 _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5698__A2 _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_1699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5402_ _1451_ _1504_ _1505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9170_ _0181_ clknet_leaf_42_i_clk core_0.execute.prev_pc_high\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_224_Right_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6382_ _1668_ _1942_ _2356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8121_ _3647_ _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5333_ _1243_ _1295_ _1316_ _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_208_3008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_2771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8052_ _3459_ _3716_ _3731_ _0454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_121_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5264_ core_0.dec_jump_cond_code\[2\] _1379_ _1382_ _1384_ _1381_ _1377_ _1385_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai222_4
XTAP_TAPCELL_ROW_110_1833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7003_ _2841_ _2931_ _2570_ _2932_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_227_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _1236_ _1256_ _1273_ _1339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5870__A2 net254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8954_ net192 core_0.decode.i_imm_pass\[9\] _1264_ _4445_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_222_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5622__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_203_2952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7905_ core_0.execute.rf.reg_outputs\[7\]\[14\] _3627_ _3636_ _3646_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6273__B _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8885_ core_0.execute.pc_high_buff_out\[4\] _4385_ _1430_ _4402_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4572__I _0765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_159_Left_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_176_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7836_ _3605_ _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_219_3137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8572__A1 _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7375__A2 core_0.execute.alu_mul_div.mul_res\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_1962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4979_ _1023_ _1158_ _1159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7883__I _3627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7767_ _3415_ _3563_ _3567_ _0333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_175_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9506_ _0516_ clknet_leaf_122_i_clk core_0.execute.alu_mul_div.mul_res\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6718_ _2648_ _2647_ _2646_ _2655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7127__A2 net277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7698_ _3512_ _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_137_2158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5138__A1 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9437_ _0447_ clknet_leaf_49_i_clk core_0.execute.rf.reg_outputs\[3\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6649_ _1912_ _1943_ _1329_ _2591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_144_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8875__A2 _4383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_2314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5689__A2 core_0.execute.sreg_priv_control.o_d\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6886__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9368_ _0378_ clknet_leaf_151_i_clk core_0.execute.rf.reg_outputs\[8\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7832__B _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_168_Left_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_8319_ _3927_ _3935_ _3936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8627__A2 _1696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9299_ _0309_ clknet_leaf_8_i_clk core_0.execute.rf.reg_outputs\[12\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__B _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_243_3433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8663__B _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7063__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_2443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6810__A1 _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5613__A2 _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_177_Left_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_243_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4482__I _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8563__A1 _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8563__B2 _2134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5377__B2 _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7118__A2 _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_2572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5019__S _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6877__A1 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_186_Left_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7742__B _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8618__A2 _2761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6358__B _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5301__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5852__A2 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_195_Left_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6801__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5951_ net88 _1813_ _1933_ _1940_ _1941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_149_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__A4 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4902_ _0891_ _1082_ _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_8670_ core_0.execute.sreg_irq_pc.o_d\[6\] _4210_ _4236_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_153_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5882_ net87 _0667_ _1872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8554__A1 _4133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4833_ _0894_ _1012_ _1013_ _1014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8799__I _4324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5368__A1 _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7621_ _3428_ _3476_ _3483_ _0271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7552_ _3397_ _3428_ _3430_ _0255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_173_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4764_ _0944_ _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__8306__A1 _1925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7109__A2 core_0.execute.alu_mul_div.mul_res\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6503_ _1753_ _2341_ _2445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_145_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5437__B _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7483_ core_0.dec_rf_ie\[10\] core_0.ew_reg_ie\[10\] _3366_ _3375_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4591__A2 _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4695_ _0667_ _0876_ _0877_ _0878_ _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_71_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_3078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6868__A1 _1309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6434_ core_0.execute.mem_stage_pc\[6\] _2395_ _2387_ _2398_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9222_ _0233_ clknet_leaf_138_i_clk core_0.ew_reg_ie\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__6868__B2 _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9153_ _0164_ clknet_leaf_67_i_clk core_0.execute.mem_stage_pc\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5540__A1 _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ _2105_ _2106_ _2107_ _2108_ _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4995__C _1026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8104_ core_0.execute.rf.reg_outputs\[1\]\[1\] _3760_ _3756_ _3762_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5316_ _1434_ net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7371__C _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9084_ _0109_ clknet_leaf_93_i_clk core_0.decode.i_imm_pass\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6296_ _2185_ _2256_ _2278_ _2229_ _0151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8035_ _3714_ _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7293__A1 _1254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6096__A2 _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__B2 _3069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _1369_ core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_194_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5843__A2 net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5178_ _1326_ _1286_ _1327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input25_I i_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_196_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8937_ _1868_ _0038_ _4436_ _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_27_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8868_ net193 _4387_ _4388_ _4389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7348__A2 _3268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8545__A1 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5359__A1 _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7819_ _3451_ _3585_ _3597_ _0355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8799_ _4324_ _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_108_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8848__A2 _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output93_I net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8658__B _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__I _0664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6087__A2 _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5834__A2 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7036__A1 _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7587__A2 core_0.ew_data\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5101__I core_0.decode.i_instr_l\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8536__A1 _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7339__A2 _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_2601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A2 _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5770__A1 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A2 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4480_ net301 core_0.dec_r_reg_sel\[1\] _0678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_80_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_144_i_clk clknet_4_1__leaf_i_clk clknet_leaf_144_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_96_1669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xmax_cap226 _1780_ net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7511__A2 _3388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5522__A1 net58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6150_ core_0.execute.alu_mul_div.cbit\[2\] _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_148_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_185_2730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7275__A1 _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5101_ core_0.decode.i_instr_l\[1\] _1257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_237_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6081_ _2055_ _2070_ _2071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5032_ _1106_ _1149_ _1203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7698__I _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7578__A2 _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8775__A1 core_0.execute.sreg_scratch.o_d\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5589__A1 _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _1337_ _2492_ core_0.decode.oc_alu_mode\[7\] _2913_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_164_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_200_2911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8722_ _4224_ _4150_ _4278_ _1662_ _4279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_87_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ _1916_ _1923_ _1924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8527__A1 _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_105_1776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_216_3107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8653_ _2822_ _4202_ _4222_ _1501_ _0564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5865_ net314 net198 _1854_ _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_196_2870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6002__A2 net322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7604_ _3387_ core_0.ew_data\[15\] _3449_ net27 _3472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_29_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4816_ core_0.execute.alu_mul_div.i_mod _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_8_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8584_ _2816_ _2868_ _4159_ _4161_ _4162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_90_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5796_ _0971_ _0943_ net328 _0958_ _1786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_173_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7750__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7535_ core_0.execute.rf.reg_outputs\[15\]\[2\] _3403_ _2404_ _3416_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4747_ _0668_ net301 _0928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5761__A1 _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7466_ _2418_ _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4678_ core_0.execute.rf.reg_outputs\[5\]\[2\] _0677_ net347 core_0.execute.rf.reg_outputs\[15\]\[2\]
+ _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7502__A2 _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8478__B _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9205_ _0216_ clknet_leaf_52_i_clk core_0.ew_addr\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6417_ _1430_ _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_3_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7397_ net212 _1974_ _3316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5681__I net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9136_ _0148_ clknet_leaf_115_i_clk core_0.execute.alu_mul_div.div_cur\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6348_ _2149_ _2317_ _2323_ _2324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_227_3236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9067_ _0092_ clknet_leaf_110_i_clk core_0.decode.i_instr_l\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6279_ _2246_ _2262_ _2263_ _2217_ _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_228_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_216_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5816__A2 _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8018_ _3465_ _3695_ _3711_ _0440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_145_2257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8518__A1 _4080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_3365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_82_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7741__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_61_i_clk clknet_4_9__leaf_i_clk clknet_leaf_61_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4555__A2 _0683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_2386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76_i_clk clknet_4_11__leaf_i_clk clknet_leaf_76_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_207_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7009__A1 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8206__B1 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8757__A1 core_0.execute.sreg_scratch.o_d\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9568__CLK clknet_leaf_21_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_180_2671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8851__B _4326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_14_i_clk clknet_4_3__leaf_i_clk clknet_leaf_14_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_187_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8509__A1 _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7980__A2 _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__A1 core_0.execute.rf.reg_outputs\[1\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4794__A2 _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5650_ _1660_ _0123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7732__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4601_ core_0.execute.rf.reg_outputs\[4\]\[8\] _0719_ net316 core_0.execute.rf.reg_outputs\[8\]\[8\]
+ _0792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_29_i_clk clknet_4_8__leaf_i_clk clknet_leaf_29_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_170_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5581_ _1139_ _1615_ _1621_ _0093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5743__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7320_ _2552_ _3240_ _3241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_170_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ _0714_ _0716_ _0723_ _0728_ _0729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_211_3048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7251_ _2536_ _3173_ core_0.decode.oc_alu_mode\[11\] _3174_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4463_ _0660_ _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_111_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ _2184_ _2189_ _2190_ _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_159_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4849__A3 _1026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7182_ _3060_ _2758_ _3106_ _3063_ _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XPHY_EDGE_ROW_15_Right_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5434__C _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6133_ _1867_ _1893_ _2122_ _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_55_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ net100 _1771_ _2046_ _2053_ _2054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_5015_ _1189_ _1146_ _1164_ _1190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_175_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6471__A2 _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8748__A1 core_0.execute.sreg_scratch.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_222_3177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7420__A1 net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7420__B2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_24_Right_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6966_ _1401_ _2894_ _2895_ _2896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7971__A2 _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8705_ core_0.execute.sreg_irq_pc.o_d\[12\] _4209_ _4265_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_191_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_132_Left_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_140_2198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ core_0.execute.rf.reg_outputs\[15\]\[9\] _0945_ _1794_ core_0.execute.rf.reg_outputs\[8\]\[9\]
+ _1907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_104_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5982__A1 _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4785__A2 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6897_ _2673_ _1411_ _2829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_75_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8636_ _1662_ core_0.execute.mem_stage_pc\[0\] _4201_ _4207_ _4208_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5848_ _1831_ _1833_ _1835_ _1837_ _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_91_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8920__A1 _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4537__A2 _0680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5734__A1 _1726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8567_ _4053_ _4145_ _4146_ _1702_ _0554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_161_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5779_ _1328_ _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XTAP_TAPCELL_ROW_118_1923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7518_ _3382_ core_0.ew_data\[0\] _3400_ _3401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_8498_ net83 _4040_ _4086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output179_I net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7449_ _2616_ _3120_ _3357_ _0225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_169_Right_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_141_Left_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_229_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7239__A1 _3156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7840__B _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4956__S _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9119_ _0131_ clknet_leaf_109_i_clk core_0.execute.sreg_long_ptr_en vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_228_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8987__A1 _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_29_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6462__A2 _0904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4473__A1 _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7411__A1 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7411__B2 _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_150_Left_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7962__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_2404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A1 core_0.execute.rf.reg_outputs\[8\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__B2 core_0.execute.rf.reg_outputs\[4\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7714__A2 _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8911__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4528__A2 net341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5725__A1 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_51_Right_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_140_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__B _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_136_Right_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_2544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__A2 net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_2700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8978__B2 _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_60_Right_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_179_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7402__A1 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6205__A2 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6820_ _1309_ _2445_ _2751_ _2076_ _2752_ _2753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_159_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7953__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6756__A3 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4767__A2 core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6751_ core_0.execute.sreg_scratch.o_d\[0\] _1686_ net227 _2683_ _2685_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_102_1735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ core_0.execute.sreg_data_page _1701_ _1705_ _1698_ _1706_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_161_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9470_ _0480_ clknet_leaf_48_i_clk core_0.execute.rf.reg_outputs\[1\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6682_ _2621_ _2622_ _2623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7705__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7925__B _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8421_ _4015_ _4024_ core_0.execute.alu_mul_div.div_res\[5\] _4025_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5633_ _1037_ _1628_ _1652_ _0114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5564_ core_0.fetch.prev_request_pc\[14\] _1082_ _1083_ net165 _1612_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8352_ core_0.execute.alu_mul_div.mul_res\[12\] _3966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4515_ net93 _0667_ _0691_ _0712_ _0713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_7303_ _1317_ _3223_ _3224_ _3225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_8283_ _1668_ _2487_ _3902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5495_ _1573_ _1551_ _1574_ _0054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8130__A2 _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_103_Right_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7234_ core_0.execute.sreg_irq_pc.o_d\[10\] _3042_ _3044_ core_0.execute.sreg_scratch.o_d\[10\]
+ _3158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_186_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_1864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7660__B _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7165_ _3087_ _3090_ _1403_ _3091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_95_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_224_3206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8969__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_30_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6116_ core_0.execute.rf.reg_outputs\[1\]\[1\] _1779_ _1794_ core_0.execute.rf.reg_outputs\[8\]\[1\]
+ _2106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7096_ _1309_ _2429_ _3023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_226_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6444__A2 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7641__A1 core_0.execute.rf.reg_outputs\[14\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6047_ _2033_ _2034_ _2035_ _2036_ _2037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_213_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_2216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_206_2983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7886__I _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8197__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9113__CLK clknet_leaf_110_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7998_ core_0.execute.rf.reg_outputs\[4\]\[4\] _3700_ _3689_ _3701_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6747__A3 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4758__A2 _0928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4524__B _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6949_ _2694_ net80 _2879_ _1403_ _2880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_64_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_238_Right_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_235_3335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8619_ _2816_ _2868_ _4192_ _4193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_107_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5707__A1 _0848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9599_ _0609_ clknet_leaf_61_i_clk core_0.execute.pc_high_out\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4930__A2 _1060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6132__A1 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8666__B _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6683__A2 _2614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7880__A1 _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4694__B2 core_0.execute.rf.reg_outputs\[3\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4485__I net297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6435__A2 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7632__A1 _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7483__I1 core_0.ew_reg_ie\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_2485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4997__A2 _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8188__A2 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7935__A2 _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4749__A2 _0675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5946__A1 core_0.execute.rf.reg_outputs\[5\]\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_205_Right_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7148__B1 _1925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7745__B _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7699__A1 core_0.execute.rf.reg_outputs\[12\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5174__A2 _1322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput206 net268 sr_bus_data_o[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4921__A2 _1023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8112__A2 _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6123__A1 core_0.execute.rf.reg_outputs\[13\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5280_ core_0.dec_sreg_irt _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_49_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7871__A1 _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4685__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4685__B2 _0869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7623__A1 _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8970_ core_0.dec_jump_cond_code\[1\] _1250_ _4453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7921_ _3421_ _3651_ _3656_ _0398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8179__A2 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7852_ _3441_ _3606_ _3616_ _0369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5237__I0 core_0.ew_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7926__A2 _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6803_ _1751_ _1898_ _2735_ _2736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_187_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5937__A1 _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7783_ _3454_ _3563_ _3576_ _0340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4995_ _1133_ _1141_ _1144_ _1026_ _1173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_175_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9522_ _0532_ clknet_leaf_118_i_clk core_0.execute.alu_mul_div.div_res\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6734_ _2662_ _2665_ _2668_ _2669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_63_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7655__B _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9453_ _0463_ clknet_leaf_23_i_clk core_0.execute.rf.reg_outputs\[2\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6665_ net315 net211 _2607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_6_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8404_ _2246_ _2216_ _4013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5616_ _1063_ _1615_ _1643_ _0106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9384_ _0394_ clknet_leaf_154_i_clk core_0.execute.rf.reg_outputs\[7\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5165__A2 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer28_I net254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ net311 _2531_ _2534_ _2537_ _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_83_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8335_ _3832_ _3949_ _3950_ _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5547_ core_0.fetch.prev_request_pc\[6\] _1595_ _1084_ net172 _1603_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_230_3276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4912__A2 _1057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8103__A2 _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5478_ core_0.fetch.out_buffer_data_instr\[8\] net67 _1559_ _1564_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8266_ _1535_ _3886_ _3887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8486__B _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input55_I i_req_data[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7217_ _2568_ _3139_ _3140_ _2563_ _3141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_111_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6665__A2 net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8197_ _1670_ _1812_ _3823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4676__B2 core_0.execute.rf.reg_outputs\[7\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7148_ _3071_ net306 _1925_ _3072_ _3073_ _3074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_226_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7614__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7079_ _2711_ _2994_ _3006_ _3007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_226_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4979__A2 _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6734__B _2668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7378__B1 _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7917__A2 _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5928__B2 core_0.execute.rf.reg_outputs\[1\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4600__A1 core_0.execute.rf.reg_outputs\[5\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7565__B _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8240__I core_0.execute.alu_mul_div.mul_res\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6353__A1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6105__A1 core_0.execute.rf.reg_outputs\[3\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7853__A1 core_0.execute.rf.reg_outputs\[8\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_2503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7456__I1 _3261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8030__A1 _3408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_177_2632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__B1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8581__A2 _2770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6041__C2 core_0.execute.rf.reg_outputs\[3\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4780_ core_0.ew_reg_ie\[10\] _0956_ _0959_ core_0.ew_reg_ie\[11\] _0960_ core_0.ew_reg_ie\[8\]
+ _0961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_172_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8333__A2 _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6450_ core_0.execute.mem_stage_pc\[12\] _2395_ _2404_ _2408_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5401_ _1502_ _1503_ _1504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6381_ net213 _2355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_140_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8120_ _3450_ _3759_ _3770_ _0483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _1241_ _1305_ _1306_ _1449_ _1450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_140_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5263_ core_0.dec_jump_cond_code\[2\] _1383_ _1384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8051_ core_0.execute.rf.reg_outputs\[3\]\[11\] _3722_ _3730_ _3731_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_208_3009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_2772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4658__A1 core_0.execute.rf.reg_outputs\[3\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7002_ net267 _2930_ _2931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_110_1834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5194_ _1337_ _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_208_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8753__C _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8953_ _1688_ _0038_ _4444_ _0642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_222_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4853__I _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7904_ _3466_ _3629_ _3645_ _0392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8884_ net203 _4387_ _4400_ _4401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_203_2953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8021__A1 core_0.execute.rf.reg_outputs\[4\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7835_ _3605_ _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_219_3138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6032__B1 _1818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6583__A1 _2428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7766_ core_0.execute.rf.reg_outputs\[10\]\[2\] _3564_ _3554_ _3567_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_121_1963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4978_ _1145_ _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_18_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9505_ _0515_ clknet_leaf_119_i_clk core_0.execute.alu_mul_div.mul_res\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6717_ _2652_ _2653_ _2654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_117_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7697_ _3428_ _3520_ _3527_ _0303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9436_ _0446_ clknet_leaf_61_i_clk core_0.execute.rf.reg_outputs\[3\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6648_ _1769_ _2589_ net270 _2590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5138__A2 _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6335__A1 _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_2315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5689__A3 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6886__A2 _2816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9367_ _0377_ clknet_leaf_151_i_clk core_0.execute.rf.reg_outputs\[8\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6579_ _2520_ _1962_ _1916_ _1923_ _2521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__4897__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8318_ _3934_ _3935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9298_ _0308_ clknet_leaf_27_i_clk core_0.execute.rf.reg_outputs\[12\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output161_I net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8249_ _3865_ _3870_ _3871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_218_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_243_3423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_243_3434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9451__CLK clknet_leaf_136_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_2444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6810__A2 _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8012__A1 _3456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_wire210_I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5377__A2 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6574__A1 _2439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_152_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5594__I _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5129__A2 _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6326__A1 _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_2573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8079__A1 _3440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7826__A1 core_0.execute.rf.reg_outputs\[9\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5301__A2 net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_77_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_232_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6801__A2 _2733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8145__I _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5950_ _1772_ _1934_ _1939_ _1940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_220_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8003__A1 _3440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4901_ _1078_ _1081_ _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_47_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ _0667_ _0886_ _0887_ _0888_ _1871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_239_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7620_ core_0.execute.rf.reg_outputs\[14\]\[4\] _3482_ _3467_ _3483_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4832_ _0894_ net48 _1013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6565__A1 _2008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4576__B1 _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7551_ core_0.execute.rf.reg_outputs\[15\]\[4\] _3429_ _3422_ _3430_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_60_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4763_ _0942_ _0943_ core_0.dec_l_reg_sel\[1\] core_0.dec_l_reg_sel\[0\] _0944_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_0_117_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8306__A2 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6502_ _2008_ _2102_ _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_43_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6317__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7482_ _3374_ _0241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4694_ core_0.execute.rf.reg_outputs\[11\]\[1\] net303 net341 core_0.execute.rf.reg_outputs\[3\]\[1\]
+ _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__9324__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_3079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9221_ _0232_ clknet_leaf_138_i_clk core_0.ew_reg_ie\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_126_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6433_ _1206_ _2385_ _2397_ _0169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4879__A1 _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9152_ _0014_ clknet_leaf_44_i_clk net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6364_ net94 _2338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8103_ _3401_ _3759_ _3761_ _0475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7817__A1 _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5315_ _1419_ core_0.execute.sreg_priv_control.o_d\[0\] _1433_ _1434_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__9474__CLK clknet_leaf_16_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6295_ core_0.execute.alu_mul_div.div_cur\[6\] _2246_ _2276_ _2277_ _2256_ _2278_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_9083_ _0108_ clknet_leaf_93_i_clk core_0.decode.i_imm_pass\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8490__A1 _1738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8034_ _3420_ _3715_ _3721_ _0446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6096__A3 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5246_ _1368_ _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_194_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_89_Right_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_243_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5177_ core_0.decode.oc_alu_mode\[11\] _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_rebuffer95_I _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8242__A1 core_0.execute.alu_mul_div.mul_res\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5056__A1 core_0.fetch.prev_request_pc\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5679__I _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I i_irq vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8936_ core_0.decode.i_imm_pass\[0\] _1293_ _4436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4803__A1 _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8867_ _0908_ _4387_ _4388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6005__B1 _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7818_ core_0.execute.rf.reg_outputs\[9\]\[8\] _3591_ _3595_ _3597_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6556__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8798_ _4326_ _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_47_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_98_Right_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_163_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4567__B1 _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7749_ core_0.execute.rf.reg_outputs\[11\]\[11\] _3548_ _3554_ _3557_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6308__A1 _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9419_ _0429_ clknet_leaf_136_i_clk core_0.execute.rf.reg_outputs\[4\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output86_I net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_18_Left_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_219_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5819__B1 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8481__A1 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7036__A2 _2954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8233__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5047__A1 core_0.fetch.prev_request_pc\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6795__A1 _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_27_Left_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6547__A1 _2439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_174_2602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__A2 _1753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7753__B _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap216 _0870_ net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_96_1659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_150_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5522__A2 _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_2731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5100_ _1255_ _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_20_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6080_ _1874_ net214 _2070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8472__A1 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_9__f_i_clk_I clknet_3_4_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7979__I _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__A1 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5031_ net83 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_189_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_224_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7027__A2 _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8224__A1 _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5038__A1 core_0.fetch.prev_request_pc\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8775__A2 _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Left_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5589__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6786__A1 _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6982_ net325 _2909_ _2911_ _2912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_200_2912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8721_ net77 _1740_ _1732_ _4205_ _4278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_220_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5933_ _1917_ _1918_ _1919_ _1922_ _1923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_76_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8652_ _1662_ core_0.execute.mem_stage_pc\[2\] _4220_ _4221_ _4201_ _4222_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_196_2860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5864_ _1518_ net182 _1854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_216_3108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_185_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7603_ _3403_ _3470_ _3471_ _0265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4549__B1 _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4815_ core_0.execute.alu_mul_div.i_div _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_91_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8583_ _4160_ _2761_ _4161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5795_ _1784_ _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_146_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7534_ _3414_ _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4746_ core_0.execute.next_ready_delayed _0927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_161_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5761__A2 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7465_ _3365_ _0233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_160_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4677_ core_0.execute.rf.reg_outputs\[1\]\[2\] net302 net321 core_0.execute.rf.reg_outputs\[12\]\[2\]
+ _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_9204_ _0215_ clknet_leaf_78_i_clk core_0.ew_data\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_114_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6416_ _1433_ _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5513__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7396_ _3020_ _3069_ _3315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_9135_ _0147_ clknet_leaf_116_i_clk core_0.execute.alu_mul_div.div_cur\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_101_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6347_ _2148_ _2323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_228_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_100_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_227_3237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8463__A1 _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7266__A2 _3188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9066_ _0091_ clknet_leaf_110_i_clk core_0.decode.i_instr_l\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6278_ core_0.execute.alu_mul_div.div_cur\[4\] _2224_ _2263_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8017_ core_0.execute.rf.reg_outputs\[4\]\[13\] _3700_ _3704_ _3711_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5229_ core_0.ew_data\[2\] core_0.ew_data\[10\] _1349_ _1360_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5816__A3 _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8215__A1 _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5029__A1 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output124_I net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6777__A1 core_0.dec_sreg_load vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8919_ _1488_ _1510_ _4423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_196_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8518__A2 _3085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6529__A1 net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_238_3366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_25_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5201__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_117_Right_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_156_2387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4488__I _0685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7799__I _3584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5268__A1 core_0.execute.alu_flag_reg.o_d\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__S _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8206__B2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8757__A2 _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_2672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6768__A1 _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5112__I _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5976__C1 _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8509__A2 core_0.execute.sreg_irq_pc.o_d\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5991__A2 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ core_0.execute.rf.reg_outputs\[5\]\[8\] net222 _0679_ core_0.execute.rf.reg_outputs\[11\]\[8\]
+ _0791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_182_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5580_ core_0.decode.i_instr_l\[4\] _1616_ _1621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _0724_ _0725_ _0726_ _0727_ _0728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4900__B _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5782__I _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_211_3049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8693__A1 _4219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7250_ _3136_ _2540_ _3173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
X_4462_ core_0.dec_r_reg_sel\[3\] _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_7_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6201_ core_0.execute.alu_mul_div.div_cur\[5\] _1851_ _2190_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4703__B1 net341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__A4 _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7181_ _2587_ _3104_ _3105_ _3060_ _3106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_111_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6132_ _1894_ _2004_ _2121_ _2122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8445__A1 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6063_ _2047_ _2048_ _2049_ _2052_ _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5014_ _0895_ _1035_ _1188_ _1189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_53_Left_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_225_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_219_Right_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_240_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8748__A2 _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_222_3178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6759__A1 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7420__A2 _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7658__B _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6965_ _1401_ core_0.execute.sreg_irq_pc.o_d\[4\] _2895_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_220_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5431__A1 _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8704_ _4263_ _4264_ _1435_ _0573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5916_ core_0.execute.rf.reg_outputs\[3\]\[9\] _1788_ _1819_ core_0.execute.rf.reg_outputs\[12\]\[9\]
+ _1906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_140_2188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clone30_I _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6896_ _2694_ _2827_ _2828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_193_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8635_ _4203_ _1226_ _4206_ _1661_ _4207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_192_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7184__A1 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ net313 net197 _1836_ _1837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_8_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8566_ net76 _4052_ _4146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5778_ _1763_ _1767_ _1768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__6931__A1 _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5734__A2 _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7517_ _3382_ _3398_ _3399_ _3400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_118_1924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4729_ core_0.execute.pc_high_out\[7\] _0901_ _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8497_ net83 _4084_ _4085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_31_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7448_ net129 _2419_ _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8684__A1 _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__A1 net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7379_ core_0.execute.sreg_priv_control.o_d\[14\] _1693_ _2996_ net6 _2689_ _3299_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_102_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9118_ _0130_ clknet_leaf_64_i_clk core_0.execute.sreg_data_page vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_229_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9049_ _0075_ clknet_leaf_85_i_clk core_0.fetch.prev_request_pc\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_216_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6998__A1 core_0.ew_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__A2 _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_143_i_clk clknet_4_1__leaf_i_clk clknet_leaf_143_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5958__C1 _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_2405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_15__f_i_clk_I clknet_3_7_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A2 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6922__A1 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__A2 _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_180_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8675__A1 _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__I _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_2545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8427__A1 _3038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_2701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8978__A2 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6989__A1 core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5110__B1 _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8354__S _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7402__A2 _2556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5413__A1 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6756__A4 _2687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7197__C _2689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ net105 _1405_ net227 _2683_ _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_57_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_147_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_102_1736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5701_ net215 _1704_ _1705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_221_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6681_ _2614_ _2620_ _2622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_193_2830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8420_ _1540_ _1543_ _3878_ _4024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__8902__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5632_ core_0.decode.i_imm_pass\[10\] _1645_ _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_rebuffer8_I net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5716__A2 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4924__B1 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8351_ _3832_ _3964_ _3965_ _0519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5563_ _1608_ _1611_ _0085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8102__B _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7302_ core_0.execute.alu_mul_div.div_cur\[12\] _2128_ _3224_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8666__A1 net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4514_ _0696_ _0701_ _0706_ _0711_ _0712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_5_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8282_ _3893_ _3895_ _3900_ _3901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_14_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5494_ net43 _1554_ _1574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6677__B1 _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7233_ core_0.execute.sreg_priv_control.o_d\[10\] _1693_ _2996_ net2 _3157_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8756__C _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7164_ _3088_ _3089_ _2673_ _3090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8969__A2 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6115_ core_0.execute.rf.reg_outputs\[12\]\[1\] _1819_ _1962_ _2105_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_225_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7095_ _2006_ _3019_ _3021_ _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7641__A2 _3475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6046_ core_0.execute.rf.reg_outputs\[2\]\[5\] net336 net226 core_0.execute.rf.reg_outputs\[10\]\[5\]
+ _2036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_241_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_60_i_clk clknet_4_11__leaf_i_clk clknet_leaf_60_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_142_2217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_206_2984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7997_ _3693_ _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5404__A1 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6747__A4 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6948_ _2875_ _2876_ _2877_ _2878_ _2879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_48_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5955__A2 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_75_i_clk clknet_4_11__leaf_i_clk clknet_leaf_75_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_235_3336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9408__CLK clknet_leaf_37_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6879_ _1894_ _2804_ _2809_ _2810_ _2811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_165_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8618_ _2123_ _2761_ _4191_ _4192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_107_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6904__A1 _2708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9598_ _0608_ clknet_leaf_61_i_clk core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_64_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5707__A2 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output191_I net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4915__B1 _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8549_ _4130_ _4131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8657__A1 _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8947__B _4441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6668__B1 _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7851__B _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8666__C _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_13_i_clk clknet_4_3__leaf_i_clk clknet_leaf_13_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7880__A2 _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4694__A2 net303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__A1 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4766__I core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7632__A2 _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8682__B _1717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_28_i_clk clknet_4_8__leaf_i_clk clknet_leaf_28_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5643__A1 _1023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_2475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_164_2486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__A2 _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7148__B2 _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8896__A1 net277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7699__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6371__A2 _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8648__A1 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput207 net207 sr_bus_data_o[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6123__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7871__A2 _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5882__A1 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8820__A1 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7623__A2 _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8592__B _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7920_ core_0.execute.rf.reg_outputs\[6\]\[3\] _3652_ _3648_ _3656_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_222_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7851_ core_0.execute.rf.reg_outputs\[8\]\[6\] _3613_ _3609_ _3616_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7387__A1 _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__I1 core_0.ew_data\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6802_ _1896_ _2731_ _2734_ _2735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7782_ core_0.execute.rf.reg_outputs\[10\]\[9\] _3570_ _3568_ _3576_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4994_ _1158_ _1155_ _1171_ _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_58_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9521_ _0531_ clknet_leaf_120_i_clk core_0.execute.alu_mul_div.div_res\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6733_ _2666_ _2667_ _2668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7936__B _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_147_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7428__S _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9452_ _0462_ clknet_leaf_16_i_clk core_0.execute.rf.reg_outputs\[2\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8887__A1 _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6664_ _2479_ _2481_ _2560_ _1326_ _2605_ _2606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_45_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8403_ _2413_ _1004_ _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_155_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5615_ core_0.decode.i_imm_pass\[2\] _1616_ _1643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9383_ _0393_ clknet_leaf_154_i_clk core_0.execute.rf.reg_outputs\[7\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6595_ _2536_ _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5165__A3 _1313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8334_ core_0.execute.alu_mul_div.mul_res\[10\] _3830_ _3950_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5546_ _1597_ _1602_ _0077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_230_3277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8265_ _3880_ _3885_ _2140_ _3886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5477_ _1563_ _0047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7216_ _2567_ _2986_ _3140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8196_ _3802_ _3821_ _3822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7862__A2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input48_I i_req_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__A2 _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7147_ core_0.decode.oc_alu_mode\[3\] _2360_ _3073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__8811__A1 _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7614__A2 _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7078_ _2711_ _3004_ _3005_ _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_198_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5625__A1 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5476__I1 net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6029_ core_0.execute.rf.reg_outputs\[15\]\[4\] _0944_ _2019_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_198_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8007__B _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7378__B2 core_0.execute.sreg_scratch.o_d\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output204_I net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5389__B1 _1494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5928__A2 _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_232_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A2 net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8878__A1 _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6889__B1 _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6353__A2 _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8677__B _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7581__B _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6105__A2 _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7853__A2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_2504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5864__A1 _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7066__B1 _2991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8802__A1 core_0.execute.pc_high_buff_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__A1 _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5467__I1 net62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8030__A2 _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_177_2633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__A1 core_0.execute.rf.reg_outputs\[6\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6041__B2 core_0.execute.rf.reg_outputs\[12\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8869__A1 core_0.execute.pc_high_buff_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_73_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7136__A4 _1865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6344__A2 _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5400_ _1262_ _1266_ _1299_ _1503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6380_ _1668_ _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_113_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5331_ _1266_ _1281_ _1449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8050_ _3647_ _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5262_ core_0.dec_jump_cond_code\[1\] core_0.dec_jump_cond_code\[0\] core_0.execute.alu_flag_reg.o_d\[0\]
+ _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7844__A2 _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_2773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7001_ _1329_ _2929_ _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4658__A2 _0698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5855__A1 _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5193_ core_0.decode.oc_alu_mode\[2\] _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7057__B1 _2978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5607__A1 core_0.decode.i_instr_l\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9253__CLK clknet_leaf_1_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8952_ core_0.decode.i_imm_pass\[8\] _1264_ _4444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5231__S _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6280__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7903_ core_0.execute.rf.reg_outputs\[7\]\[13\] _3634_ _3636_ _3645_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8883_ _0912_ _4383_ _4400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_203_2943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_203_2954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4830__A2 net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7834_ core_0.ew_reg_ie\[8\] _3395_ _3605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_210_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6032__A1 core_0.execute.rf.reg_outputs\[9\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_219_3139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7666__B _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7765_ _3409_ _3563_ _3566_ _0332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4977_ core_0.fetch.prev_request_pc\[15\] _1156_ _1157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_191_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_175_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_1964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7780__A1 core_0.execute.rf.reg_outputs\[10\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6583__A2 _2054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6716_ core_0.execute.rf.reg_outputs\[7\]\[5\] _2611_ _2612_ core_0.execute.rf.reg_outputs\[5\]\[5\]
+ _2653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9504_ _0514_ clknet_leaf_123_i_clk core_0.execute.alu_mul_div.mul_res\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4594__A1 core_0.execute.rf.reg_outputs\[2\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_rebuffer40_I net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7696_ core_0.execute.rf.reg_outputs\[12\]\[4\] _3526_ _3513_ _3527_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9435_ _0445_ clknet_leaf_45_i_clk core_0.execute.rf.reg_outputs\[3\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6647_ _2000_ _1957_ _2589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7532__A1 _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__A3 _1289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5543__B1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9366_ _0376_ clknet_leaf_151_i_clk core_0.execute.rf.reg_outputs\[8\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_2316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6578_ net101 _2520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4897__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8317_ core_0.execute.alu_mul_div.mul_res\[9\] _3933_ _3934_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_42_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5529_ _0896_ _1367_ _1591_ _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8088__A2 _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9297_ _0307_ clknet_leaf_31_i_clk core_0.execute.rf.reg_outputs\[12\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8248_ _3862_ _3869_ _3870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5846__A1 _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output154_I net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8179_ _1543_ _1894_ _3805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_243_3424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7599__A1 _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_213_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8260__A2 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_2445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8012__A2 _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6023__A1 core_0.execute.rf.reg_outputs\[8\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7523__A1 net36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_172_2574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9126__CLK clknet_leaf_108_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8079__A2 _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7826__A2 _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5837__A1 _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9276__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5301__A3 _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4890__S _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4900_ core_0.fetch.pc_flush_override _1079_ _1080_ _1081_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8003__A2 _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5880_ _0881_ _0882_ _0883_ _0884_ _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_153_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__A1 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4831_ core_0.fetch.out_buffer_data_instr\[1\] _1012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_185_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_173_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6565__A2 _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7762__A1 core_0.execute.rf.reg_outputs\[10\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7550_ _3396_ _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_28_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4762_ core_0.dec_l_reg_sel\[2\] _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__4576__B2 core_0.execute.rf.reg_outputs\[3\]\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6501_ _2442_ _2443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7481_ core_0.dec_rf_ie\[9\] core_0.ew_reg_ie\[9\] _3366_ _3374_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4693_ core_0.execute.rf.reg_outputs\[2\]\[1\] net250 _0695_ core_0.execute.rf.reg_outputs\[10\]\[1\]
+ _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_126_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6317__A2 _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9220_ _0231_ clknet_leaf_92_i_clk net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6432_ core_0.execute.mem_stage_pc\[5\] _2395_ _2387_ _2397_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4879__A2 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9151_ _0163_ clknet_leaf_41_i_clk net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6363_ _2334_ _1962_ _2335_ _2336_ _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_8102_ core_0.execute.rf.reg_outputs\[1\]\[0\] _3760_ _3756_ _3761_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5314_ _1006_ _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_140_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9082_ _0107_ clknet_leaf_101_i_clk core_0.decode.i_imm_pass\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7817__A2 _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6294_ _1547_ _2268_ _2224_ _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_178_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5828__A1 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8033_ core_0.execute.rf.reg_outputs\[3\]\[3\] _3716_ _3718_ _3721_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5245_ _0895_ _0896_ _1008_ _1367_ _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__6096__A4 _0980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8764__C _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ _1267_ _1319_ _1323_ _1324_ _1325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_199_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_242_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_235_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer88_I _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8935_ _2709_ _1486_ _4435_ _4307_ _0633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_210_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10__f_i_clk clknet_3_5_0_i_clk clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8866_ _4383_ _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_38_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7817_ _3447_ _3585_ _3596_ _0354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8797_ _1433_ _4325_ _4326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_109_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__B2 core_0.execute.rf.reg_outputs\[12\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7748_ _3457_ _3543_ _3556_ _0325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_163_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7679_ _3466_ _3498_ _3516_ _0296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9418_ _0428_ clknet_leaf_137_i_clk core_0.execute.rf.reg_outputs\[4\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5644__B _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9299__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9349_ _0359_ clknet_leaf_152_i_clk core_0.execute.rf.reg_outputs\[9\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_246_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output79_I net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8481__A2 _4040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8674__C _4201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6492__A1 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_21_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__A2 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4774__I core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7992__A1 _3408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_174_2603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5770__A3 _1757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap217 _0859_ net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_52_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4730__A1 core_0.execute.pc_high_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_2732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6483__A1 net264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5286__A2 net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5030_ _1086_ _1200_ _1201_ _1162_ net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_209_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8224__A2 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7283__I0 core_0.ew_data\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6981_ _2009_ _1960_ _2910_ _2006_ _2911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_177_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7983__A1 _3469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8720_ _4276_ _4277_ _0576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4797__A1 core_0.ew_reg_ie\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5932_ _1920_ _1921_ _1922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_200_2913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4797__B2 core_0.ew_reg_ie\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8651_ _4203_ _4060_ _1661_ _4221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_180_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5863_ net314 net199 _1852_ _1853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__4633__B _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7735__A1 _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_196_2861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_216_3109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7602_ core_0.execute.rf.reg_outputs\[15\]\[14\] _3396_ _3467_ _3471_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4814_ core_0.ew_submit _0927_ _0994_ _0995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__4549__A1 core_0.execute.rf.reg_outputs\[3\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8582_ _2123_ _4160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5794_ _0942_ _0947_ net329 _0958_ _1784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_146_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7533_ _3382_ core_0.ew_data\[2\] _3413_ _3414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__7944__B _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4745_ _0925_ _0926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_32_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7464_ core_0.dec_rf_ie\[1\] core_0.ew_reg_ie\[1\] _2419_ _3365_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4676_ core_0.execute.rf.reg_outputs\[4\]\[2\] _0720_ _0683_ core_0.execute.rf.reg_outputs\[7\]\[2\]
+ _0861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_126_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8160__A1 _3453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9203_ _0214_ clknet_leaf_77_i_clk core_0.ew_data\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_189_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6415_ _1433_ _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_43_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7395_ _3313_ _3312_ _3314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_102_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__C _2217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9134_ _0146_ clknet_leaf_116_i_clk core_0.execute.alu_mul_div.div_cur\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6346_ _2321_ _2322_ _0157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9065_ _0090_ clknet_leaf_114_i_clk core_0.decode.i_instr_l\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_227_3238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8463__A2 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6277_ _2249_ _2261_ _2141_ _2262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8016_ _3462_ _3695_ _3710_ _0439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5277__A2 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5228_ _1359_ net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5816__A4 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input30_I i_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_243_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_2248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5159_ _1244_ _1310_ _1264_ _1311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5029__A2 _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6226__A1 _2206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6777__A2 _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7974__A1 _3456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__A1 _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8918_ _1231_ _1455_ _4422_ _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8849_ _4335_ _4370_ _4371_ _4372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6529__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7726__A1 _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_3367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8015__B _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_2388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8151__A1 net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7145__I core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__A1 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4476__B1 _0673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6217__A1 core_0.execute.alu_mul_div.div_cur\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_180_2673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6768__A2 _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7965__A1 core_0.execute.rf.reg_outputs\[5\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4779__A1 core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5976__B1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7717__A1 core_0.execute.rf.reg_outputs\[12\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8390__A1 core_0.execute.alu_mul_div.mul_res\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7764__B _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4530_ core_0.execute.rf.reg_outputs\[13\]\[14\] net284 _0710_ core_0.execute.rf.reg_outputs\[8\]\[14\]
+ _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8142__A1 _3408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_211_3039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6200_ _2186_ _2188_ _2189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7180_ _2586_ _2932_ _3105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4703__B2 core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6131_ _2006_ _2120_ _2121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5504__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_55_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _2050_ _2051_ _2052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5013_ _0895_ net55 _1188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_0_Left_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_183_Right_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6208__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_222_3179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6759__A2 net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7956__A1 _3414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_5_Right_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_37_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6964_ net81 _2829_ _2892_ _2893_ _2894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_177_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5431__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8703_ core_0.execute.sreg_irq_pc.o_d\[11\] _4202_ _4264_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_193_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5915_ core_0.execute.rf.reg_outputs\[14\]\[9\] _1802_ _1781_ core_0.execute.rf.reg_outputs\[10\]\[9\]
+ _1905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_140_2189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6895_ _2823_ _2824_ _2825_ _2826_ _2827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7708__A1 _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8905__B1 _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6134__I core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5846_ _1518_ net181 _1836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8634_ _1226_ _1699_ _4204_ _4205_ _4206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_8_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7184__A2 _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8381__A1 core_0.execute.alu_mul_div.mul_res\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7674__B _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5195__A1 _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8565_ _4144_ _4145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5777_ _1765_ _1766_ _1767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_106_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6931__A2 _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7516_ net21 _1349_ _3399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4728_ core_0.execute.prev_pc_high\[2\] _0904_ _0905_ core_0.execute.prev_pc_high\[1\]
+ _0909_ _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_210_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_1925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8496_ net82 _4076_ _4084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8133__A1 _3469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7447_ _3356_ _0224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4659_ _0842_ _0843_ _0844_ _0845_ _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_142_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5498__A2 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7378_ core_0.execute.sreg_irq_pc.o_d\[14\] _3042_ _3044_ core_0.execute.sreg_scratch.o_d\[14\]
+ _3298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9117_ _0129_ clknet_leaf_64_i_clk core_0.execute.sreg_priv_control.o_d\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6329_ _2161_ _2307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8436__A2 _4031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6447__A1 _1185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9048_ _0074_ clknet_leaf_83_i_clk core_0.fetch.prev_request_pc\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__6998__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_150_Right_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_203_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7849__B _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7947__A1 _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__B1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5958__C2 core_0.execute.rf.reg_outputs\[3\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_2406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4630__B1 net312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8372__A1 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_205_Left_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4933__A1 core_0.fetch.prev_request_pc\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_239_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5489__A2 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_2535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_2546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_219_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_182_2702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_214_Left_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_207_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6989__A2 core_0.execute.alu_mul_div.mul_res\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5110__A1 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__B1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5413__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5700_ _1417_ _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_102_1737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6680_ _2614_ _2620_ _2621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_193_2831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7166__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_223_Left_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_143_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8363__A1 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5631_ _1049_ _1628_ _1651_ _0113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_214_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8350_ core_0.execute.alu_mul_div.mul_res\[11\] _3830_ _3965_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5562_ core_0.fetch.prev_request_pc\[13\] _1082_ _1083_ net164 _1611_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__4924__A1 core_0.fetch.prev_request_pc\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8115__A1 core_0.execute.rf.reg_outputs\[1\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4924__B2 core_0.fetch.prev_request_pc\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ core_0.execute.alu_mul_div.div_res\[12\] _1742_ _3222_ _3223_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4513_ core_0.execute.rf.reg_outputs\[13\]\[15\] _0708_ _0710_ core_0.execute.rf.reg_outputs\[8\]\[15\]
+ _0711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8281_ core_0.execute.alu_mul_div.mul_res\[6\] _3894_ _3900_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8666__A2 _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5493_ core_0.fetch.out_buffer_data_instr\[14\] _1573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_130_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6677__A1 core_0.execute.rf.reg_outputs\[1\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7232_ _1683_ core_0.execute.sreg_irq_pc.o_d\[10\] _3156_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6677__B2 core_0.execute.rf.reg_outputs\[3\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4688__B1 net347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7163_ core_0.execute.sreg_priv_control.o_d\[8\] _1693_ _2996_ net15 _2689_ _3089_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_113_1866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6114_ _2091_ _2103_ _2104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_244_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8969__A3 _1272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7094_ _1894_ _3020_ _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6045_ core_0.execute.rf.reg_outputs\[5\]\[5\] net225 _1801_ core_0.execute.rf.reg_outputs\[14\]\[5\]
+ _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_241_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_68_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_9_i_clk clknet_4_2__leaf_i_clk clknet_leaf_9_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_240_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_206_2985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7996_ _3420_ _3694_ _3699_ _0430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ core_0.execute.alu_flag_reg.o_d\[3\] _2770_ _2774_ core_0.execute.sreg_irq_pc.o_d\[3\]
+ _2878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4612__B1 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_235_3337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6878_ _1749_ _2005_ _2810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7157__A2 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8617_ _2989_ _3035_ _4190_ _4191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5168__A1 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5829_ _1818_ _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_9597_ _0607_ clknet_leaf_61_i_clk core_0.execute.pc_high_out\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_146_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4915__A1 core_0.fetch.prev_request_pc\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__B2 core_0.fetch.prev_request_pc\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8548_ _1736_ _4127_ _4128_ _4129_ _4130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8106__A1 core_0.execute.rf.reg_outputs\[1\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_2347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output184_I net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6117__B1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5208__I _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8479_ _2393_ _4058_ _4069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6668__A1 core_0.execute.rf.reg_outputs\[1\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6668__B2 core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A1 _1294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_246_3466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7093__A1 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8682__C _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5643__A2 _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_2476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__I net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8254__I core_0.execute.alu_mul_div.mul_res\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7396__A2 _3069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_72_Left_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_200_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7148__A2 net306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6930__C _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A1 _1244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8896__A2 _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6108__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8648__A2 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput208 net245 sr_bus_data_o[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_81_Left_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5331__A1 _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6377__C core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5882__A2 _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8873__B _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8820__A2 _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5634__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_210_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_90_Left_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7850_ _3435_ _3606_ _3615_ _0368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7387__A2 _3297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8584__A1 _2816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6801_ _1895_ _2733_ _2734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_187_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5398__A1 _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4993_ core_0.fetch.prev_request_pc\[13\] _1154_ _1171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7781_ _3451_ _3563_ _3575_ _0339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9520_ _0530_ clknet_leaf_120_i_clk core_0.execute.alu_mul_div.div_res\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6732_ core_0.execute.rf.reg_outputs\[1\]\[7\] _2608_ _2609_ core_0.execute.rf.reg_outputs\[3\]\[7\]
+ _2667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_147_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8336__A1 _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6663_ _1765_ _1866_ _2603_ _2604_ _2605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_9451_ _0461_ clknet_leaf_136_i_clk core_0.execute.rf.reg_outputs\[2\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8887__A2 _4383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4641__B _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5229__S _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8113__B _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6898__A1 net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8402_ _4000_ _3832_ _4010_ _4012_ _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5614_ _1043_ _1615_ _1642_ _0105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_139_2180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9382_ _0392_ clknet_leaf_154_i_clk core_0.execute.rf.reg_outputs\[7\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6594_ _2465_ _2535_ _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5545_ core_0.fetch.prev_request_pc\[5\] _1595_ _1084_ net171 _1602_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_8333_ _3940_ _3833_ _3948_ _3828_ _3949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_171_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_230_3267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_230_3278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8767__C _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8264_ _3882_ _3884_ _1669_ _3885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5476_ core_0.fetch.out_buffer_data_instr\[7\] net66 _1559_ _1563_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_142_i_clk clknet_4_1__leaf_i_clk clknet_leaf_142_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7215_ _2592_ _2575_ _2588_ _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8195_ _1743_ core_0.execute.alu_mul_div.comp _3812_ _3820_ _3821_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_245_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6287__C _2217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5873__A2 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7146_ _1766_ _1886_ _1887_ _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_226_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7075__A1 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7077_ _2963_ _3003_ _3005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5625__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6822__A1 core_0.decode.oc_alu_mode\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6028_ core_0.execute.rf.reg_outputs\[14\]\[4\] _0957_ _0958_ _0980_ _2018_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_EDGE_ROW_129_Left_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8575__A1 _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7378__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__A1 core_0.decode.i_imm_pass\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5389__B2 core_0.decode.i_instr_l\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7979_ _3647_ _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_193_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_166_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8327__A1 _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9649_ _0659_ clknet_leaf_140_i_clk core_0.dec_rf_ie\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6889__A1 core_0.execute.alu_mul_div.div_cur\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_138_Left_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7862__B _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__A1 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8677__C _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__A2 _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4777__I core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_2505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__A2 net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7066__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_147_Left_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_205_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8566__A1 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6026__C1 _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6941__B _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6041__A2 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_2634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6660__C _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8869__A2 _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_16_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6232__I _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7772__B _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5552__A1 _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4888__S _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5330_ _1445_ _1447_ _1448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ core_0.dec_jump_cond_code\[1\] _1380_ _1381_ core_0.dec_jump_cond_code\[0\]
+ _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_227_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_2763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_2774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_8__f_i_clk clknet_3_4_0_i_clk clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7000_ _1899_ net218 _2732_ _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5855__A2 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_74_i_clk clknet_4_11__leaf_i_clk clknet_leaf_74_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5192_ _1231_ _1335_ _1336_ _0006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_110_1836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7057__A1 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6804__A1 _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5607__A2 _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8951_ _1839_ _0038_ _4443_ _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_222_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8108__B _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_89_i_clk clknet_4_15__leaf_i_clk clknet_leaf_89_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7012__B core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7902_ _3463_ _3629_ _3644_ _0391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6280__A2 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8882_ _4386_ _4398_ _4399_ _0616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5311__I _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_203_2944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8557__A1 _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_210_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7833_ _3473_ _3586_ _3604_ _0362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_188_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6032__A2 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7764_ core_0.execute.rf.reg_outputs\[10\]\[1\] _3564_ _3554_ _3566_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4976_ core_0.fetch.prev_request_pc\[14\] _1155_ _1156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7780__A2 _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_121_1965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9503_ _0513_ clknet_leaf_125_i_clk core_0.execute.alu_mul_div.mul_res\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6715_ core_0.execute.rf.reg_outputs\[1\]\[5\] _2608_ _2609_ core_0.execute.rf.reg_outputs\[3\]\[5\]
+ _2652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_117_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4594__A2 _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7695_ _3519_ _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9434_ _0444_ clknet_leaf_37_i_clk core_0.execute.rf.reg_outputs\[3\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_18_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6646_ _2582_ _2588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7682__B _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_27_i_clk clknet_4_2__leaf_i_clk clknet_leaf_27_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5543__A1 core_0.fetch.prev_request_pc\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9365_ _0375_ clknet_leaf_150_i_clk core_0.execute.rf.reg_outputs\[8\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_150_2317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5543__B2 net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _2516_ _2517_ _2518_ _2519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_30_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8316_ _1679_ _1539_ _3880_ _3932_ _3933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__4751__C1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5528_ _0895_ _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_41_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input60_I i_req_data[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9296_ _0306_ clknet_leaf_32_i_clk core_0.execute.rf.reg_outputs\[12\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5459_ net38 _1552_ _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8247_ _1535_ _3868_ _3869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_246_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A2 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8178_ _1534_ _3803_ _3804_ _0507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_243_3425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7048__A1 _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7129_ core_0.ew_data\[7\] _2642_ _3056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7599__A2 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_2446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6271__A2 _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8548__A1 _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_87_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7857__B _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6761__B _2694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7220__A1 net247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6023__A2 net345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5534__A1 _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_172_2575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6731__B1 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_1691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7287__A1 _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8484__B1 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_155_Left_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_207_3000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8787__A1 core_0.execute.sreg_irq_flags.o_d\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6655__C _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5131__I _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8539__A1 _1180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7211__A1 _2480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_164_Left_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4830_ _0894_ net38 _1010_ _1011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_157_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7762__A2 _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4761_ core_0.dec_l_reg_sel\[3\] _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4576__A2 net297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6970__B1 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6500_ _2074_ _2090_ _2442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7480_ _3373_ _0240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4692_ core_0.execute.rf.reg_outputs\[6\]\[1\] _0670_ net318 core_0.execute.rf.reg_outputs\[4\]\[1\]
+ core_0.execute.rf.reg_outputs\[1\]\[1\] _0693_ _0876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__8711__A1 net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6431_ _1211_ _2385_ _2396_ _0168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6722__B1 _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ _2097_ _2098_ _2099_ _2100_ _2336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_9150_ _0162_ clknet_leaf_96_i_clk core_0.de_jmp_pred vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_178_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5313_ _1432_ _0014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8101_ _3758_ _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_141_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9220__CLK clknet_leaf_92_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_173_Left_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6293_ _2221_ _2275_ _2276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9081_ _0106_ clknet_leaf_101_i_clk core_0.decode.i_imm_pass\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_228_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5828__A2 _1790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8032_ _3414_ _3715_ _3720_ _0445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5244_ core_0.decode.i_flush core_0.fetch.flush_event_invalidate _1367_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_228_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4887__I0 net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5175_ _1234_ _1236_ _1269_ _1324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_236_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_194_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8934_ _1482_ _1490_ _1522_ _4435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_78_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8780__C _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8865_ _4385_ _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_94_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6005__A2 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8352__I core_0.execute.alu_mul_div.mul_res\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7816_ core_0.execute.rf.reg_outputs\[9\]\[7\] _3591_ _3595_ _3596_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8796_ _4322_ _4323_ _4324_ _4325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7753__A2 _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4567__A2 _0685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7747_ core_0.execute.rf.reg_outputs\[11\]\[10\] _3548_ _3554_ _3556_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4959_ _1071_ _1139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6961__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7678_ core_0.execute.rf.reg_outputs\[13\]\[13\] _3504_ _3513_ _3516_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_151_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7505__A2 core_0.ew_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8702__A1 _4249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5516__A1 net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9417_ _0427_ clknet_leaf_14_i_clk core_0.execute.rf.reg_outputs\[4\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6629_ _2570_ _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_117_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9348_ _0358_ clknet_leaf_6_i_clk core_0.execute.rf.reg_outputs\[9\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_197_Right_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9279_ _0289_ clknet_leaf_32_i_clk core_0.execute.rf.reg_outputs\[13\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5819__A2 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6492__A2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8769__A1 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_214_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7992__A2 _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8941__A1 _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_2604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4558__A2 _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5755__A1 _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5770__A4 _1759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9243__CLK clknet_leaf_2_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_213_3070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_164_Right_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4730__A2 net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_2733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7680__A1 core_0.execute.rf.reg_outputs\[13\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__A3 net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8881__B _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7432__A1 net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7283__I1 _3205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6980_ _2009_ _2073_ _2074_ _2910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_205_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7983__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5931_ core_0.execute.rf.reg_outputs\[6\]\[8\] net219 _1787_ core_0.execute.rf.reg_outputs\[3\]\[8\]
+ _1921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4797__A2 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_200_2914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8650_ _2391_ _4217_ _4218_ _4219_ _4220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7196__B1 _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5862_ _1518_ net183 _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XTAP_TAPCELL_ROW_196_2862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8932__A1 core_0.dec_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7735__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7601_ _3469_ _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5746__A1 _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4549__A2 _0698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4813_ _0993_ _0994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_91_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8581_ _1419_ _2770_ _4159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_200_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5793_ _1771_ _1774_ _1777_ _1782_ _1783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_28_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7532_ _3381_ _3411_ _3412_ _3413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_28_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4744_ core_0.execute.hold_valid core_0.decode.o_submit _0923_ _0924_ _0925_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_28_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7463_ _3364_ _0232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4675_ core_0.execute.rf.reg_outputs\[6\]\[2\] _0670_ net250 core_0.execute.rf.reg_outputs\[2\]\[2\]
+ _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5237__S _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8160__A2 _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9202_ _0213_ clknet_leaf_77_i_clk core_0.ew_data\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_43_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__I net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6414_ _1226_ _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6171__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7394_ _2483_ _3279_ _3313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_3_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6710__A3 _2640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9133_ _0145_ clknet_leaf_116_i_clk core_0.execute.alu_mul_div.div_cur\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_141_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4721__A2 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_131_Right_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6345_ core_0.execute.alu_mul_div.div_cur\[13\] _2218_ _0999_ _2322_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5036__I net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9064_ _0089_ clknet_leaf_114_i_clk core_0.decode.i_instr_l\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6276_ _2211_ _2260_ _2261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_227_3239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5227_ core_0.ew_data\[1\] core_0.ew_data\[9\] _1349_ _1359_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8015_ core_0.execute.rf.reg_outputs\[4\]\[12\] _3700_ _3704_ _3710_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7671__A1 _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_138_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6295__C _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5158_ _1243_ _1273_ _1310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_243_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input23_I i_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5089_ core_0.decode.i_instr_l\[5\] _1245_ _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7974__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8917_ core_0.dec_sreg_load _1286_ _4422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8848_ core_0.execute.pc_high_buff_out\[6\] _4335_ _4371_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7726__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_238_3368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8779_ core_0.execute.sreg_scratch.o_d\[15\] _4293_ _4314_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_2389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8031__B _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4960__A2 _1139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8151__A2 _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output91_I net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7870__B _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__A2 _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7662__A1 core_0.execute.rf.reg_outputs\[13\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4476__A1 core_0.execute.rf.reg_outputs\[6\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6217__A2 net239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_180_2674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7965__A2 _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5976__A1 core_0.execute.rf.reg_outputs\[6\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4779__A2 core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5976__B2 core_0.execute.rf.reg_outputs\[12\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7717__A2 _3519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__A1 _0765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_233_Right_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8390__A2 _2375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5057__S _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8142__A2 _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7780__B _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5900__A1 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4703__A2 net303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ _2011_ _2073_ _2075_ _2119_ _2120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_194_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8167__I _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6061_ core_0.execute.rf.reg_outputs\[6\]\[7\] net219 _1787_ core_0.execute.rf.reg_outputs\[3\]\[7\]
+ _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_225_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5012_ _1158_ _1152_ _1186_ _1187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_225_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6208__A2 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7956__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6759__A3 _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6963_ _2694_ _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_37_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8702_ _4249_ core_0.execute.mem_stage_pc\[11\] _4260_ _4262_ _4209_ _4263_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6415__I _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ core_0.execute.rf.reg_outputs\[9\]\[9\] _1815_ _1799_ core_0.execute.rf.reg_outputs\[6\]\[9\]
+ core_0.execute.rf.reg_outputs\[1\]\[9\] _1779_ _1904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_220_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6894_ core_0.execute.irq_en _1692_ _2777_ core_0.execute.sreg_irq_flags.o_d\[2\]
+ _2826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_191_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7708__A2 _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7955__B _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8633_ core_0.dec_wfi _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5719__A1 _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5845_ net313 net195 _1834_ _1835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XPHY_EDGE_ROW_200_Right_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8381__A2 _2375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8630__I _4201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8564_ _1736_ _4141_ _4142_ _4143_ _4144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_173_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5195__A2 _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5776_ _1328_ core_0.decode.oc_alu_mode\[13\] _1766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_clkbuf_leaf_64_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_101_Left_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_133_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7515_ net35 _1347_ _3398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4727_ core_0.execute.prev_pc_high\[0\] _0908_ _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_133_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8495_ _4051_ _4083_ _0545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_118_1926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8133__A2 _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6150__I core_0.execute.alu_mul_div.cbit\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7446_ net128 _3085_ _2415_ _3356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4658_ core_0.execute.rf.reg_outputs\[3\]\[4\] _0698_ _0716_ _0845_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7892__A1 _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7377_ _2142_ _0997_ _3295_ _3296_ _3297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_4589_ core_0.execute.rf.reg_outputs\[7\]\[9\] net297 _0697_ core_0.execute.rf.reg_outputs\[3\]\[9\]
+ _0781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9116_ _0128_ clknet_leaf_119_i_clk core_0.execute.alu_mul_div.cbit\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6328_ _2299_ _2256_ _2306_ _2229_ _0155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_229_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6447__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7644__A1 _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9047_ _0073_ clknet_leaf_83_i_clk core_0.fetch.prev_request_pc\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6259_ _2219_ _2244_ _2245_ _2229_ _0147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_244_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_110_Left_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_212_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7947__A2 _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__B2 core_0.execute.rf.reg_outputs\[12\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8026__B _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_2407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6383__A1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5186__A2 _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4933__A2 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8124__A2 _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6135__A1 _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_239_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_2536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_238_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Right_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6438__A2 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_246_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5110__A2 _1254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9431__CLK clknet_leaf_144_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7938__A2 _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8060__A1 _3472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6235__I _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9581__CLK clknet_leaf_21_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_102_1738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7166__A3 _3091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_2832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8363__A2 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5630_ core_0.decode.i_imm_pass\[9\] _1645_ _1651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5561_ _1608_ _1610_ _0084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4924__A2 _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8115__A2 _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7300_ _1743_ _3220_ _3221_ _0996_ _3222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_26_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6126__A1 _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4512_ _0709_ _0710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8280_ _3899_ _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5492_ _1571_ _1551_ _1572_ _0053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6677__A2 _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7231_ core_0.execute.alu_mul_div.div_cur\[10\] _1317_ _3152_ _3154_ _3155_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_111_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4688__A1 core_0.execute.rf.reg_outputs\[5\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7162_ core_0.execute.sreg_irq_pc.o_d\[8\] _3042_ _3044_ core_0.execute.sreg_scratch.o_d\[8\]
+ _3088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_113_1867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6113_ _1875_ _2102_ _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7093_ _2009_ _2561_ _2716_ _3020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7477__I1 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6044_ core_0.execute.rf.reg_outputs\[1\]\[5\] _1778_ _1803_ core_0.execute.rf.reg_outputs\[11\]\[5\]
+ _2034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_119_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8625__I core_0.execute.irq_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7929__A2 _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8051__A1 core_0.execute.rf.reg_outputs\[3\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_206_2986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7995_ core_0.execute.rf.reg_outputs\[4\]\[3\] _3695_ _3689_ _3699_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6601__A2 _2366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6946_ core_0.execute.pc_high_buff_out\[3\] _2771_ _2777_ core_0.execute.sreg_irq_flags.o_d\[3\]
+ _2877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_135_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4612__A1 core_0.execute.rf.reg_outputs\[10\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_235_3327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5984__I _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6877_ _1751_ _2806_ _2808_ _1894_ _2809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_147_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_235_3338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8616_ _2918_ _2949_ _4190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5168__A2 _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5828_ _0950_ _1790_ _1818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_162_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9596_ _0606_ clknet_leaf_61_i_clk core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_63_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8547_ _1685_ core_0.execute.sreg_irq_pc.o_d\[12\] net196 _2134_ _2136_ _4129_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_173_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4915__A2 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5759_ _1748_ _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_134_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8106__A2 _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_2348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6117__A1 core_0.execute.rf.reg_outputs\[7\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8478_ _4066_ _4068_ _4051_ _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6668__A2 _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7865__A1 _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output177_I net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7429_ _3347_ _0215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_246_3467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8290__A1 core_0.execute.alu_mul_div.mul_res\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6764__B _2135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_2477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8042__A1 core_0.execute.rf.reg_outputs\[3\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7305__B1 _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput209 net209 sr_bus_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7856__A1 _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7608__A1 core_0.ew_reg_ie\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8281__A1 core_0.execute.alu_mul_div.mul_res\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5095__A1 core_0.decode.oc_alu_mode\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_128_2052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6831__A2 core_0.execute.alu_mul_div.i_div vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4842__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8033__A1 core_0.execute.rf.reg_outputs\[3\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6044__B1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_172_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6800_ _1882_ net214 _2732_ _2733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8584__A2 _2868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7780_ core_0.execute.rf.reg_outputs\[10\]\[8\] _3570_ _3568_ _3575_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5398__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4992_ net75 _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_148_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ core_0.execute.rf.reg_outputs\[7\]\[7\] _2611_ _2612_ core_0.execute.rf.reg_outputs\[5\]\[7\]
+ _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_187_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8336__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9450_ _0460_ clknet_leaf_136_i_clk core_0.execute.rf.reg_outputs\[2\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_63_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6662_ core_0.decode.oc_alu_mode\[13\] _1763_ _2604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8401_ _4011_ _4012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6898__A2 _2829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5613_ core_0.decode.i_imm_pass\[1\] _1616_ _1642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9381_ _0391_ clknet_leaf_155_i_clk core_0.execute.rf.reg_outputs\[7\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_139_2181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6593_ _2155_ _1942_ _2535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8332_ _3945_ _3947_ _3948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5544_ _1597_ _1601_ _0076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_230_3268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7847__A1 core_0.execute.rf.reg_outputs\[8\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9477__CLK clknet_leaf_145_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8263_ _1541_ _2040_ _3883_ _3884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5475_ _1562_ _0046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_197_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7214_ _2795_ _3136_ _3137_ _3138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_111_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8194_ _1537_ _3819_ _3820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4530__B1 _0710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7145_ core_0.decode.oc_alu_mode\[7\] _3071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__7460__S _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8272__A1 core_0.execute.alu_mul_div.mul_res\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7076_ _2963_ _3003_ _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_225_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6027_ core_0.execute.rf.reg_outputs\[1\]\[4\] _0954_ _0955_ _0962_ _2017_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4833__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5389__A2 _1488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7978_ _3462_ _3673_ _3688_ _0423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_221_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6929_ _2076_ _2738_ _2860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_193_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8304__B _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8327__A2 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9648_ _0658_ clknet_leaf_139_i_clk core_0.dec_rf_ie\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6889__A2 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9579_ _0589_ clknet_leaf_21_i_clk core_0.execute.sreg_scratch.o_d\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_242_Left_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7838__A1 _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6510__A1 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_2506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4521__B1 net303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7066__A2 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_216_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__A1 core_0.dec_wfi vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8015__A1 core_0.execute.rf.reg_outputs\[4\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6026__B1 net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8566__A2 _4052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4588__B1 net316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_2635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7609__I _3475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5001__A1 _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_8_i_clk clknet_4_2__leaf_i_clk clknet_leaf_8_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_23_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7829__A1 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_239_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5260_ core_0.execute.alu_flag_reg.o_d\[2\] core_0.execute.alu_flag_reg.o_d\[0\]
+ _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_188_2764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5191_ core_0.decode.oc_alu_mode\[3\] _1286_ _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_110_1837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7057__A2 _2438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6804__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8950_ core_0.decode.i_imm_pass\[7\] _1264_ _4443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_222_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7901_ core_0.execute.rf.reg_outputs\[7\]\[12\] _3634_ _3636_ _3644_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8006__A1 _3446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8881_ core_0.execute.pc_high_buff_out\[3\] _4385_ _3797_ _4399_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_203_2945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7832_ core_0.execute.rf.reg_outputs\[9\]\[15\] _3584_ _3595_ _3604_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6568__A1 _1759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4579__B1 _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7763_ _3402_ _3563_ _3565_ _0331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4975_ core_0.fetch.prev_request_pc\[13\] _1154_ _1155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_59_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8124__B _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7519__I _3401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9502_ _0512_ clknet_leaf_124_i_clk core_0.execute.alu_mul_div.mul_res\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6714_ _2422_ _2650_ _2651_ _0195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_1966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6423__I net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7694_ _3421_ _3520_ _3525_ _0302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_178_Right_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7963__B _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9433_ _0443_ clknet_leaf_25_i_clk core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_190_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6645_ _2586_ _2587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8778__C _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9364_ _0374_ clknet_leaf_7_i_clk core_0.execute.rf.reg_outputs\[8\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5543__A2 _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6576_ _2439_ _2488_ _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6740__A1 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_2307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer26_I _1745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_2318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8315_ _1538_ _3930_ _3931_ _1679_ _3932_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5527_ _1021_ _1552_ _1590_ _0070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4751__B1 _0930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4751__C2 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9295_ _0305_ clknet_leaf_31_i_clk core_0.execute.rf.reg_outputs\[12\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8493__A1 _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8246_ _2139_ _3823_ _3867_ _3868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5458_ _1550_ _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input53_I i_req_data[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8794__B _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4503__B1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8177_ _1543_ _1534_ _3804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5389_ core_0.decode.i_imm_pass\[0\] _1488_ _1494_ core_0.decode.i_instr_l\[11\]
+ _1495_ _1496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_243_3426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7128_ _2709_ _3053_ _3054_ _3055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5059__A1 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__B _2710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7059_ _2587_ _2813_ _2987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_199_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_161_2447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6559__A1 _2433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7220__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_145_Right_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_181_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5534__A2 net160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6731__A1 core_0.execute.rf.reg_outputs\[7\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_2576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6731__B2 core_0.execute.rf.reg_outputs\[5\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8484__A1 net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8484__B2 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_207_3001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8787__A2 _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6798__A1 _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9172__CLK clknet_leaf_42_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_141_i_clk clknet_4_4__leaf_i_clk clknet_leaf_141_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_158_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_218_3130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _0935_ _0940_ net293 _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6970__B2 _1865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_60_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_112_Right_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4691_ _0871_ _0872_ _0873_ _0874_ _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_70_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8711__A2 _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6430_ core_0.execute.mem_stage_pc\[4\] _2395_ _2387_ _2396_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6722__A1 core_0.execute.rf.reg_outputs\[1\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6722__B2 core_0.execute.rf.reg_outputs\[3\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6361_ _2092_ _2093_ _2094_ _2095_ _2335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XPHY_EDGE_ROW_49_Right_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8100_ _3758_ _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5312_ _1431_ _1428_ _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__8475__A1 _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9080_ _0105_ clknet_leaf_100_i_clk core_0.decode.i_imm_pass\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_140_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6292_ _2186_ _2274_ _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5289__A1 net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8031_ core_0.execute.rf.reg_outputs\[3\]\[2\] _3716_ _3718_ _3720_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5243_ net17 net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_87_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8227__A1 _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5174_ _1321_ _1322_ _1323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8119__B _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7023__B _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8778__A2 _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6789__A1 _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5322__I core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_2280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7450__A2 _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7958__B _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8933_ _1231_ _1493_ _4434_ _0632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Right_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8633__I core_0.dec_wfi vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8864_ _4383_ _4384_ _1400_ _4385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_149_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_109_i_clk clknet_4_12__leaf_i_clk clknet_leaf_109_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7202__A2 _3126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7815_ _3512_ _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8795_ core_0.dec_sreg_store _2775_ _4324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_59_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__A1 core_0.ew_data\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8950__A2 _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7746_ _3454_ _3542_ _3555_ _0324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_164_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4958_ _1134_ _1135_ _1136_ _1137_ _1138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__6961__A1 core_0.execute.alu_flag_reg.o_d\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_134_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6961__B2 net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7693__B _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7677_ _3463_ _3498_ _3515_ _0295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_191_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4889_ _1068_ _1069_ _1070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9416_ _0426_ clknet_leaf_136_i_clk core_0.execute.rf.reg_outputs\[5\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6628_ _1895_ _2569_ _2570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_117_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5516__A2 _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_67_Right_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__B1 _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9347_ _0357_ clknet_leaf_6_i_clk core_0.execute.rf.reg_outputs\[9\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6559_ _2433_ _2435_ _2501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_120_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7269__A2 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8466__A1 net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9278_ _0288_ clknet_leaf_28_i_clk core_0.execute.rf.reg_outputs\[13\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_219_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8229_ _1535_ core_0.execute.alu_mul_div.cbit\[2\] _3846_ _2344_ _3852_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_218_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8029__B _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8769__A2 _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5232__I _1361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_199_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7868__B _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_214_Right_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_198_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8941__A2 _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_2605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_73_i_clk clknet_4_14__leaf_i_clk clknet_leaf_73_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_194_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_85_Right_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8211__C _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_213_3071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xmax_cap219 _1798_ net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_88_i_clk clknet_4_15__leaf_i_clk clknet_leaf_88_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_150_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__A1 _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_2734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_237_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8209__A1 core_0.execute.alu_mul_div.mul_res\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__A4 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7680__A2 _3496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_94_Right_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5691__A1 _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4494__A2 _0675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7432__A2 _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7778__B _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_26_i_clk clknet_4_8__leaf_i_clk clknet_leaf_26_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5930_ core_0.execute.rf.reg_outputs\[9\]\[8\] net224 _1818_ core_0.execute.rf.reg_outputs\[12\]\[8\]
+ _1920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_200_2915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ _1850_ _0836_ _1519_ _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XANTENNA__7196__A1 core_0.execute.sreg_irq_pc.o_d\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7196__B2 core_0.execute.sreg_scratch.o_d\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7600_ _3387_ core_0.ew_data\[14\] _3449_ net26 _3469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__8932__A2 _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_196_2863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4812_ core_0.dec_used_operands\[1\] _0941_ _0992_ core_0.dec_used_operands\[0\]
+ _0993_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_200_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8580_ _2918_ _2949_ _4158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5746__A2 _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6943__A1 _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5792_ core_0.execute.rf.reg_outputs\[1\]\[0\] _1779_ _1781_ core_0.execute.rf.reg_outputs\[10\]\[0\]
+ _1782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_29_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7531_ net29 _1348_ _3412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4743_ core_0.decode.i_flush _0924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_28_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8696__A1 _4249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7462_ core_0.dec_rf_ie\[0\] core_0.ew_reg_ie\[0\] _2419_ _3364_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5745__C _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4674_ net217 net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_113_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9201_ _0212_ clknet_leaf_76_i_clk core_0.ew_data\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_43_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6413_ _2382_ _1004_ _2383_ _1501_ _0163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7018__B core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7393_ _2557_ _2559_ _3312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5317__I _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6171__A2 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9132_ _0144_ clknet_leaf_58_i_clk net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_3_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6344_ core_0.execute.alu_mul_div.div_cur\[12\] _2220_ _2256_ _2320_ _2321_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_11_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9063_ _0088_ clknet_leaf_94_i_clk core_0.fetch.out_buffer_data_pred vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_23_Left_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_228_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7120__A1 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6275_ _2183_ _2248_ _2259_ _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7120__B2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8014_ _3459_ _3695_ _3709_ _0438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5226_ _1358_ net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_228_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7671__A2 _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_60_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5157_ core_0.decode.oc_alu_mode\[9\] _1309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_4_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7423__A2 _3341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5088_ core_0.decode.i_instr_l\[6\] core_0.decode.i_instr_l\[4\] _1245_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input16_I i_core_int_sreg[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__A1 _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6084__S _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8916_ _1231_ _1489_ _4421_ _0628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5985__A2 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8847_ core_0.execute.pc_high_out\[6\] _4369_ _4370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_195_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_238_3369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5198__B1 _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6934__A1 _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8778_ _1729_ _4295_ _4313_ _4307_ _0598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_176_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7729_ core_0.execute.rf.reg_outputs\[11\]\[2\] _3543_ _3539_ _3546_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_2379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8687__A1 net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8231__S0 core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6162__A2 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8439__A1 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5370__B1 _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output84_I net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7662__A2 _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4476__A2 _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_192_Left_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_199_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7598__B _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8611__A1 _3293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7414__A2 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_2675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5976__A2 net322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_230_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_202_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7110__C _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7178__A1 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5028__I1 _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6925__A1 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__A2 _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8678__A1 _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6689__B1 _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7350__A1 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5361__B1 _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5900__A2 _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8448__I _4040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7102__A1 _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8850__A1 _4324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7653__A2 _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6060_ core_0.execute.rf.reg_outputs\[9\]\[7\] net224 _1818_ core_0.execute.rf.reg_outputs\[12\]\[7\]
+ _2050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input8_I i_core_int_sreg[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5664__A1 _1001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__A2 net301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5011_ core_0.fetch.prev_request_pc\[10\] _1151_ _1186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8602__A1 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6962_ _2888_ _2889_ _2890_ _2891_ _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5967__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8701_ _4224_ _4261_ _4249_ _4262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5913_ _1771_ _1900_ _1901_ _1902_ _1903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__7169__A1 _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6893_ core_0.execute.alu_flag_reg.o_d\[2\] _2770_ _2778_ net104 _2825_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__I1 _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8905__A2 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8632_ _0890_ _1704_ _4204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_174_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5844_ _1517_ net179 _1834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_146_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__A2 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4927__B1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8563_ _1685_ core_0.execute.sreg_irq_pc.o_d\[14\] net198 _2134_ _2136_ _4143_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_118_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5775_ _1749_ _1764_ _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__8132__B _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__A2 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7527__I _3408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7514_ _3396_ _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4726_ core_0.execute.pc_high_out\[0\] net104 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8669__A1 _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8494_ _4079_ _4082_ _4083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7971__B _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7445_ _2616_ _3040_ _3355_ _0223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7341__A1 _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6144__A2 _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4657_ core_0.execute.rf.reg_outputs\[5\]\[4\] _0677_ _0686_ core_0.execute.rf.reg_outputs\[14\]\[4\]
+ _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_114_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7892__A2 _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7376_ core_0.execute.alu_mul_div.div_res\[14\] _1742_ _0997_ _3296_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4588_ core_0.execute.rf.reg_outputs\[4\]\[9\] _0720_ net316 core_0.execute.rf.reg_outputs\[8\]\[9\]
+ _0780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9115_ _0127_ clknet_leaf_121_i_clk core_0.execute.alu_mul_div.cbit\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_12_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6327_ core_0.execute.alu_mul_div.div_cur\[10\] _2246_ _2304_ _2305_ _2256_ _2306_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_244_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9046_ _0072_ clknet_leaf_82_i_clk core_0.fetch.prev_request_pc\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__8841__A1 _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7644__A2 _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6258_ core_0.execute.alu_mul_div.div_cur\[3\] _2218_ _2245_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_228_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5655__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5209_ core_0.ew_data\[0\] net156 _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8294__S _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6189_ core_0.execute.alu_mul_div.div_cur\[2\] _2011_ _2075_ core_0.execute.alu_mul_div.div_cur\[3\]
+ _2177_ _2178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_231_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output122_I net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__A2 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6080__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_2408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4630__A2 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_8__f_i_clk_I clknet_3_4_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8042__B _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7881__B _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7332__A1 _2468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6135__A2 core_0.execute.alu_mul_div.mul_res\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_210_3030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8696__C _4209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5894__A1 _1755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_2537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8832__A1 core_0.execute.pc_high_buff_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7635__A2 _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5646__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6843__B1 _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5110__A3 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8060__A2 _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_221_3170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5949__A2 _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8899__A1 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_193_2833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5560_ core_0.fetch.prev_request_pc\[12\] _1082_ _1083_ net163 _1610_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_171_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7791__B _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4511_ _0661_ net263 _0688_ _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__6126__A2 _2115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5491_ net42 _1554_ _1572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7283__S _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7230_ _3153_ _1314_ _2128_ _3154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_123_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4688__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7161_ net85 _2995_ _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_22_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6112_ net95 _1772_ _2096_ _2101_ _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XTAP_TAPCELL_ROW_113_1868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8823__A1 core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7092_ _2075_ _3017_ _3018_ _3019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5637__A1 _1020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6685__I0 _2625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6043_ core_0.execute.rf.reg_outputs\[15\]\[5\] _0944_ _1773_ core_0.execute.rf.reg_outputs\[7\]\[5\]
+ _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_213_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_206_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6426__I net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8051__A2 _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_206_2987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7994_ _3414_ _3694_ _3698_ _0429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6945_ core_0.execute.sreg_long_ptr_en _1692_ _2780_ net10 _2673_ _2876_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_48_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7458__S _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4612__A2 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8641__I _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _2076_ _2104_ _2807_ _1857_ _2808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_124_1997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_rebuffer56_I _1759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_235_3328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5827_ _1814_ _1816_ _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8615_ _4186_ _4187_ _4188_ _4189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_9595_ _0605_ clknet_leaf_62_i_clk core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_91_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7562__A1 _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8546_ _4080_ _3225_ _4128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5758_ net314 net203 _1747_ _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_134_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_153_2349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4709_ net70 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_12
X_8477_ _4047_ _4067_ _4068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6117__A2 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5689_ core_0.dec_sreg_store core_0.execute.sreg_priv_control.o_d\[0\] _1693_ _1694_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_121_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7428_ core_0.ew_data\[15\] _3346_ _2415_ _3347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7865__A2 _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5876__A1 _1760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7206__B _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7359_ _2550_ _2553_ _2483_ _3278_ _3279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_217_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8814__A1 _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7617__A2 _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_246_3479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5628__A1 core_0.decode.i_imm_pass\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9029_ _0056_ clknet_leaf_89_i_clk core_0.fetch.out_buffer_data_instr\[17\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_217_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_2478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8042__A2 _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5240__I _1365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__A1 core_0.execute.rf.reg_outputs\[7\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7553__A1 net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5564__B1 _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7305__A1 net4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6108__A2 _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7305__B2 core_0.execute.sreg_scratch.o_d\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6939__C _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclone94 _0697_ net341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7856__A2 _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7069__B1 _2768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8805__A1 _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7608__A2 _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5095__A2 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4842__A2 net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8033__A2 _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6044__A1 core_0.execute.rf.reg_outputs\[1\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_159_Right_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_203_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8584__A3 _4159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7786__B _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4991_ _1163_ _1165_ _1168_ _1169_ _1080_ net165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__7792__A1 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _2627_ _2660_ _2665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8461__I _4052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_147_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6661_ _2564_ _2585_ _2602_ _1765_ _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_63_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7544__A1 _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8400_ _1974_ _3827_ _3863_ _4011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5612_ _1054_ _1615_ _1641_ _0104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5555__B1 _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9380_ _0390_ clknet_leaf_6_i_clk core_0.execute.rf.reg_outputs\[7\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6592_ _2532_ _2533_ _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8331_ _3927_ _3935_ _3946_ _3947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_60_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ core_0.fetch.prev_request_pc\[4\] _1595_ _1084_ net170 _1601_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__8410__B _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_230_3269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8262_ _1541_ net218 _3883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5474_ core_0.fetch.out_buffer_data_instr\[6\] net65 _1559_ _1562_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7847__A2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5858__A1 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7213_ _2528_ _2531_ _2534_ _3137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8193_ _3814_ _3815_ _3817_ _3818_ _3819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_4_14__f_i_clk_I clknet_3_7_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4530__A1 core_0.execute.rf.reg_outputs\[13\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7144_ net306 _1925_ _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4530__B2 core_0.execute.rf.reg_outputs\[8\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6865__B _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7075_ _1683_ _3001_ _3002_ _3003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6357__S _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6026_ core_0.execute.rf.reg_outputs\[5\]\[4\] net225 net226 core_0.execute.rf.reg_outputs\[10\]\[4\]
+ _1796_ core_0.execute.rf.reg_outputs\[2\]\[4\] _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_146_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6035__A1 net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_126_Right_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_179_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Left_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7696__B _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7977_ core_0.execute.rf.reg_outputs\[5\]\[12\] _3679_ _3677_ _3688_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7783__A1 _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8980__B1 _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4597__A1 net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6928_ _2716_ _2856_ _2858_ _2010_ _2859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_194_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9647_ _0657_ clknet_leaf_139_i_clk core_0.dec_rf_ie\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6859_ _2444_ _2791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6338__A2 _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9578_ _0588_ clknet_leaf_20_i_clk core_0.execute.sreg_scratch.o_d\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8529_ net86 net85 _4099_ _4113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_32_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8320__B _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9421__CLK clknet_leaf_21_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7838__A2 _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6510__A2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_2507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4521__B2 core_0.execute.rf.reg_outputs\[11\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8263__A2 _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_129_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5077__A2 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4824__A2 core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8015__A2 _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6026__A1 core_0.execute.rf.reg_outputs\[5\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6026__B2 core_0.execute.rf.reg_outputs\[10\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7774__A1 core_0.execute.rf.reg_outputs\[10\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4588__A1 core_0.execute.rf.reg_outputs\[4\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_177_2636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__B1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7829__A2 _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_2765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_228_Right_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_239_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5190_ _1247_ _1310_ _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_110_1827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4984__I net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6265__A1 _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7900_ _3460_ _3629_ _3643_ _0390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8006__A2 _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8880_ net202 _4387_ _4397_ _4398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_183_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6017__A1 net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_203_2946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7831_ _3470_ _3586_ _3603_ _0361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_203_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7765__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6568__A2 _2349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4974_ core_0.fetch.prev_request_pc\[12\] _1153_ _1154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_58_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7762_ core_0.execute.rf.reg_outputs\[10\]\[0\] _3564_ _3554_ _3565_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9501_ _0511_ clknet_leaf_125_i_clk core_0.execute.alu_mul_div.mul_res\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6713_ net134 _2642_ _2651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_121_1967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7693_ core_0.execute.rf.reg_outputs\[12\]\[3\] _3521_ _3513_ _3525_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9432_ _0442_ clknet_leaf_137_i_clk core_0.execute.rf.reg_outputs\[4\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6644_ _2009_ _2566_ _2586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_128_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8190__A1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6575_ _2438_ _2490_ _2517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9363_ _0373_ clknet_leaf_7_i_clk core_0.execute.rf.reg_outputs\[8\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_2308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6740__A2 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5526_ net61 _1556_ _1590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8314_ _1538_ _3885_ _3931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4751__A1 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4751__B2 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9294_ _0304_ clknet_leaf_28_i_clk core_0.execute.rf.reg_outputs\[12\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_rebuffer19_I _1833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8245_ _2139_ _3866_ _3867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5457_ _1550_ _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7471__S _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8176_ _2354_ _0999_ _3802_ _3803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5388_ _1437_ _1495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_239_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input46_I i_req_data[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7127_ _2708_ net277 _3054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_243_3427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8245__A2 _3866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_130_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7058_ _2579_ _2573_ _2570_ _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_214_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ net90 _1813_ _1991_ _1998_ _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_214_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_2448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6008__A1 _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7756__A1 _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output202_I net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7508__A1 core_0.ew_reg_ie\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4990__A1 _1016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8181__A1 _1674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_55_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8181__B2 _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6731__A2 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_172_2577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5393__C _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4742__A1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8484__A2 _4048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_237_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6495__A1 _2433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_207_3002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6247__A1 _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9317__CLK clknet_leaf_1_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Left_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_244_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6798__A2 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_218_3131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4981__A1 net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4690_ core_0.execute.rf.reg_outputs\[14\]\[1\] net262 net321 core_0.execute.rf.reg_outputs\[12\]\[1\]
+ _0874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_78_Left_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8172__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_136_2141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6722__A2 _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6399__C _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6360_ net95 _2334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5930__B1 _1818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ _1430_ _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__8387__S _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6291_ _2273_ _2267_ _2187_ _2274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8030_ _3408_ _3715_ _3719_ _0444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5289__A2 net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5242_ _1366_ core_0.ew_mem_width net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_229_3260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8227__A2 _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_87_Left_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5173_ _1279_ _1266_ _1288_ _1322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_71_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7986__A1 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_2281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput1 i_core_int_sreg[0] net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8932_ core_0.dec_mem_we _1286_ _4434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8863_ _2673_ _0901_ _4384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_195_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_210_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7814_ _3441_ _3585_ _3594_ _0353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_176_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8794_ net76 _1738_ _1415_ _4323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_149_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5213__A2 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4957_ net67 core_0.fetch.out_buffer_data_instr\[8\] _0895_ _1137_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_47_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_96_Left_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7745_ core_0.execute.rf.reg_outputs\[11\]\[9\] _3548_ _3554_ _3555_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_191_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6961__A2 _2770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4972__A1 core_0.fetch.prev_request_pc\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4888_ net64 core_0.fetch.out_buffer_data_instr\[5\] _0894_ _1069_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7676_ core_0.execute.rf.reg_outputs\[13\]\[12\] _3504_ _3513_ _3515_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8163__A1 net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9415_ _0425_ clknet_4_1__leaf_i_clk core_0.execute.rf.reg_outputs\[5\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6627_ _1328_ _1757_ _2569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6713__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7910__A1 _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6558_ _2489_ _2491_ _2499_ _2500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
X_9346_ _0356_ clknet_leaf_27_i_clk core_0.execute.rf.reg_outputs\[9\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5509_ _1581_ _0061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8297__S _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6489_ _2428_ _2360_ _2431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9277_ _0287_ clknet_leaf_28_i_clk core_0.execute.rf.reg_outputs\[13\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8466__A2 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8228_ _1535_ core_0.execute.alu_mul_div.cbit\[2\] _2344_ _3846_ _3851_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_2_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8096__I _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9132__D _0144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8159_ net102 _3787_ _3785_ _3793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7977__A1 core_0.execute.rf.reg_outputs\[5\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5988__B1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_7_i_clk clknet_4_2__leaf_i_clk clknet_leaf_7_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_241_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_26_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5204__A2 core_0.ew_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6401__A1 _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7884__B _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_174_2606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4963__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8154__A1 _3440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6704__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4715__A1 net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_213_3072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5912__B1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6468__A1 net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4748__B _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_185_2735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_218_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7417__B1 _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_217_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7968__A1 _3446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5979__B1 _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6640__A1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5579__B _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4651__B1 _0683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_200_2916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ net188 _1850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_158_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7196__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8393__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _0945_ _0946_ _0977_ _0991_ _0992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_158_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_196_2864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _1780_ _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_173_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7530_ net22 _1347_ _3411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4742_ _0900_ _0922_ _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_113_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7461_ _3363_ _0231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4673_ net96 _0667_ _0853_ _0858_ _0859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_154_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9200_ _0211_ clknet_leaf_54_i_clk core_0.ew_data\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6412_ core_0.execute.sreg_data_page _1004_ _2383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4502__I _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4706__A1 _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7392_ _2478_ _2556_ _3311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_43_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6343_ _2221_ _2318_ _2319_ _2224_ _2320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_9131_ _0143_ clknet_leaf_104_i_clk core_0.execute.sreg_priv_control.o_d\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9062_ core_0.fetch.submitable clknet_leaf_106_i_clk core_0.decode.i_submit vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6274_ _2179_ _2259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_116_1899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7120__A2 _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4658__B _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5225_ core_0.ew_data\[0\] core_0.ew_data\[8\] net156 _1358_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6429__I _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8013_ core_0.execute.rf.reg_outputs\[4\]\[11\] _3700_ _3704_ _3709_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_228_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7969__B _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _1308_ _0007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7959__A1 _3420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_208_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5087_ _1232_ _1241_ _1243_ _1244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA_rebuffer86_I net331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6631__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8915_ _1419_ _1286_ _4421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_196_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8846_ core_0.execute.pc_high_out\[5\] core_0.execute.pc_high_out\[4\] _4349_ _4369_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_66_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5198__A1 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8777_ core_0.execute.sreg_scratch.o_d\[14\] _4293_ _4313_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5989_ _1977_ _1978_ _1979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_191_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7728_ _3409_ _3542_ _3545_ _0316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_170_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8136__A1 core_0.ew_reg_ie\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8687__A2 _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8231__S1 core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7659_ _3428_ _3497_ _3505_ _0287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_172_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9329_ _0339_ clknet_leaf_39_i_clk core_0.execute.rf.reg_outputs\[10\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_95_1652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7723__I _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone100_I _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_140_i_clk clknet_4_1__leaf_i_clk clknet_leaf_140_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4568__B _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output77_I net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5122__A1 _1272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput190 net190 sr_bus_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_100_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7879__B _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_155_i_clk clknet_4_0__leaf_i_clk clknet_leaf_155_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8611__A2 _3330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_180_2676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5830__C1 _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8503__B _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8127__A1 _3459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6689__A1 core_0.execute.rf.reg_outputs\[1\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6689__B2 core_0.execute.rf.reg_outputs\[3\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5361__B2 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_108_i_clk clknet_4_12__leaf_i_clk clknet_leaf_108_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7102__A2 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew212 _1853_ net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_237_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_226_3230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ net72 _1185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__6861__A1 _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5664__A2 _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__I net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8602__A2 _3330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_2240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5416__A2 _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6961_ core_0.execute.alu_flag_reg.o_d\[4\] _2770_ _2780_ net11 _2891_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_191_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8700_ net73 _1740_ _1723_ _4261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_177_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5912_ core_0.execute.rf.reg_outputs\[5\]\[9\] _1785_ _1797_ core_0.execute.rf.reg_outputs\[2\]\[9\]
+ _1902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7169__A2 _3085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6892_ net9 _2780_ _2768_ core_0.execute.sreg_scratch.o_d\[2\] _2824_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_192_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8631_ core_0.dec_wfi _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5843_ net313 net194 _1832_ _1833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__8413__B _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7808__I _3584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__B2 _1106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8562_ _4080_ _3297_ _4142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8118__A1 _3446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5774_ _1328_ _1760_ _1764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7513_ core_0.ew_reg_ie\[15\] _3395_ _3396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_133_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4725_ _0903_ _0906_ _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8493_ _4039_ _4081_ _4082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_118_1928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7444_ net127 _3168_ _3355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4656_ core_0.execute.rf.reg_outputs\[2\]\[4\] _0673_ _0710_ core_0.execute.rf.reg_outputs\[8\]\[4\]
+ _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_142_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7341__A2 _3261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput70 i_rst net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__8639__I _4209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5352__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7375_ _1290_ core_0.execute.alu_mul_div.mul_res\[14\] _3294_ core_0.execute.alu_mul_div.i_div
+ _3295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4587_ core_0.execute.rf.reg_outputs\[5\]\[9\] net222 _0679_ core_0.execute.rf.reg_outputs\[11\]\[9\]
+ _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_142_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9114_ _0126_ clknet_leaf_121_i_clk core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6326_ _1547_ _2294_ _2224_ _2305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9045_ core_0.fetch.current_req_branch_pred clknet_leaf_93_i_clk core_0.fetch.prev_req_branch_pred
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6257_ core_0.execute.alu_mul_div.div_cur\[2\] _2220_ _2243_ _2244_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5208_ _1349_ net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6852__A1 _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7699__B _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6188_ _2173_ _2175_ _2176_ _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ core_0.decode.oc_alu_mode\[4\] _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_165_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4615__B1 _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_87_i_clk clknet_4_15__leaf_i_clk clknet_leaf_87_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_output115_I net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6080__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8357__A1 _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_158_2409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8829_ core_0.execute.pc_high_out\[3\] _4327_ _4354_ _4355_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6622__I _2563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_10_i_clk clknet_4_2__leaf_i_clk clknet_leaf_10_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_137_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8109__A1 _3420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5591__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5238__I _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8977__C _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_25_i_clk clknet_4_9__leaf_i_clk clknet_leaf_25_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_210_3031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_169_2538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_219_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7096__A1 _1309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8832__A2 _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__A1 core_0.execute.sreg_irq_pc.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5646__A2 core_0.fetch.dbg_out vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6843__B2 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_42_Left_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7399__A2 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8596__A1 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_3160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_203_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4606__B1 _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__A2 net336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7020__A1 _2759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_193_2823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_2834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4909__A1 core_0.fetch.prev_request_pc\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5582__A1 _1069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Left_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4510_ _0707_ _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_124_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5490_ core_0.fetch.out_buffer_data_instr\[13\] _1571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8520__A1 _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5334__A1 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Right_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7160_ _1683_ core_0.execute.sreg_irq_pc.o_d\[8\] _3086_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_21_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6111_ _2097_ _2098_ _2099_ _2100_ _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_95_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7091_ _2010_ _2863_ _3018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_226_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_107_Right_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6834__A1 _2694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5637__A2 _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6042_ _1771_ _2031_ _2032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_225_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_206_2988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7993_ core_0.execute.rf.reg_outputs\[4\]\[2\] _3695_ _3689_ _3698_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6944_ core_0.execute.pc_high_out\[3\] _2775_ _2768_ core_0.execute.sreg_scratch.o_d\[3\]
+ net80 _1411_ _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__8339__A1 _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__B _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6875_ _2076_ _2042_ _2011_ _2807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8143__B _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_1998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6442__I net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7011__A1 _1759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_235_3329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8614_ _3220_ _3256_ _4188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5826_ core_0.execute.rf.reg_outputs\[13\]\[15\] _1792_ _1815_ core_0.execute.rf.reg_outputs\[9\]\[15\]
+ _1816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_158_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9594_ _0604_ clknet_leaf_40_i_clk core_0.execute.sreg_irq_flags.o_d\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7982__B _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8545_ net74 _4126_ _4127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5573__A1 _1011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5757_ _1518_ net187 _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_146_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4708_ _0890_ net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_8476_ net217 _4048_ _2873_ _2133_ _2874_ _4067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_115_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8511__A1 _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5688_ _1692_ _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_79_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7427_ _2672_ _3344_ _3345_ _3346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5325__A1 _1244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4639_ core_0.execute.rf.reg_outputs\[6\]\[5\] _0670_ net347 core_0.execute.rf.reg_outputs\[15\]\[5\]
+ _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_92_1611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5876__A2 _1865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7358_ _2423_ _2482_ _3278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7078__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6309_ _2221_ _2288_ _2289_ _2246_ _2290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_229_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7289_ _3209_ _2544_ _3210_ _3211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_246_3469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5628__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9028_ _0055_ clknet_leaf_89_i_clk core_0.fetch.out_buffer_data_instr\[16\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_243_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_2479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__A2 _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5800__A2 core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8053__B _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4581__B _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_125_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8750__A1 core_0.execute.sreg_scratch.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5564__B2 net165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_209_Right_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_11_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclone40 _0699_ net321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_106_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8502__A1 _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7305__A2 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclone73 core_0.dec_r_reg_sel\[0\] net301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_180_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7069__A1 net13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7069__B2 core_0.execute.sreg_scratch.o_d\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7132__B _2480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_2043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_141_2210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7241__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6044__A2 _1778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4990_ _1016_ _1146_ _1165_ _1169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7792__A2 _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5587__B _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6660_ _2587_ _2594_ _2601_ _2564_ _2602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_39_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7544__A2 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5611_ core_0.decode.i_imm_pass\[0\] _1616_ _1641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5555__A1 core_0.fetch.prev_request_pc\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5555__B2 net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6591_ _1846_ _2355_ _2533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_144_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_139_2183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8330_ core_0.execute.alu_mul_div.mul_res\[9\] _3933_ _3946_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5542_ _1597_ _1600_ _0075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5307__A1 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _1561_ _0045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8261_ _1541_ _2349_ _3881_ _3882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4510__I _0707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7212_ net276 _2531_ _2534_ _3136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5858__A2 net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8192_ _1674_ net306 _2372_ net234 _1540_ _3818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_10_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7143_ _2006_ _2075_ _3069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__4530__A2 net284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6807__A1 _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7074_ _1683_ core_0.execute.sreg_irq_pc.o_d\[6\] _3002_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_225_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6025_ _1770_ _2012_ _2013_ _2014_ _2015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_198_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7977__B _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_241_3399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7469__S _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7232__A1 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6035__A2 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7976_ _3459_ _3673_ _3687_ _0422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8980__A1 core_0.dec_rf_ie\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7783__A2 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8980__B2 _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6927_ _1896_ _2725_ _2857_ _2858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5794__A1 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4597__A2 _0666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_13__f_i_clk clknet_3_6_0_i_clk clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_9646_ _0656_ clknet_leaf_139_i_clk core_0.dec_rf_ie\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6858_ _2422_ _2789_ _2790_ _0201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7535__A2 _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5546__A1 _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5809_ _1798_ _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_29_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9577_ _0587_ clknet_leaf_19_i_clk core_0.execute.sreg_scratch.o_d\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_146_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6789_ _1898_ _2720_ _2721_ _2722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8528_ _4110_ _4112_ _4051_ _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_162_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7299__A1 _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output182_I net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8459_ _4045_ _4050_ _4051_ _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_107_Left_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_166_2508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4521__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8048__B _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7887__B _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4824__A3 _1001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6026__A2 net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_116_Left_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7774__A2 _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8971__A1 _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5785__A1 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4588__A2 _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_177_2637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7526__A2 core_0.ew_data\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8723__A1 _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__A1 core_0.fetch.prev_request_pc\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5537__B2 net167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9246__CLK clknet_leaf_37_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_125_Left_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9396__CLK clknet_leaf_3_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_192_Right_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_188_2766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_208_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_134_Left_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_162_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7214__A1 _2795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7830_ core_0.execute.rf.reg_outputs\[9\]\[14\] _3584_ _3595_ _3603_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_203_2947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7765__A2 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5776__A1 _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7761_ _3562_ _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__A2 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4973_ core_0.fetch.prev_request_pc\[11\] _1152_ _1153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_199_2895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9500_ _0510_ clknet_4_4__leaf_i_clk core_0.execute.alu_mul_div.mul_res\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6712_ _2646_ _2649_ _2650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4505__I _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7692_ _3415_ _3520_ _3524_ _0301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_1968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8714__A1 core_0.execute.sreg_irq_pc.o_d\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9431_ _0441_ clknet_leaf_144_i_clk core_0.execute.rf.reg_outputs\[4\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6643_ _2568_ _2577_ _2584_ _2585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_46_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8190__A2 _2155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_143_Left_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_9362_ _0372_ clknet_leaf_27_i_clk core_0.execute.rf.reg_outputs\[8\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6574_ _2439_ _2488_ _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_171_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6740__A3 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_2309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8313_ _3903_ _3929_ _3878_ _3930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5525_ _1589_ _0069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9293_ _0303_ clknet_leaf_28_i_clk core_0.execute.rf.reg_outputs\[12\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8244_ net218 _2090_ _2102_ _2115_ core_0.execute.alu_mul_div.cbit\[0\] core_0.execute.alu_mul_div.cbit\[1\]
+ _3866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_5456_ _1008_ _1549_ _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_67_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8647__I _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4503__A2 _0698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8175_ _3801_ _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5387_ _1489_ _1493_ _1494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_100_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _2711_ _3040_ _3050_ _3052_ _3053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_10_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_243_3428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input39_I i_req_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7453__A1 _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_5_0_i_clk clknet_0_i_clk clknet_3_5_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7057_ _1880_ _2438_ _2978_ _2980_ _2984_ _2985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_241_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6008_ _1813_ _1992_ _1997_ _1998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_241_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_2449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7205__A1 _2708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8315__C _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7756__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5767__A1 _1755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7959_ _3420_ _3672_ _3678_ _0414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7508__A2 core_0.ew_reg_ie\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9629_ _0639_ clknet_leaf_114_i_clk net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_135_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6716__B1 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4990__A2 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8181__A2 _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_21_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_2578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4742__A2 _0922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5246__I _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_1694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7692__A1 _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_217_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7995__A2 _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8244__I0 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7747__A2 _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5758__A1 net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_218_3132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6707__B1 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4981__A2 _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4733__A2 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5310_ _0891_ _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6290_ _2167_ _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7683__A1 _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6486__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5241_ core_0.ew_addr\[0\] _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_229_3261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6891__C1 _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5172_ _1232_ _1320_ _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7435__A1 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6238__A2 _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_2271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7986__A2 _3394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_2282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput2 i_core_int_sreg[10] net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8931_ _4433_ _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8862_ _1419_ _2771_ _4383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_78_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8935__A1 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7738__A2 _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7813_ core_0.execute.rf.reg_outputs\[9\]\[6\] _3591_ _3580_ _3594_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5749__A1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8793_ _0901_ _4322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6946__B1 _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7744_ _3512_ _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4956_ net39 core_0.fetch.out_buffer_data_instr\[10\] _0894_ _1136_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7675_ _3460_ _3498_ _3514_ _0294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8151__B _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4887_ net65 core_0.fetch.out_buffer_data_instr\[6\] _0893_ _1068_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8163__A2 _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9414_ _0424_ clknet_leaf_24_i_clk core_0.execute.rf.reg_outputs\[5\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6626_ _2567_ _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_117_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer31_I _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7910__A2 _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9345_ _0355_ clknet_leaf_31_i_clk core_0.execute.rf.reg_outputs\[9\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4724__A2 _0904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6557_ _2494_ _2497_ _2498_ _2499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5921__A1 net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5066__I _0904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5508_ core_0.fetch.out_buffer_data_instr\[22\] net51 _1559_ _1581_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9276_ _0286_ clknet_leaf_8_i_clk core_0.execute.rf.reg_outputs\[13\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6488_ _1843_ net214 _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8466__A3 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8227_ _3802_ _3832_ _3849_ _3850_ _0510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__7674__A1 core_0.execute.rf.reg_outputs\[13\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5524__I1 net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5439_ core_0.execute.alu_mul_div.comp _1001_ _1533_ _0923_ _1534_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_246_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8158_ _3450_ _3780_ _3792_ _0499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_227_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7426__A1 core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ _1290_ core_0.execute.alu_mul_div.mul_res\[7\] _3036_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8089_ _3459_ _3738_ _3752_ _0470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7977__A2 _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5988__B2 core_0.execute.rf.reg_outputs\[9\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7230__B _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7729__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8926__A1 _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_239_Left_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_46_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__A2 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8154__A2 _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6360__I net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7901__A2 _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__A1 core_0.execute.rf.reg_outputs\[5\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5912__B2 core_0.execute.rf.reg_outputs\[2\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_213_3073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__B1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6468__A2 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7665__A1 _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_2736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_218_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9434__CLK clknet_leaf_37_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7417__B2 core_0.execute.sreg_scratch.o_d\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5640__S _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7968__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5979__B2 core_0.execute.rf.reg_outputs\[10\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8917__A1 core_0.dec_sreg_load vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9584__CLK clknet_leaf_108_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4651__B2 core_0.execute.rf.reg_outputs\[7\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_200_2917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7440__I1 _2954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4810_ _0981_ _0984_ _0987_ _0990_ _0991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_185_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_196_2865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _0971_ core_0.dec_l_reg_sel\[2\] _0953_ core_0.dec_l_reg_sel\[0\] _1780_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_145_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4741_ _0907_ _0910_ _0921_ _0922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_29_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7460_ net120 _3335_ _2415_ _3363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6156__A1 _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4672_ _0854_ _0855_ _0856_ _0857_ _0858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_114_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6411_ net103 _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7391_ _2839_ _3309_ _3310_ _0214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_153_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9130_ _0142_ clknet_leaf_106_i_clk core_0.execute.sreg_priv_control.o_d\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6342_ _2141_ _2311_ _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7656__A1 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7315__B core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9061_ _0087_ clknet_leaf_91_i_clk core_0.fetch.prev_request_pc\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6273_ _2254_ _2257_ _2258_ _0148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_149_2300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8012_ _3456_ _3695_ _3708_ _0437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5224_ _1357_ net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_209_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7408__A1 _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5155_ _1292_ _1251_ _1293_ _1307_ _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7959__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8081__A1 _3446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5086_ _1242_ core_0.decode.i_instr_l\[2\] _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_224_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8146__B _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_98_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6631__A2 _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8914_ _4419_ _4420_ _0627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_196_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8908__A1 _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer79_I _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8845_ _4316_ _4368_ _0610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_149_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7477__S _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8384__A2 _3995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_1__f_i_clk clknet_3_0_0_i_clk clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_149_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6395__A1 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5198__A2 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8776_ _1726_ _4295_ _4312_ _4307_ _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5988_ core_0.execute.rf.reg_outputs\[13\]\[13\] _1792_ _1815_ core_0.execute.rf.reg_outputs\[9\]\[13\]
+ _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7727_ core_0.execute.rf.reg_outputs\[11\]\[1\] _3543_ _3539_ _3545_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4939_ _1107_ _1118_ _1119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7276__I _3198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8136__A2 _3394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6147__A1 _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7658_ core_0.execute.rf.reg_outputs\[13\]\[4\] _3504_ _3500_ _3505_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7344__B1 _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7895__A1 core_0.execute.rf.reg_outputs\[7\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6609_ _2548_ _2551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_160_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7589_ core_0.execute.rf.reg_outputs\[15\]\[11\] _3429_ _3422_ _3461_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9328_ _0338_ clknet_leaf_39_i_clk core_0.execute.rf.reg_outputs\[10\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5370__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9259_ _0269_ clknet_leaf_1_i_clk core_0.execute.rf.reg_outputs\[14\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A2 _1276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput180 net180 sr_bus_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput191 net191 sr_bus_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_215_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4881__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_2677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4633__A1 core_0.execute.rf.reg_outputs\[15\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5830__B1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_230_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7895__B _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8127__A2 _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6689__A2 _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7638__A1 _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7489__I1 core_0.ew_reg_ie\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_3220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4872__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_144_2241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6074__B1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7810__A1 _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6960_ core_0.execute.sreg_priv_control.o_d\[4\] _1692_ _2768_ core_0.execute.sreg_scratch.o_d\[4\]
+ _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_108_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5821__B1 _1783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5911_ core_0.execute.rf.reg_outputs\[13\]\[9\] _1792_ _1901_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_221_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6891_ core_0.execute.pc_high_buff_out\[2\] _2771_ _2774_ core_0.execute.sreg_irq_pc.o_d\[2\]
+ _2775_ core_0.execute.pc_high_out\[2\] _2823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_177_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clone39_A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8630_ _4201_ _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_186_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6377__A1 _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ _1517_ net178 _1832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_57_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_237_3360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8561_ net76 _4133_ _4141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4927__A2 _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5773_ net255 _1762_ _1763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__8118__A2 _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7512_ _3394_ _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_127_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4724_ core_0.execute.prev_pc_high\[2\] _0904_ _0905_ core_0.execute.prev_pc_high\[1\]
+ _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6129__A1 _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8492_ _1685_ core_0.execute.sreg_irq_pc.o_d\[5\] net204 _2134_ _2954_ _4080_ _4081_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_127_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7443_ _2616_ _2994_ _3354_ _0222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7877__A1 core_0.execute.rf.reg_outputs\[7\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_2370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4655_ core_0.execute.rf.reg_outputs\[1\]\[4\] _0693_ _0703_ core_0.execute.rf.reg_outputs\[15\]\[4\]
+ _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_142_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput60 i_req_data[30] net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_6_i_clk clknet_4_2__leaf_i_clk clknet_leaf_6_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5352__A2 _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7374_ _2124_ _3293_ _3294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4586_ core_0.execute.rf.reg_outputs\[10\]\[9\] net221 net220 core_0.execute.rf.reg_outputs\[9\]\[9\]
+ _0778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_9_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9113_ _0003_ clknet_leaf_110_i_clk core_0.decode.oc_alu_mode\[13\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6325_ _2221_ _2303_ _2304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9044_ _0071_ clknet_leaf_91_i_clk core_0.fetch.out_buffer_valid vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6256_ _2241_ _2242_ _2224_ _2243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5207_ _1348_ _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__8655__I _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6187_ core_0.execute.alu_mul_div.div_cur\[2\] _2008_ _2176_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_90_1594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8054__A1 _3462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5138_ _1230_ _1256_ _1289_ _1291_ _0011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_input21_I i_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7801__A1 _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5069_ _0914_ net113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_211_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4615__A1 core_0.execute.rf.reg_outputs\[7\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4615__B2 core_0.execute.rf.reg_outputs\[3\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8604__B _3329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8828_ net217 _4328_ _4326_ _4353_ _4354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_183_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8759_ core_0.execute.sreg_scratch.o_d\[6\] _4300_ _4303_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5040__A1 _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8109__A2 _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5591__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7868__A1 core_0.execute.rf.reg_outputs\[8\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_210_3032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4551__B1 _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5894__A3 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_2539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8293__A1 _2054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__A2 _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_121_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8045__A1 _3450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_203_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6085__I _2074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_221_3161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6359__A1 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7020__A2 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_2824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4909__A2 _1026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_214_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5582__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_46_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6906__I0 core_0.ew_data\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4542__B1 _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ core_0.execute.rf.reg_outputs\[7\]\[2\] _1821_ _1785_ core_0.execute.rf.reg_outputs\[5\]\[2\]
+ _2100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_186_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8284__A1 _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7090_ _1751_ _2858_ _3017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_237_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__A2 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6041_ core_0.execute.rf.reg_outputs\[6\]\[5\] net219 _1819_ core_0.execute.rf.reg_outputs\[12\]\[5\]
+ _1787_ core_0.execute.rf.reg_outputs\[3\]\[5\] _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_119_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4845__A1 _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8036__A1 core_0.execute.rf.reg_outputs\[3\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7992_ _3408_ _3694_ _3697_ _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_68_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_206_2989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6943_ _1401_ core_0.execute.sreg_irq_pc.o_d\[3\] _2874_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6874_ _1930_ _1927_ _2805_ _2806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_193_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_1999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7011__A2 _2939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8613_ _3188_ _3150_ _4187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5825_ net340 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_146_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9593_ _0603_ clknet_leaf_63_i_clk core_0.execute.sreg_irq_flags.o_d\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5022__A1 core_0.fetch.prev_request_pc\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8544_ net73 _4121_ _4126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5756_ core_0.dec_r_bus_imm _1746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_146_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6770__A1 _2130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5573__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4707_ net87 _0667_ _0885_ _0889_ _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_162_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8475_ _4039_ _4065_ _4066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5687_ _1686_ _1689_ _1691_ _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xclkbuf_leaf_154_i_clk clknet_4_0__leaf_i_clk clknet_leaf_154_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7426_ core_0.dec_mem_access net232 _3345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6522__A1 net247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4638_ core_0.execute.rf.reg_outputs\[11\]\[5\] net303 net257 core_0.execute.rf.reg_outputs\[8\]\[5\]
+ _0826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_input69_I i_req_data_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7357_ _2423_ _2476_ _3276_ _3277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_102_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5074__I _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4569_ _0759_ _0760_ _0761_ _0762_ _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_229_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8275__A1 core_0.execute.alu_mul_div.mul_res\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _2141_ _2280_ _2289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_228_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7288_ _3209_ _2544_ _1326_ _3210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_246_3459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9027_ _0054_ clknet_leaf_102_i_clk core_0.fetch.out_buffer_data_instr\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_217_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6239_ core_0.decode.o_submit _0998_ _2228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5802__I _1791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8027__A1 _3401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_107_i_clk clknet_4_12__leaf_i_clk clknet_leaf_107_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_137_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5249__I _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5013__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8750__A2 _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5564__A2 _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6761__A1 _2691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_173_Right_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclone30 _0719_ net318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_11_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclone41 net337 net322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_118_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclone74 _0692_ net302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_152_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_189_Left_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7069__A2 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8266__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_235_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9175__CLK clknet_leaf_42_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8018__A1 _3465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8569__A2 _4048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7241__A2 _3155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__B _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_198_Left_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__C net293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5610_ _1638_ _1640_ _0103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8741__A2 _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5555__A2 _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6590_ _2464_ _2532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_27_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_71_i_clk clknet_4_12__leaf_i_clk clknet_leaf_71_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_140_Right_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4998__I net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5541_ core_0.fetch.prev_request_pc\[3\] _1595_ _1084_ net169 _1600_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_60_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_152_2340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8260_ _1541_ _2102_ _3881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5472_ core_0.fetch.out_buffer_data_instr\[5\] net64 _1559_ _1561_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_170_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6504__A1 _1755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7211_ _2480_ _3134_ _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_86_i_clk clknet_4_15__leaf_i_clk clknet_leaf_86_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8191_ _2354_ _1835_ _3816_ _1545_ _3817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_22_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7142_ _3065_ _2526_ _2795_ _3068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8419__B _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6807__A2 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7323__B _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7073_ net83 _2995_ _3000_ _2893_ _3001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_226_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4818__A1 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8009__A1 core_0.execute.rf.reg_outputs\[4\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ core_0.execute.rf.reg_outputs\[13\]\[4\] _1791_ net331 core_0.execute.rf.reg_outputs\[4\]\[4\]
+ _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_226_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5491__A1 net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7975_ core_0.execute.rf.reg_outputs\[5\]\[11\] _3679_ _3677_ _3687_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_24_i_clk clknet_4_9__leaf_i_clk clknet_leaf_24_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7549__I _3427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8980__A2 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6926_ _1930_ _2715_ _2857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_221_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_rebuffer61_I net288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5794__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7993__B _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ core_0.ew_data\[1\] _2642_ _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9645_ _0655_ clknet_leaf_139_i_clk core_0.dec_rf_ie\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5069__I _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_202_Left_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7485__S _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8732__A2 _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5808_ _0942_ _0947_ _0954_ _0955_ _1798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_39_i_clk clknet_4_8__leaf_i_clk clknet_leaf_39_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_9576_ _0586_ clknet_leaf_19_i_clk core_0.execute.sreg_scratch.o_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5546__A2 _1602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6788_ _1899_ _1942_ _2721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_1_0_i_clk clknet_0_i_clk clknet_3_1_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_162_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8527_ _4047_ _4111_ _4112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5739_ core_0.execute.sreg_priv_control.o_d\[14\] _1700_ _1730_ _1697_ _1731_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_150_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7299__A2 core_0.execute.alu_mul_div.mul_res\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8496__A1 net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8458_ _1702_ _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7217__C _2563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7409_ _2564_ _3326_ _3327_ _3063_ _3328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA_output175_I net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8389_ core_0.execute.alu_mul_div.mul_res\[15\] _4000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_166_2509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_211_Left_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__A1 _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__A4 _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_242_Right_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8420__A1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8064__B _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_240_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8971__A2 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6982__A1 net325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5785__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_220_Left_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_177_2638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8184__B1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__A2 _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4611__I _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8487__A1 _1211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8239__A1 _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_188_2767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6538__I core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8954__S _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5442__I _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_222_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8411__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_203_2948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7760_ _3562_ _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_230_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4972_ core_0.fetch.prev_request_pc\[10\] _1151_ _1152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_188_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5776__A2 core_0.decode.oc_alu_mode\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_199_2896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6711_ _2647_ _2648_ _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7691_ core_0.execute.rf.reg_outputs\[12\]\[2\] _3521_ _3513_ _3524_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_121_1969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8714__A2 _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9430_ _0440_ clknet_leaf_144_i_clk core_0.execute.rf.reg_outputs\[4\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6642_ _2568_ _2583_ _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9361_ _0371_ clknet_leaf_29_i_clk core_0.execute.rf.reg_outputs\[8\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6573_ _2502_ _2511_ _2513_ _2514_ _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_26_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8312_ _1668_ net213 _3928_ _3929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5524_ core_0.fetch.out_buffer_data_instr\[30\] net60 _1550_ _1589_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6740__A4 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9292_ _0302_ clknet_leaf_8_i_clk core_0.execute.rf.reg_outputs\[12\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9340__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8243_ _3853_ _3857_ _3864_ _3865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5455_ _0891_ _0896_ _1367_ _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_41_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7150__A1 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6876__C _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8174_ core_0.decode.o_submit _1743_ _3801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_100_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5386_ _1282_ _1301_ _1491_ _1492_ _1493_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__8149__B _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7125_ _2711_ _3051_ _3052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7053__B _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9490__CLK clknet_leaf_21_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_243_3429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_238_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7453__A2 _3192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7056_ net214 _1889_ _2981_ net260 _2983_ _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_157_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6007_ core_0.execute.rf.reg_outputs\[15\]\[12\] _0945_ _1821_ core_0.execute.rf.reg_outputs\[7\]\[12\]
+ _1996_ _1997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_214_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_161_2439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8953__A2 _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7958_ core_0.execute.rf.reg_outputs\[5\]\[3\] _3673_ _3677_ _3678_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6964__A1 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5767__A2 _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6964__B2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6909_ _1329_ _2740_ _2737_ _2840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_166_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_194_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7889_ core_0.execute.rf.reg_outputs\[7\]\[6\] _3634_ _3636_ _3638_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8705__A2 _4209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7508__A3 core_0.ew_reg_ie\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5519__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9628_ _0638_ clknet_leaf_94_i_clk net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6716__A1 core_0.execute.rf.reg_outputs\[7\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__B2 core_0.execute.rf.reg_outputs\[5\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9559_ _0569_ clknet_leaf_75_i_clk core_0.execute.sreg_irq_pc.o_d\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_21_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8469__A1 _1738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_172_2579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_1684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7692__A2 _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8059__B _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7444__A2 _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5455__A1 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_220_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8244__I1 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__B1 _2375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6955__A1 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5758__A2 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_1791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_218_3133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6707__A1 core_0.execute.rf.reg_outputs\[7\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6707__B2 core_0.execute.rf.reg_outputs\[5\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9363__CLK clknet_leaf_7_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_136_2143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5930__A2 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _1365_ net144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_228_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8880__A1 net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7683__A2 _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_229_3262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6891__B1 _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Right_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5171_ _1233_ _1236_ _1269_ _1320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_236_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_194_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7435__A2 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8632__A1 _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_2272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8930_ _1431_ _4432_ _4433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput3 i_core_int_sreg[11] net3 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8861_ _4376_ _4327_ _4382_ _1431_ _0612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7199__A1 net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7199__B2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5121__B _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8935__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4516__I _0713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7812_ _3435_ _3585_ _3593_ _0352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8792_ _4316_ _4321_ _0604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_188_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5749__A2 _1738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6946__A1 core_0.execute.pc_high_buff_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7743_ _3451_ _3542_ _3553_ _0323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4955_ net68 core_0.fetch.out_buffer_data_instr\[9\] _0894_ _1135_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_27_Right_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8699__A1 _4219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7674_ core_0.execute.rf.reg_outputs\[13\]\[11\] _3504_ _3513_ _3514_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4886_ _1015_ _1066_ _1067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_82_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9413_ _0423_ clknet_leaf_35_i_clk core_0.execute.rf.reg_outputs\[5\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6625_ _1751_ _2566_ _2567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_74_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5347__I _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7371__A1 _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_94_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6556_ _2453_ _2493_ _2498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9344_ _0354_ clknet_leaf_30_i_clk core_0.execute.rf.reg_outputs\[9\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_rebuffer24_I net251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5921__A2 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5507_ _1580_ _0060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6379__S _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9275_ _0285_ clknet_leaf_5_i_clk core_0.execute.rf.reg_outputs\[13\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6487_ _2428_ _2360_ _2429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8226_ _3802_ _2740_ _3830_ core_0.execute.alu_mul_div.mul_res\[2\] _3850_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_112_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8871__A1 _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7674__A2 _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5438_ core_0.decode.i_flush net70 _1533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_36_Right_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input51_I i_req_data[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8157_ net101 _3787_ _3785_ _3792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5369_ _1439_ core_0.decode.i_instr_l\[8\] core_0.decode.i_instr_l\[7\] _1480_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7108_ _3013_ _3016_ _3027_ _3034_ _3035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__8623__A1 core_0.execute.alu_flag_reg.o_d\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8088_ core_0.execute.rf.reg_outputs\[2\]\[11\] _3743_ _3745_ _3752_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_214_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7511__B _3393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7039_ core_0.ew_data\[5\] _2967_ _0199_ _2968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5988__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8326__C _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Right_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6937__A1 _2759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9386__CLK clknet_leaf_1_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_46_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5373__B1 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_213_3063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5912__A2 _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_213_3074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7114__A1 core_0.execute.sreg_priv_control.o_d\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7114__B2 net14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Right_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8862__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7665__A2 _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5676__A1 _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_2737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7417__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8614__A1 _3220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5428__A1 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8090__A2 _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A2 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Right_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4651__A2 _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8917__A2 _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_200_2907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_200_2918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7647__I _3496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_196_2866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5600__A1 _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4740_ _0916_ _0920_ _0921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_116_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4671_ core_0.execute.rf.reg_outputs\[11\]\[3\] net303 _0716_ _0857_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7353__A1 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5167__I core_0.execute.alu_mul_div.i_mod vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6156__A2 _0713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6410_ _2381_ _0162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7390_ core_0.ew_data\[14\] _3168_ _3310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5364__B1 _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_72_Right_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6341_ _2150_ _2317_ _2318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9060_ _0086_ clknet_leaf_89_i_clk core_0.fetch.prev_request_pc\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8853__A1 _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7656__A2 _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6272_ _2229_ _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_12_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_2301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5667__A1 _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9259__CLK clknet_leaf_1_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8011_ core_0.execute.rf.reg_outputs\[4\]\[10\] _3700_ _3704_ _3708_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_121_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5223_ core_0.ew_data\[7\] net156 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8605__A1 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5154_ _1300_ _1304_ _1305_ _1306_ _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__8427__B _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5085_ core_0.decode.i_instr_l\[3\] _1242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__8081__A2 _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_81_Right_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_223_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6092__B2 core_0.execute.rf.reg_outputs\[5\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7050__C _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8913_ _1293_ _1267_ _1274_ _4420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_78_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8908__A2 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8844_ core_0.execute.pc_high_out\[5\] _4327_ _4367_ _4368_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5987_ core_0.execute.rf.reg_outputs\[8\]\[13\] _1794_ _1776_ core_0.execute.rf.reg_outputs\[4\]\[13\]
+ _1977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8775_ core_0.execute.sreg_scratch.o_d\[13\] _4300_ _4312_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7557__I _3434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4938_ _1108_ _1117_ _1118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7726_ _3402_ _3542_ _3544_ _0315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4869_ _1043_ _1046_ _1049_ _1050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7344__A1 core_0.execute.sreg_irq_pc.o_d\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6147__A2 _2134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7657_ _3496_ _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7344__B2 core_0.execute.sreg_scratch.o_d\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7493__S _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_90_Right_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6608_ _2538_ _2542_ _2545_ _2549_ _2550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_6_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7895__A2 _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7588_ _3459_ _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_43_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9327_ _0337_ clknet_leaf_40_i_clk core_0.execute.rf.reg_outputs\[10\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6539_ net212 _1974_ _2480_ _2481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_95_1654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9258_ _0268_ clknet_leaf_1_i_clk core_0.execute.rf.reg_outputs\[14\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5658__A1 _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5026__B core_0.fetch.prev_request_pc\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8209_ core_0.execute.alu_mul_div.mul_res\[0\] _3823_ _3824_ _3834_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xoutput170 net170 o_req_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9189_ _0200_ clknet_leaf_53_i_clk core_0.ew_data\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_219_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput181 net181 sr_bus_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput192 net192 sr_bus_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_199_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6083__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_2667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_2678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4633__A2 _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5830__A1 core_0.execute.rf.reg_outputs\[6\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_161_Left_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6386__A2 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7583__B2 net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_194_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7335__A1 _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__A1 core_0.decode.oc_alu_mode\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_170_Left_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5715__I _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8835__A1 net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7638__A2 _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6846__B1 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A2 _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_226_3221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8962__S _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_42_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5450__I _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_2242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6074__A1 core_0.execute.rf.reg_outputs\[14\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7271__B1 _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7810__A2 _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A1 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5821__B2 _1810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_187_Right_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5910_ core_0.execute.rf.reg_outputs\[7\]\[9\] _1821_ _1900_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6890_ core_0.execute.sreg_irq_pc.o_d\[2\] _2822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_88_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone39_A2 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ net313 net196 _1830_ _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_220_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6377__A2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8560_ _4053_ _4139_ _4140_ _1702_ _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5772_ _1328_ _1761_ _1762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_237_3361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4723_ core_0.execute.pc_high_out\[1\] _0901_ _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_29_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7511_ _3386_ _3388_ _3393_ _3394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_8491_ _1419_ _1685_ _4080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_44_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6129__A2 _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7442_ net126 _3168_ _3354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7877__A2 _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4654_ _0837_ _0838_ _0839_ _0840_ _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_155_2371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput50 i_req_data[21] net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput61 i_req_data[31] net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7373_ _3277_ _3282_ _3287_ _3292_ _3293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_3_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4585_ _0777_ net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__5352__A3 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9112_ _0002_ clknet_leaf_127_i_clk core_0.decode.oc_alu_mode\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6324_ _2163_ _2302_ _2303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7629__A2 _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9043_ _0070_ clknet_leaf_90_i_clk core_0.fetch.out_buffer_data_instr\[31\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6255_ _1546_ _2233_ _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6301__A2 _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5206_ _1347_ _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
X_6186_ _2170_ _2174_ _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_243_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8157__B _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_1595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8054__A2 _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5137_ _1290_ _1286_ _1291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6456__I net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer91_I _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6065__A1 _1757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5068_ _0917_ net112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7801__A2 _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input14_I i_core_int_sreg[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4615__A2 net297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_154_Right_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8827_ _4324_ _4352_ _4353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7565__A1 core_0.execute.rf.reg_outputs\[15\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_0_Right_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_176_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8758_ _0836_ _4294_ _4302_ _4287_ _0589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5040__A2 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7709_ core_0.execute.rf.reg_outputs\[12\]\[10\] _3526_ _3528_ _3534_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7317__A1 core_0.ew_data\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8689_ _4224_ _4250_ _4251_ _4249_ _4252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_62_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7868__A2 _3605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__A1 _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_160_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_210_3033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__A2 _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__A3 _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8817__A1 core_0.execute.pc_high_buff_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4551__A1 core_0.execute.rf.reg_outputs\[5\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4551__B2 core_0.execute.rf.reg_outputs\[4\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output82_I net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8293__A2 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_235_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8045__A2 _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6056__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4606__A2 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5803__A1 _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_221_3162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_121_Right_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_159_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_2825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7308__A1 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7308__B2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5873__C _1862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7859__A2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_232_3291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5445__I _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6531__A2 _2371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8808__A1 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6477__S _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8284__A2 _2054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6295__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6040_ _2028_ _2029_ _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_238_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_237_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input6_I i_core_int_sreg[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4845__A2 net58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8036__A2 _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7795__A1 core_0.execute.rf.reg_outputs\[10\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7991_ core_0.execute.rf.reg_outputs\[4\]\[1\] _3695_ _3689_ _3697_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_206_2979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6942_ core_0.execute.alu_mul_div.div_cur\[3\] _1317_ _2870_ _2872_ _2873_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_88_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7547__A1 _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6873_ _1898_ _1930_ _2055_ _2070_ _2805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_88_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9447__CLK clknet_leaf_145_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8612_ _3079_ _3115_ _4186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_157_2400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5558__B1 _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5824_ core_0.execute.rf.reg_outputs\[8\]\[15\] _1794_ _1776_ core_0.execute.rf.reg_outputs\[4\]\[15\]
+ _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_147_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9592_ _0602_ clknet_leaf_40_i_clk core_0.execute.sreg_irq_flags.o_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8543_ _4053_ _4124_ _4125_ _4051_ _0551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_173_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5755_ _1519_ net253 _1744_ _1745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_60_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6770__A2 _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7835__I _3605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ _0667_ _0886_ _0887_ _0888_ _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_8474_ _4041_ _4063_ _4064_ _4065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5686_ _1690_ net177 _1421_ _1691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_44_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7425_ _2703_ _3335_ _3343_ _3344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_60_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4637_ _0825_ net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_142_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6522__A2 _1941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7356_ _2423_ _2476_ _1292_ _3276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4568_ core_0.execute.rf.reg_outputs\[15\]\[11\] _0702_ _0715_ _0762_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_92_1613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ _2160_ _2287_ _2288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7287_ _2538_ _2542_ _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_12_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4499_ _0671_ _0678_ _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__6286__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_223_Right_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6238_ core_0.execute.alu_mul_div.div_cur\[1\] _2218_ _2227_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9026_ _0053_ clknet_leaf_102_i_clk core_0.fetch.out_buffer_data_instr\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_244_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8027__A2 _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6169_ core_0.execute.alu_mul_div.div_cur\[8\] net306 _2158_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_243_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output120_I net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8735__B1 _1418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5549__B1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5013__A2 net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6761__A2 _2692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclone42 _1863_ net270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_11_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone75 _0679_ net303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_105_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5265__I core_0.execute.alu_flag_reg.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7710__A1 _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4524__A1 core_0.execute.rf.reg_outputs\[4\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_239_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8266__A2 _3886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7413__C _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_234_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8018__A2 _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6029__A1 core_0.execute.rf.reg_outputs\[15\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7777__A1 _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_5_i_clk clknet_4_2__leaf_i_clk clknet_leaf_5_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7529__A1 _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6201__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_234_3320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8741__A3 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5540_ _1597_ _1599_ _0074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4763__A1 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5960__B1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5471_ _1560_ _0044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_170_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_2341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7701__A1 core_0.execute.rf.reg_outputs\[12\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7210_ _2459_ _2463_ _2532_ _3134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4515__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4515__B2 _0712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8190_ _2354_ _2155_ _3816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7141_ _3066_ _3067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6268__A1 _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7072_ _2997_ _2998_ _2999_ _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_4_7__f_i_clk_I clknet_3_3_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4818__A2 _0998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6023_ core_0.execute.rf.reg_outputs\[8\]\[4\] net345 _2013_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8009__A2 _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4519__I _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5491__A2 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8435__B _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_163_2470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7974_ _3456_ _3673_ _3686_ _0421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_221_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6925_ _2009_ _2565_ _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_221_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9644_ _0654_ clknet_leaf_66_i_clk core_0.dec_jump_cond_code\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6856_ _2709_ net200 _2788_ _2789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5807_ _1796_ _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__8170__B _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9575_ _0585_ clknet_leaf_19_i_clk core_0.execute.sreg_scratch.o_d\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6787_ _1875_ net213 _2720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7940__A1 core_0.execute.rf.reg_outputs\[6\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6743__A2 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8526_ _0789_ _4048_ _3120_ _2133_ _3125_ _4111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_91_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5738_ _1729_ _1704_ _1730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8496__A2 _4076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8457_ _4047_ _4049_ _4050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ _1671_ _1675_ _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_5_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4506__A1 _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7408_ _2564_ _3033_ _3327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8388_ _3999_ _0522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output168_I net168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7339_ core_0.execute.alu_mul_div.div_cur\[13\] _2128_ _3260_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6259__A1 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4809__A2 _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9009_ _0036_ clknet_leaf_111_i_clk core_0.dec_r_bus_imm vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_216_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7759__A1 core_0.ew_reg_ie\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__B1 net321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_89_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8420__A2 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6431__A1 _1211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8971__A3 _1272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6982__A2 _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5785__A3 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_2639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4993__A1 core_0.fetch.prev_request_pc\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8184__A1 _1674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8080__B _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5942__B1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__A1 _2438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Left_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5170__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_2768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9292__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6670__A1 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4681__B1 _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_153_i_clk clknet_4_0__leaf_i_clk clknet_leaf_153_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8411__A2 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_3390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_203_2949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ core_0.fetch.prev_request_pc\[9\] core_0.fetch.prev_request_pc\[8\] _1150_
+ _1151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_48_Left_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_176_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6710_ _2627_ _2634_ _2640_ _2648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_199_2897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7690_ _3409_ _3520_ _3523_ _0300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_132_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_1959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8702__C _4209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6641_ _2579_ _2581_ _2582_ _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_184_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6725__A2 _2654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer4_I net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9360_ _0370_ clknet_leaf_30_i_clk core_0.execute.rf.reg_outputs\[8\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _2489_ _2491_ _2514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_41_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8311_ _1668_ _2521_ _3928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5523_ _1024_ _1552_ _1588_ _0068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9291_ _0301_ clknet_leaf_5_i_clk core_0.execute.rf.reg_outputs\[12\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6489__A1 _2428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8242_ core_0.execute.alu_mul_div.mul_res\[3\] _3856_ _3864_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5454_ _1534_ _1548_ _0039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5161__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5385_ _1267_ _1331_ _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8173_ _3472_ _3781_ _3800_ _0506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_239_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7124_ _3004_ _3049_ _3051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_106_i_clk clknet_4_12__leaf_i_clk clknet_leaf_106_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7055_ _1885_ _2982_ _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6110__B1 _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8650__A2 _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clone74_I _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6661__A1 _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _1993_ _1994_ _1995_ _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_207_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8165__B _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_90_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_206_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8402__A2 _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7957_ _3647_ _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6964__A2 _2829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6908_ _2421_ _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4975__A1 core_0.fetch.prev_request_pc\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7888_ _3435_ _3628_ _3637_ _0384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8166__A1 _3462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7508__A4 core_0.ew_reg_ie\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9627_ _0637_ clknet_leaf_110_i_clk net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_119_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6839_ core_0.execute.alu_flag_reg.o_d\[1\] _2770_ _2771_ core_0.execute.pc_high_buff_out\[1\]
+ _2772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6716__A2 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4712__I _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9558_ _0568_ clknet_leaf_75_i_clk core_0.execute.sreg_irq_pc.o_d\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7228__C _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8509_ _1685_ core_0.execute.sreg_irq_pc.o_d\[7\] _4096_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9489_ _0499_ clknet_leaf_24_i_clk net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_122_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5455__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_70_i_clk clknet_4_12__leaf_i_clk clknet_leaf_70_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_232_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4663__B1 net321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8244__I2 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8803__B _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_85_i_clk clknet_4_15__leaf_i_clk clknet_leaf_85_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_233_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_1792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_13__f_i_clk_I clknet_3_6_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8157__A1 net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_218_3123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_218_3134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6707__A2 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7904__A1 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5915__B1 _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__A1 _0675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7933__I _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_23_i_clk clknet_4_9__leaf_i_clk clknet_leaf_23_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5143__A1 _1294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8880__A2 _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6891__A1 core_0.execute.pc_high_buff_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5170_ _1232_ _1241_ _1270_ _1319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_229_3263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_112_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8632__A2 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_i_clk clknet_4_8__leaf_i_clk clknet_leaf_38_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6643__A1 _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_147_2273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput4 i_core_int_sreg[12] net4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_223_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_56_Left_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_127_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8860_ net269 _4328_ _4327_ _4381_ _4382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7199__A2 _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6217__C _2205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7811_ core_0.execute.rf.reg_outputs\[9\]\[5\] _3591_ _3580_ _3593_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_204_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8791_ core_0.execute.irq_en net19 _4217_ core_0.execute.sreg_irq_flags.o_d\[4\]
+ _4321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_149_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8713__B _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6946__A2 _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7742_ core_0.execute.rf.reg_outputs\[11\]\[8\] _3548_ _3539_ _3553_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4954_ net66 core_0.fetch.out_buffer_data_instr\[7\] _0895_ _1134_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_143_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7673_ _3512_ _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_191_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4885_ _1051_ _1065_ _1066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9412_ _0422_ clknet_leaf_38_i_clk core_0.execute.rf.reg_outputs\[5\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_62_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8004__I _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6624_ _1328_ _2565_ _2566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_37_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Left_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5382__A1 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9343_ _0353_ clknet_leaf_31_i_clk core_0.execute.rf.reg_outputs\[9\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6555_ _2495_ _2496_ _2497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_6_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5506_ core_0.fetch.out_buffer_data_instr\[21\] net50 _1559_ _1580_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9274_ _0284_ clknet_leaf_155_i_clk core_0.execute.rf.reg_outputs\[13\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6486_ _1746_ _1839_ _2427_ _2428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_131_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6459__I _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8225_ _3846_ _3847_ _3848_ _3849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5437_ _1531_ _1532_ _1435_ _0037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8871__A2 _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5368_ _1464_ _1479_ _0021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8156_ _3446_ _3780_ _3791_ _0498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input44_I i_req_data[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7107_ _1768_ _2563_ _3033_ _3034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_227_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8087_ _3456_ _3738_ _3751_ _0469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5299_ _0995_ _1005_ _1399_ _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_0_214_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6634__A1 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7038_ _2672_ _2965_ _2966_ _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_74_Left_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4645__B1 net341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8989_ _0016_ clknet_leaf_141_i_clk core_0.dec_rf_ie\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6937__A2 net281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8623__B _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output200_I net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8139__A1 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_83_Left_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5373__B2 _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5474__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_213_3064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8311__A1 _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8862__A2 _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6873__A1 _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5676__A2 _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_2727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_2738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_168_Right_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_228_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8614__A2 _3256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5428__A2 _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6625__A1 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6318__B _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8378__A1 _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9330__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_200_2908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6928__A2 _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_196_2867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9480__CLK clknet_leaf_144_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5448__I _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4670_ core_0.execute.rf.reg_outputs\[6\]\[3\] _0670_ _0695_ core_0.execute.rf.reg_outputs\[10\]\[3\]
+ _0856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_113_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8550__A1 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5364__B2 _1476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6340_ _2153_ _2307_ _2309_ _2152_ _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__8302__A1 core_0.execute.alu_mul_div.mul_res\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6271_ core_0.execute.alu_mul_div.div_cur\[4\] _2256_ _2257_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5183__I _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5222_ _1356_ net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5667__A2 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8010_ _3453_ _3694_ _3707_ _0436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_149_2302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5153_ _1261_ _1246_ _1280_ _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__8605__A2 _4179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_135_Right_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5084_ core_0.decode.i_instr_l\[0\] _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_236_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4627__B1 net316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8912_ _2673_ _1251_ _4419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6092__A2 _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8843_ net252 _4328_ _4326_ _4366_ _4367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_84_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8774_ _4310_ _4295_ _4311_ _4307_ _0596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5986_ _1882_ _1973_ _1975_ _1897_ _1976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_47_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7725_ core_0.execute.rf.reg_outputs\[11\]\[0\] _3543_ _3539_ _3544_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4937_ _1111_ _1116_ _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ _3421_ _3497_ _3503_ _0286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4868_ _1017_ net54 _1048_ _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__6898__B _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7344__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8541__A1 _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5355__A1 core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6607_ _2547_ _2548_ _2549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_31_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7587_ _3387_ core_0.ew_data\[11\] _3449_ net23 _3459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_172_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4799_ _0942_ _0943_ _0980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
X_9326_ _0336_ clknet_leaf_40_i_clk core_0.execute.rf.reg_outputs\[10\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6538_ core_0.decode.oc_alu_mode\[4\] _2480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XTAP_TAPCELL_ROW_95_1655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9257_ _0267_ clknet_leaf_3_i_clk core_0.execute.rf.reg_outputs\[14\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__8844__A2 _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6469_ _2414_ _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_88_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6855__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8208_ _3828_ _1875_ _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_112_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput160 net160 o_req_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9188_ _0199_ clknet_leaf_44_i_clk core_0.ew_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xoutput171 net171 o_req_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput182 net182 sr_bus_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput193 net193 sr_bus_data_o[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8139_ net87 _3781_ _3771_ _3782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_102_Right_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_214_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__B1 net286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7280__A1 _2710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_214_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6853__S _2785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_214_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_180_2668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5830__A2 net322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_39_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7032__A1 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_214_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8780__A1 _0713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8532__A1 net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire210 net211 net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_25_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5346__A1 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_237_Right_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5897__A2 core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7099__A1 core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_238_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8835__A2 _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6846__A1 core_0.execute.sreg_irq_flags.o_d\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6846__B2 core_0.execute.trap_flag vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8528__B _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_226_3222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8599__A1 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclone100 _0702_ net347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_218_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A2 _1801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7271__B2 core_0.execute.sreg_scratch.o_d\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6990__C _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A2 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4791__B _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ _1518_ net180 _1830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_88_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7574__A2 core_0.ew_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8771__A1 _0765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_237_3351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5771_ _1749_ _1760_ _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_130_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_237_3362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7510_ _3389_ _3390_ _3391_ _3392_ _3393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
X_4722_ core_0.execute.pc_high_out\[2\] _0901_ _0904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_173_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8490_ _1738_ _4077_ _4078_ _4047_ _4079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7326__A2 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7441_ _3353_ _0221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5337__A1 _1239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ core_0.execute.rf.reg_outputs\[10\]\[4\] _0695_ _0700_ core_0.execute.rf.reg_outputs\[12\]\[4\]
+ _0840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5906__I _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_2372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_204_Right_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput40 i_req_data[11] net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput51 i_req_data[22] net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7372_ _2564_ _3288_ _3291_ _1768_ _3292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_114_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput62 i_req_data[3] net62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4584_ net88 _0666_ _0776_ _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_141_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9111_ _0001_ clknet_leaf_130_i_clk core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_114_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6323_ _2198_ _2301_ _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_0_i_clk_I i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6837__A1 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9042_ _0069_ clknet_leaf_90_i_clk core_0.fetch.out_buffer_data_instr\[30\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6254_ _2221_ _2240_ _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _1346_ _1347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6185_ core_0.execute.alu_mul_div.div_cur\[0\] _1883_ _2174_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_90_1596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5136_ core_0.execute.alu_mul_div.i_mul _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_35_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7262__A1 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6065__A2 _2054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5067_ _0902_ net110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7262__B2 core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer84_I _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_212_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7014__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8826_ _4349_ _4350_ _4351_ _4352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7565__A2 _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5576__A1 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8757_ core_0.execute.sreg_scratch.o_d\[5\] _4300_ _4302_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5969_ _1930_ _1958_ _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_43_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7708_ _3454_ _3520_ _3533_ _0308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_62_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8688_ _4203_ _4108_ _4251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7317__A2 _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5328__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7639_ core_0.execute.rf.reg_outputs\[14\]\[13\] _3482_ _3486_ _3493_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output198_I net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6421__B _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__A2 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_210_3034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9309_ _0319_ clknet_leaf_26_i_clk core_0.execute.rf.reg_outputs\[11\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4551__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output75_I net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5500__A1 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_2_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5803__A2 _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_3163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7005__A1 _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8753__A1 _0859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A1 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_193_2826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8505__A1 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7308__A2 _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_232_3292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8808__A2 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A2 net296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6819__A1 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6295__A2 _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__I _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8772__I net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7990_ _3401_ _3694_ _3696_ _0427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_135_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7795__A2 _3562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_68_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6941_ _2871_ _1314_ _2128_ _2872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_88_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6872_ _2010_ _2801_ _2803_ _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_44_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8611_ _3293_ _3330_ _4185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5558__A1 core_0.fetch.prev_request_pc\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5823_ _1772_ _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_157_2401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5558__B2 net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9591_ _0601_ clknet_leaf_41_i_clk core_0.execute.sreg_irq_flags.o_d\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_146_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8542_ net73 _4053_ _4125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5754_ _1518_ net188 _1744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4705_ core_0.execute.rf.reg_outputs\[6\]\[0\] _0670_ net318 core_0.execute.rf.reg_outputs\[4\]\[0\]
+ core_0.execute.rf.reg_outputs\[1\]\[0\] net302 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_8473_ net80 _4041_ _4064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4781__A2 _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5685_ net184 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_161_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7424_ _2703_ _3342_ _3343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4636_ net99 net324 _0824_ _0825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_79_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7355_ _2839_ _3274_ _3275_ _0213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5730__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4567_ core_0.execute.rf.reg_outputs\[14\]\[11\] _0685_ _0699_ core_0.execute.rf.reg_outputs\[12\]\[11\]
+ _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_92_1614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6306_ _2286_ _2279_ _2158_ _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7286_ _2480_ _3207_ _3208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_168_2530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4498_ core_0.execute.rf.reg_outputs\[1\]\[15\] _0693_ _0695_ core_0.execute.rf.reg_outputs\[10\]\[15\]
+ _0696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__8168__B _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6286__A2 _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9025_ _0052_ clknet_leaf_102_i_clk core_0.fetch.out_buffer_data_instr\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6237_ core_0.execute.alu_mul_div.div_cur\[0\] _2220_ _2225_ _2226_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_229_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_216_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_243_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6168_ core_0.execute.alu_mul_div.div_cur\[8\] net306 _2157_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7499__S _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7800__B _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6038__A2 net345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5119_ _1270_ _1273_ _1274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6099_ _2081_ _2082_ _2083_ _2088_ _2089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__8983__A1 _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7786__A2 _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5797__A1 _0960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8735__B2 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5549__A1 core_0.fetch.prev_request_pc\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8809_ core_0.execute.pc_high_buff_out\[1\] _4335_ _4337_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5549__B2 net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclone43 core_0.dec_r_reg_sel\[2\] net271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_62_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclone65 core_0.dec_r_reg_sel\[3\] net293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_85_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7710__A2 _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4524__A2 net318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5721__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5482__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__I _3562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8078__B _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_112_1861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5281__I _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6029__A2 _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_2202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7777__A2 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5788__A1 _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6326__B _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4835__I0 net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5252__A3 core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8726__A1 net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7529__A2 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6201__A2 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_234_3321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4763__A2 _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_2331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5470_ core_0.fetch.out_buffer_data_instr\[4\] net63 _1559_ _1560_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7162__B1 _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_2342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7701__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5712__A1 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4515__A2 _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7140_ _3065_ _2526_ _3066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7071_ core_0.execute.sreg_priv_control.o_d\[6\] _1692_ _2775_ core_0.execute.pc_high_out\[6\]
+ _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_74_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_245_3450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6022_ core_0.execute.rf.reg_outputs\[7\]\[4\] _1773_ _2012_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8716__B _1730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7217__A1 _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7620__B _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_2471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7973_ core_0.execute.rf.reg_outputs\[5\]\[10\] _3679_ _3677_ _3686_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6440__A2 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6924_ _2795_ _2848_ _2850_ _2480_ _2854_ _2855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_89_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8717__A1 _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5794__A4 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9643_ _0653_ clknet_leaf_129_i_clk core_0.dec_jump_cond_code\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6855_ _2711_ _2766_ _2787_ _2788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7846__I _3605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5806_ _0953_ _0955_ _0951_ _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_9574_ _0584_ clknet_leaf_19_i_clk core_0.execute.sreg_scratch.o_d\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6786_ _1896_ _2715_ _2718_ _2719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_119_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7940__A2 _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_107_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6743__A3 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8525_ _4041_ _4108_ _4109_ _4110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5951__A1 net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5737_ net198 _1729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8456_ net215 _4048_ _2766_ _2133_ _2784_ _4049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_33_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5668_ _1540_ _1674_ _1675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_33_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7407_ _2587_ _3179_ _3323_ _3325_ _3326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_60_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4619_ core_0.execute.rf.reg_outputs\[14\]\[7\] net310 net308 core_0.execute.rf.reg_outputs\[1\]\[7\]
+ _0809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4506__A2 _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5703__A1 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8387_ core_0.execute.alu_mul_div.mul_res\[14\] _3998_ _3863_ _3999_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5599_ core_0.decode.i_instr_l\[12\] _1616_ _1632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7338_ core_0.execute.alu_mul_div.div_res\[13\] _1742_ _3258_ _3259_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_40_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7269_ core_0.execute.alu_mul_div.div_cur\[11\] _1317_ _3191_ _3192_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_229_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9008_ _0035_ clknet_leaf_131_i_clk core_0.dec_alu_flags_ie vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7759__A2 _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4690__B2 core_0.execute.rf.reg_outputs\[12\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8420__A3 _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6431__A2 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8708__A1 _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8184__A2 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7931__A2 _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__A2 _2439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8587__I _4159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7705__B _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_2769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7998__A2 _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6670__A2 _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4681__A1 core_0.execute.rf.reg_outputs\[9\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6958__B1 _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8411__A3 _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_240_3391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6422__A2 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4970_ core_0.fetch.prev_request_pc\[7\] core_0.fetch.prev_request_pc\[6\] _1149_
+ _1150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_230_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_103_Left_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_199_2898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6640_ _1929_ _2569_ _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_156_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5233__I0 core_0.ew_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4736__A2 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6571_ _2497_ _2512_ _2513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8310_ _3919_ _3921_ _3926_ _3927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5522_ net58 _1556_ _1588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9290_ _0300_ clknet_leaf_155_i_clk core_0.execute.rf.reg_outputs\[12\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8241_ _3829_ _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_42_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7615__B _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6489__A2 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5453_ _1001_ _1547_ _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_152_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8172_ net93 _3779_ _3797_ _3800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5161__A2 _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5384_ _1241_ _1490_ _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7123_ _3004_ _3049_ _3050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7438__A1 net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7989__A2 _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7054_ net260 net214 _2982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6110__A1 core_0.execute.rf.reg_outputs\[7\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6110__B2 core_0.execute.rf.reg_outputs\[5\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6005_ core_0.execute.rf.reg_outputs\[2\]\[12\] _1797_ _1781_ core_0.execute.rf.reg_outputs\[10\]\[12\]
+ _1995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_157_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_214_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_33_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8938__A1 core_0.decode.i_imm_pass\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__A2 _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7956_ _3414_ _3672_ _3676_ _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_179_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6907_ _2838_ _0202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7887_ core_0.execute.rf.reg_outputs\[7\]\[5\] _3634_ _3636_ _3637_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7576__I _3450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8166__A2 _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6480__I _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9626_ _0636_ clknet_leaf_132_i_clk net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6838_ _1405_ _1691_ _2692_ _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_175_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__C _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4727__A2 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9557_ _0567_ clknet_leaf_74_i_clk core_0.execute.sreg_irq_pc.o_d\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_190_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5924__A1 core_0.execute.rf.reg_outputs\[13\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _2699_ _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_18_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8508_ _4039_ _4094_ _4095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9488_ _0498_ clknet_leaf_24_i_clk net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_162_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output180_I net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7677__A1 _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_149_Right_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_8439_ _2230_ _4035_ _0537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_98_1686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_4_i_clk clknet_4_2__leaf_i_clk clknet_leaf_4_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5152__A2 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6101__A1 _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7260__B core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4663__A1 core_0.execute.rf.reg_outputs\[3\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4663__B2 core_0.execute.rf.reg_outputs\[12\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8244__I3 _2115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__A2 _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_212_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_218_3124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8157__A2 _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__I _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7904__A2 _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_116_Right_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8110__I _3758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6891__A2 _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_229_3264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8093__A1 _3465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_242_3420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_147_2274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 i_core_int_sreg[13] net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_189_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_189_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_160_2430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7810_ _3428_ _3585_ _3592_ _0351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_188_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8790_ _4249_ _4320_ _1435_ _0603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_231_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7741_ _3447_ _3542_ _3552_ _0322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4953_ _1128_ _1132_ _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7329__C _3073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7672_ _0891_ _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4884_ _1011_ _1014_ _1064_ _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_157_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9411_ _0421_ clknet_leaf_38_i_clk core_0.execute.rf.reg_outputs\[5\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_46_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_82_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6623_ _1929_ _1874_ _2565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_7_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9342_ _0352_ clknet_leaf_28_i_clk core_0.execute.rf.reg_outputs\[9\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6554_ _2074_ _2349_ _2496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5505_ _1579_ _0059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7659__A1 _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_171_2570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9273_ _0283_ clknet_leaf_4_i_clk core_0.execute.rf.reg_outputs\[13\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6485_ net314 net206 _2427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8224_ _1537_ _1540_ _2344_ _3848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5436_ core_0.dec_pc_inc _1438_ _1532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8155_ net100 _3787_ _3785_ _3791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_227_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5367_ core_0.dec_rf_ie\[11\] _1438_ _1472_ _1478_ _1479_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4893__A1 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7106_ _2586_ _3031_ _3032_ _3033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__8084__A1 core_0.execute.rf.reg_outputs\[2\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8086_ core_0.execute.rf.reg_outputs\[2\]\[10\] _3743_ _3745_ _3751_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8176__B _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5298_ core_0.dec_sreg_store _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_input37_I i_mem_exception vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ core_0.dec_mem_access net204 _2966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7831__A1 _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4645__B2 core_0.execute.rf.reg_outputs\[3\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6398__A1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8988_ _0015_ clknet_leaf_138_i_clk core_0.dec_rf_ie\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_218_Right_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_194_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7939_ _3460_ _3652_ _3666_ _0406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6424__B _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8139__A2 _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9609_ _0619_ clknet_leaf_60_i_clk core_0.execute.pc_high_buff_out\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7898__A1 _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5373__A2 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_208_Left_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_213_3065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8311__A2 _2521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_152_i_clk clknet_4_0__leaf_i_clk clknet_leaf_152_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_104_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8865__I _4385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6873__A2 _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_2728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4884__A1 _1011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8086__B _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5428__A3 _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4636__A1 net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_217_Left_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5833__B1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_109_1822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8378__A2 _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6389__A1 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_200_2909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8533__C _4046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9625__CLK clknet_leaf_133_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_196_2868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7889__A1 core_0.execute.rf.reg_outputs\[7\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_226_Left_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8550__A2 _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5364__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7165__B _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5464__I _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6270_ core_0.execute.alu_mul_div.comp _0998_ _2255_ _2256_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__5116__A2 _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5221_ core_0.ew_data\[6\] net156 _1356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_149_2303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4875__A1 _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8708__C _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5152_ _1260_ _1247_ _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_209_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_235_Left_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7813__A1 core_0.execute.rf.reg_outputs\[9\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5083_ _1239_ _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_223_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5824__B1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__B2 core_0.execute.rf.reg_outputs\[8\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8911_ _1231_ _1529_ _4418_ _0626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8724__B _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8842_ _4324_ _4365_ _4366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_195_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8773_ core_0.execute.sreg_scratch.o_d\[12\] _4300_ _4311_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5985_ _1882_ _1974_ _1975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5052__A1 core_0.fetch.prev_request_pc\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7724_ _3541_ _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4936_ _1112_ _1113_ _1114_ _1115_ _1116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_93_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_244_Left_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_10 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7655_ core_0.execute.rf.reg_outputs\[13\]\[3\] _3498_ _3500_ _3503_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4867_ _0892_ _1047_ _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6606_ _2546_ _1999_ _2469_ _2548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_34_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5355__A2 core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6552__A1 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7586_ _3403_ _3457_ _3458_ _0261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_132_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4798_ core_0.ew_reg_ie\[14\] _0959_ _0960_ core_0.ew_reg_ie\[15\] _0979_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_6_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9325_ _0335_ clknet_leaf_32_i_clk core_0.execute.rf.reg_outputs\[10\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6537_ net212 _1974_ _2478_ _2479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4563__B1 _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9256_ _0266_ clknet_leaf_150_i_clk core_0.execute.rf.reg_outputs\[15\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_95_1656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6304__A1 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ net70 _1371_ _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5307__C _0922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8207_ _3830_ _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6855__A2 _2766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5419_ _1516_ _0035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput150 net150 o_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_84_i_clk clknet_4_14__leaf_i_clk clknet_leaf_84_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_9187_ _0198_ clknet_leaf_47_i_clk net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput161 net161 o_req_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6399_ _1674_ _2370_ _2371_ _2372_ _1539_ _2373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xoutput172 net172 o_req_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput183 net183 sr_bus_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8138_ _3779_ _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput194 net194 sr_bus_data_o[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6068__B1 net331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_215_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7804__A1 core_0.execute.rf.reg_outputs\[9\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8069_ _3414_ _3737_ _3741_ _0461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_242_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__B2 core_0.execute.rf.reg_outputs\[13\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_99_i_clk clknet_4_13__leaf_i_clk clknet_leaf_99_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_3_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_2669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5291__A1 core_0.dec_sreg_store vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_22_i_clk clknet_4_3__leaf_i_clk clknet_leaf_22_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_194_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8780__A2 _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6791__A1 _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_2_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8532__A2 _2134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire211 _2606_ net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_81_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_37_i_clk clknet_4_10__leaf_i_clk clknet_leaf_37_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_155_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6543__A1 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4554__B1 _0693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5897__A3 core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8296__A1 _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7099__A2 _2439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6846__A2 _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7713__B _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8048__A1 core_0.execute.rf.reg_outputs\[3\]\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_226_3223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_245_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7271__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8220__A1 core_0.execute.alu_mul_div.mul_res\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7023__A2 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5034__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8771__A2 _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5770_ _1751_ _1753_ _1757_ _1759_ _1760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__6782__A1 _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_237_3352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4721_ core_0.execute.prev_pc_high\[3\] _0902_ _0903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5990__C1 _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8523__A2 _4107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7440_ net125 _2954_ _2415_ _3353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6534__A1 _2468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4652_ core_0.execute.rf.reg_outputs\[4\]\[4\] _0720_ _0708_ core_0.execute.rf.reg_outputs\[13\]\[4\]
+ _0839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_2373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput30 i_mem_data[3] net30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput41 i_req_data[12] net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7371_ _2568_ _3289_ _3290_ _2564_ _3291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xinput52 i_req_data[23] net52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5194__I _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4583_ _0770_ _0775_ _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_142_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput63 i_req_data[4] net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9110_ _0000_ clknet_leaf_113_i_clk core_0.execute.alu_mul_div.i_mod vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6322_ _2300_ _2293_ _2301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8719__B _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9041_ _0068_ clknet_leaf_90_i_clk core_0.fetch.out_buffer_data_instr\[29\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6253_ _2210_ _2239_ _2240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6837__A2 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4848__A1 _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8039__A1 _3434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5204_ core_0.ew_addr\[0\] core_0.ew_mem_width _1346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6184_ core_0.execute.alu_mul_div.div_cur\[1\] _2076_ _2172_ _2173_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_237_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5135_ _1261_ _1288_ _1289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_90_1597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _0904_ net109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_rebuffer77_I net304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8211__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8825_ core_0.execute.pc_high_buff_out\[3\] _4335_ _4351_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5025__A1 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8762__A2 _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6773__A1 core_0.ew_data\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5576__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5968_ _1897_ _1943_ _1957_ _1958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8756_ net243 _4294_ _4301_ _4287_ _0588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_149_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ core_0.fetch.prev_request_pc\[12\] _1020_ _1026_ core_0.fetch.prev_request_pc\[13\]
+ _1099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_192_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7707_ core_0.execute.rf.reg_outputs\[12\]\[9\] _3526_ _3528_ _3533_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8687_ net86 _1740_ _1719_ _4250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5899_ core_0.decode.oc_alu_mode\[3\] _1888_ _1889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7584__I _3456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6525__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7638_ _3463_ _3477_ _3492_ _0279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5328__A2 _1313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4536__B1 _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7569_ _3381_ _3443_ _3444_ _3445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_160_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_210_3035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8278__A1 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9308_ _0318_ clknet_leaf_9_i_clk core_0.execute.rf.reg_outputs\[11\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9239_ _0013_ clknet_leaf_106_i_clk core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__4839__A1 _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5500__A2 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6149__B _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8450__A1 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_6_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_81_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5803__A3 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_221_3164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5016__A1 _1185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8753__A2 _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A2 _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_193_2827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4527__B1 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_3293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8441__A1 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6940_ core_0.execute.alu_mul_div.div_res\[3\] _2871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_89_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6871_ _2010_ _2802_ _2803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_240_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5007__A1 _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5822_ _1811_ _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
X_8610_ _4184_ _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_159_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9590_ _0600_ clknet_leaf_41_i_clk core_0.execute.sreg_irq_flags.o_d\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_33_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5558__A2 _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6755__A1 _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_2402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8721__C _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8541_ _1736_ _4120_ _4123_ _4124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5753_ core_0.execute.alu_mul_div.i_mul _1743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_8_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9536__D _0546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4704_ core_0.execute.rf.reg_outputs\[2\]\[0\] net250 _0695_ core_0.execute.rf.reg_outputs\[10\]\[0\]
+ _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7337__C _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8472_ net80 _4058_ _4063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5684_ _1687_ _1688_ _1423_ _1424_ _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_32_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7423_ _3304_ _3341_ _3342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_154_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4635_ _0818_ _0823_ _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_71_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7354_ core_0.ew_data\[13\] _3168_ _3275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4566_ core_0.execute.rf.reg_outputs\[6\]\[11\] _0669_ _0692_ core_0.execute.rf.reg_outputs\[1\]\[11\]
+ _0760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_130_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6305_ _2157_ _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_130_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7285_ _2468_ _2472_ _3207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5652__I _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4497_ net221 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_228_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_168_2531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9024_ _0051_ clknet_leaf_102_i_clk core_0.fetch.out_buffer_data_instr\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6236_ _2221_ _2222_ _2223_ _2224_ _2225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8680__A1 _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5494__A1 net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6167_ core_0.execute.alu_mul_div.div_cur\[10\] _2155_ _2156_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_176_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_103_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5118_ core_0.decode.i_instr_l\[1\] core_0.decode.i_instr_l\[0\] _1273_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6098_ _2084_ _2085_ _2086_ _2087_ _2088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_240_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__B _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5049_ net80 _1085_ _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_224_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6994__A1 _2710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5797__A2 _0951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8735__A2 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8808_ core_0.execute.pc_high_out\[1\] core_0.execute.pc_high_out\[0\] _4336_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5549__A2 _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_2660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6746__A1 net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7528__B _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8739_ _4289_ _4290_ _1435_ _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6432__B _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4731__I _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8499__A1 _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclone22 _0672_ net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_164_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_28_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7171__A1 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8671__A1 net279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5485__A1 net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_158_Left_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_216_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_128_2047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8423__A1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8094__B _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8974__A2 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4906__I _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_215_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_19_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6985__A1 _1254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5788__A2 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6985__B2 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_205_2970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8726__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6737__A1 _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_167_Left_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_1991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_234_3322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5737__I net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7157__C core_0.execute.alu_mul_div.i_mod vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5960__A2 _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4763__A3 core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_152_2332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7162__B2 core_0.execute.sreg_scratch.o_d\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7070_ core_0.execute.pc_high_buff_out\[6\] _2771_ _2774_ core_0.execute.sreg_irq_pc.o_d\[6\]
+ _2998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_176_Left_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8662__A1 _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_226_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_245_3451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6021_ _2010_ _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_238_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8783__I _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7901__B _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8716__C _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8414__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_234_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4816__I core_0.execute.alu_mul_div.i_mod vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_2472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7972_ _3453_ _3672_ _3685_ _0420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6236__C _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6923_ _1880_ _2510_ _2853_ _2854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8732__B _4283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_185_Left_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_9642_ _0652_ clknet_leaf_129_i_clk core_0.dec_jump_cond_code\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__6728__A1 net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6854_ core_0.dec_mem_access _2786_ _2787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4739__B1 _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5805_ core_0.execute.rf.reg_outputs\[13\]\[0\] _1792_ _1794_ core_0.execute.rf.reg_outputs\[8\]\[0\]
+ _1795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_9573_ _0583_ clknet_leaf_63_i_clk net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6785_ _2716_ _2717_ _2718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8524_ _2403_ _4041_ _1735_ _1433_ _4109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_134_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ _1714_ _1728_ _0141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5951__A2 _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8455_ _1419_ _1403_ _4048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_33_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5667_ _1542_ _1544_ _1674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4618_ core_0.execute.rf.reg_outputs\[12\]\[7\] _0699_ net286 core_0.execute.rf.reg_outputs\[13\]\[7\]
+ _0808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7406_ _2588_ _3324_ _2587_ _3325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8386_ _2370_ _3827_ _3996_ _3997_ _3998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_170_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4506__A3 core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5598_ _1629_ _1631_ _0100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input67_I i_req_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4911__B1 _1057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7337_ _1743_ _3256_ _3257_ _0996_ _3258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XPHY_EDGE_ROW_194_Left_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4549_ core_0.execute.rf.reg_outputs\[3\]\[12\] _0698_ _0708_ core_0.execute.rf.reg_outputs\[13\]\[12\]
+ _0744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_102_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7268_ _3170_ _1314_ _3189_ _3190_ core_0.execute.alu_mul_div.i_mod _3191_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_96_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9007_ _0034_ clknet_leaf_131_i_clk core_0.dec_alu_carry_en vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6219_ _2180_ _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7811__B _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7199_ net86 _2995_ _3123_ _2893_ _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_244_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8405__A1 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6427__B _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__A2 net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5050__C _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8642__B _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6719__A1 _2654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5927__C1 net336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5557__I _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5942__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__A1 net306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5155__B1 _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8644__A1 _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8536__C _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4681__A2 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8947__A2 _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6958__A1 core_0.execute.sreg_irq_flags.o_d\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_3392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A1 core_0.decode.i_imm_pass\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_2899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7383__A1 _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5233__I1 core_0.ew_data\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6570_ _2495_ _2496_ _2512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5394__B1 _1494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5521_ _1018_ _1552_ _1587_ _0067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8240_ core_0.execute.alu_mul_div.mul_res\[4\] _3862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_124_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ _1546_ _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__8883__A1 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5697__A1 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6894__B1 _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8171_ _3469_ _3781_ _3799_ _0505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5383_ _1236_ _1316_ _1490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7122_ _1683_ core_0.execute.sreg_irq_pc.o_d\[7\] _3048_ _3049_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_239_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7438__A2 _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8635__A1 _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ _1337_ _2487_ _1285_ _2981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7631__B _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6110__A2 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6004_ core_0.execute.rf.reg_outputs\[5\]\[12\] _1785_ _1802_ core_0.execute.rf.reg_outputs\[14\]\[12\]
+ _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__9531__CLK clknet_leaf_74_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8938__A2 _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4546__I _0741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6949__A1 _2694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7071__B1 _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4990__B _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7955_ core_0.execute.rf.reg_outputs\[5\]\[2\] _3673_ _3663_ _3676_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5621__A1 _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5472__I1 net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6906_ core_0.ew_data\[2\] _2837_ _0199_ _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8181__C _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7886_ _3512_ _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_77_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_2630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9625_ _0635_ clknet_leaf_133_i_clk net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_108_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _1686_ net227 _1410_ _2770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
Xclkbuf_4_4__f_i_clk clknet_3_2_0_i_clk clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7374__A1 _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9556_ _0566_ clknet_leaf_69_i_clk core_0.execute.sreg_irq_pc.o_d\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6768_ _2673_ _2698_ _2701_ _2702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5924__A2 _1791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8507_ _4041_ _4092_ _4093_ _4094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7806__B _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7126__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5719_ _0801_ _1704_ _1717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6699_ core_0.execute.rf.reg_outputs\[1\]\[3\] _2608_ _2609_ core_0.execute.rf.reg_outputs\[3\]\[3\]
+ _2638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7592__I _3462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9487_ _0497_ clknet_leaf_62_i_clk net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__8874__A1 _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7677__A2 _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8438_ _4022_ _4031_ core_0.execute.alu_mul_div.div_res\[12\] _4035_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_98_1687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output173_I net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5326__B _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8369_ _3981_ _3982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8626__A1 _1696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6101__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8356__C _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__A2 _0698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_202_2940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5612__A1 _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_218_3125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7365__A1 _2370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6168__A2 net306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7365__B2 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5915__A2 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__B _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7668__A2 _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9554__CLK clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_229_3265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8093__A2 _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5750__I _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_242_3421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_223_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7840__A2 _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_2275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5851__A1 net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput6 i_core_int_sreg[14] net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_160_2431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5603__A1 core_0.decode.i_instr_l\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4952_ _1115_ _1127_ _1129_ _1131_ _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
X_7740_ core_0.execute.rf.reg_outputs\[11\]\[7\] _3548_ _3539_ _3552_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4883_ _1054_ _1057_ _1060_ _1063_ _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_7671_ _3457_ _3498_ _3511_ _0293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6159__A2 _1837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9410_ _0420_ clknet_leaf_37_i_clk core_0.execute.rf.reg_outputs\[5\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_117_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5367__B1 _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6622_ _2563_ _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_6_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6553_ _1748_ _2492_ _2495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_9341_ _0351_ clknet_leaf_28_i_clk core_0.execute.rf.reg_outputs\[9\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5504_ core_0.fetch.out_buffer_data_instr\[20\] net49 _1559_ _1579_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_171_2560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7345__C _2689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6484_ net248 _1942_ _2425_ _2426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9272_ _0282_ clknet_leaf_149_i_clk core_0.execute.rf.reg_outputs\[14\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7659__A2 _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8223_ _3834_ _3840_ _3838_ _3847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5435_ _1528_ _1529_ _1530_ _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5861__S _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8608__A1 core_0.execute.alu_flag_reg.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ core_0.decode.i_instr_l\[9\] _1465_ _1440_ _1478_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8154_ _3440_ _3780_ _3790_ _0497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4893__A2 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7361__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7105_ _2586_ _2843_ _3032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8084__A2 _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8085_ _3453_ _3737_ _3750_ _0468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_226_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5297_ _1417_ _1415_ _1418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__5660__I core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7036_ _2703_ _2954_ _2962_ _2964_ _2965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7831__A2 _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4645__A2 net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__A1 _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8987_ _1497_ _4461_ _0659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6398__A2 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7595__B2 net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_182_Right_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7938_ core_0.execute.rf.reg_outputs\[6\]\[11\] _3657_ _3663_ _3666_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4802__C1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7869_ _3470_ _3607_ _3625_ _0377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_46_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9427__CLK clknet_leaf_16_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9608_ _0618_ clknet_leaf_60_i_clk core_0.execute.pc_high_buff_out\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5358__B1 _1470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7898__A2 _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__I0 net39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_122_Left_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_9539_ _0549_ clknet_leaf_77_i_clk net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_46_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6440__B _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_213_3066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output98_I net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_2729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Right_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5570__I _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_131_Left_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7822__A2 _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_151_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4636__A2 net324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5833__B2 core_0.execute.rf.reg_outputs\[14\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_224_3195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6615__B _2556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7586__A1 _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Right_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_196_2869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4850__S _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8322__S _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Left_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7889__A2 _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6010__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8121__I _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8838__A1 core_0.execute.pc_high_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_76_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7960__I _3671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _1355_ net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Right_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_2304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5151_ _1301_ _1303_ _1304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8066__A2 _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5413__C _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5082_ core_0.decode.i_instr_l\[6\] _1238_ core_0.decode.i_instr_l\[5\] _1239_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__7813__A2 _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5824__A1 core_0.execute.rf.reg_outputs\[8\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__A2 _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5824__B2 core_0.execute.rf.reg_outputs\[4\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8910_ _1685_ _1286_ _4418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7026__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8841_ _4335_ _4363_ _4364_ _4365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_189_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9539__D _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_50_Right_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_3_i_clk clknet_4_2__leaf_i_clk clknet_leaf_3_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8772_ net196 _4310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_177_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5984_ _1828_ _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7723_ _3541_ _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4935_ core_0.fetch.prev_request_pc\[0\] _1054_ _1043_ core_0.fetch.prev_request_pc\[1\]
+ core_0.fetch.prev_request_pc\[2\] _1063_ _1115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_176_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7329__A1 _2371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__B1 _3120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7329__B2 net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4760__S net293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_11 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7654_ _3415_ _3497_ _3502_ _0285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4866_ core_0.fetch.out_buffer_data_instr\[25\] _1047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6605_ _2546_ _1999_ _2469_ _2547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7356__B _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5355__A3 core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4797_ core_0.ew_reg_ie\[12\] _0950_ _0956_ core_0.ew_reg_ie\[13\] _0978_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7585_ core_0.execute.rf.reg_outputs\[15\]\[10\] _3429_ _3422_ _3458_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_31_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8829__A1 core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9324_ _0334_ clknet_leaf_8_i_clk core_0.execute.rf.reg_outputs\[10\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6536_ _2423_ _2476_ _2477_ _2478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4563__B2 core_0.execute.rf.reg_outputs\[3\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer22_I _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9255_ _0265_ clknet_leaf_150_i_clk core_0.execute.rf.reg_outputs\[15\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7501__A1 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6467_ _2413_ _0911_ _0187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8206_ _3822_ _3826_ _3827_ _1812_ _3831_ _0508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xoutput140 net140 o_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5418_ core_0.dec_alu_flags_ie _1251_ _1293_ _1506_ _1516_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_101_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput151 net151 o_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9186_ _0197_ clknet_leaf_46_i_clk net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6398_ _2354_ _1544_ _2372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_140_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput162 net162 o_req_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput173 net173 o_req_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput184 net184 sr_bus_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5349_ _1439_ _1465_ core_0.decode.i_instr_l\[7\] _1466_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__8057__A2 _3714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8137_ _3779_ _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput195 net304 sr_bus_data_o[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5390__I _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6068__A1 core_0.execute.rf.reg_outputs\[13\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7804__A2 _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8068_ core_0.execute.rf.reg_outputs\[2\]\[2\] _3738_ _3730_ _3741_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4618__A2 _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output136_I net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7019_ _2501_ _2946_ _2947_ _2948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_3_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8634__C _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5291__A2 _1411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6791__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_191_2799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4554__B2 core_0.execute.rf.reg_outputs\[1\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5897__A4 core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8296__A2 _1680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8097__B _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6396__I _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8048__A2 _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_226_3224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_2245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7559__A1 _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6345__B _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8220__A2 _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5034__A2 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_237_3353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6782__A2 _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4720_ core_0.execute.pc_high_out\[3\] _0901_ _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__4793__A1 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5990__B1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5990__C2 core_0.execute.rf.reg_outputs\[3\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7176__B _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4651_ core_0.execute.rf.reg_outputs\[6\]\[4\] _0670_ _0683_ core_0.execute.rf.reg_outputs\[7\]\[4\]
+ _0838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7731__A1 core_0.execute.rf.reg_outputs\[11\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput20 i_mem_ack net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_2374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput31 i_mem_data[4] net31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4545__A1 _0730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7370_ _2568_ _3139_ _3290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4582_ _0771_ _0772_ _0773_ _0774_ _0775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_126_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput42 i_req_data[13] net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput53 i_req_data[24] net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput64 i_req_data[5] net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6321_ _2156_ _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__8287__A2 _3854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9040_ _0067_ clknet_leaf_88_i_clk core_0.fetch.out_buffer_data_instr\[28\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6252_ _2176_ _2232_ _2238_ _2239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__9122__CLK clknet_leaf_108_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6837__A3 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5203_ _1345_ core_0.fetch.current_req_branch_pred vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8039__A2 _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6183_ _2170_ _2171_ _2172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5134_ _1242_ _1235_ _1288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_90_1587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _0905_ net108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8824_ core_0.execute.pc_high_out\[3\] _4342_ _4329_ _4350_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_151_i_clk clknet_4_0__leaf_i_clk clknet_leaf_151_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8211__A2 _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clone42_I _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8755_ core_0.execute.sreg_scratch.o_d\[4\] _4300_ _4301_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_181_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _1882_ _1956_ _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6773__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7970__A1 _3450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7706_ _3451_ _3520_ _3532_ _0307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4918_ _1094_ _1097_ _1098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8686_ _1661_ _4249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_35_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5981__B1 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4784__B2 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5898_ _1766_ _1886_ _1887_ _1888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_192_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7637_ core_0.execute.rf.reg_outputs\[14\]\[12\] _3482_ _3486_ _3492_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4849_ _1020_ _1023_ _1026_ _1029_ _1030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7722__A1 core_0.ew_reg_ie\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4536__A1 core_0.execute.rf.reg_outputs\[3\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5584__I0 _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7568_ net34 _1348_ _3444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9307_ _0317_ clknet_leaf_4_i_clk core_0.execute.rf.reg_outputs\[11\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_210_3036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8278__A2 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6519_ net319 _1925_ _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_120_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7499_ core_0.dec_mem_width core_0.ew_mem_width _2421_ _3384_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6289__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9238_ _0249_ clknet_leaf_133_i_clk core_0.ew_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_113_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9169_ _0180_ clknet_leaf_43_i_clk core_0.execute.prev_pc_high\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_104_i_clk clknet_4_12__leaf_i_clk clknet_leaf_104_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_227_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_227_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7789__A1 _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8645__B _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8986__B1 _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8450__A2 _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_24_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__A1 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_3165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_119_i_clk clknet_4_5__leaf_i_clk clknet_leaf_119_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5016__A2 _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_183_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7961__A1 core_0.execute.rf.reg_outputs\[5\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_193_2828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4775__A1 _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7713__A1 core_0.execute.rf.reg_outputs\[12\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4527__A1 core_0.execute.rf.reg_outputs\[1\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__B2 core_0.execute.rf.reg_outputs\[10\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_232_3294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_234_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _2001_ _1958_ _1930_ _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6204__A1 _2165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ net87 _1772_ _1783_ _1810_ _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_201_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_233_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7952__A1 _3401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7685__I _3519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6755__A2 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_83_i_clk clknet_4_14__leaf_i_clk clknet_leaf_83_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_159_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8540_ _4039_ _4122_ _4123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5963__B1 _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ _0996_ _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_174_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4703_ core_0.execute.rf.reg_outputs\[11\]\[0\] net303 net341 core_0.execute.rf.reg_outputs\[3\]\[0\]
+ _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_8471_ _1702_ _4054_ _4062_ _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_173_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5683_ net191 _1688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_151_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7704__A1 _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7422_ _1685_ _3339_ _3340_ _3341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_4_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4634_ _0819_ _0820_ _0821_ _0822_ _0823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_32_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_98_i_clk clknet_4_13__leaf_i_clk clknet_leaf_98_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7353_ _2672_ net295 _3273_ _3274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4565_ core_0.execute.rf.reg_outputs\[2\]\[11\] _0672_ _0707_ core_0.execute.rf.reg_outputs\[13\]\[11\]
+ _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5191__A1 core_0.decode.oc_alu_mode\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6304_ _2219_ _2284_ _2285_ _0152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7284_ _3206_ _0211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4496_ _0661_ _0662_ _0668_ _0664_ _0694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_228_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_i_clk clknet_4_9__leaf_i_clk clknet_leaf_21_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_9023_ _0050_ clknet_leaf_80_i_clk core_0.fetch.out_buffer_data_instr\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_168_2532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Right_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6235_ _2215_ _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_228_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5494__A2 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6166_ _1833_ _2155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_243_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_225_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5117_ _1271_ _1272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__8432__A2 _4031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6097_ core_0.execute.rf.reg_outputs\[3\]\[3\] _0948_ _0962_ _2087_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_36_i_clk clknet_4_8__leaf_i_clk clknet_leaf_36_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8184__C _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5048_ _1215_ _1060_ _1145_ _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_197_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input12_I i_core_int_sreg[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6994__A2 _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_212_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8196__A1 _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8807_ _4334_ _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_67_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7809__B _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_2661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6999_ _2839_ _2927_ _2928_ _0204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7943__A1 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__A2 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4757__A1 core_0.ew_reg_ie\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8738_ core_0.execute.sreg_jtr_buff.o_d\[1\] _4217_ _1415_ _4290_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_192_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8669_ _1658_ _4232_ _4235_ _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_35_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclone34 _0685_ net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_145_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4509__A1 core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone56 _0707_ net284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_145_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclone78 net313 net207 _1847_ net306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_106_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5182__A1 _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output80_I net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8120__A1 _3450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8671__A2 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_1852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5485__A2 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4693__B1 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6674__I _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8423__A2 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_141_2204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A3 _0951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_205_2971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4996__A1 _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8187__A1 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4748__A1 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_123_1992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5945__B1 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_234_3323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4763__A4 core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7162__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_2333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__I core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8111__A1 core_0.execute.rf.reg_outputs\[1\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__B1 _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6673__A1 _2607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6020_ _2009_ _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_245_3452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I i_core_int_sreg[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_207_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8414__A2 _1670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7971_ core_0.execute.rf.reg_outputs\[5\]\[9\] _3679_ _3677_ _3685_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_163_2473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6922_ _2075_ _2851_ _2852_ _2853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8178__A1 _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9310__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9641_ _0651_ clknet_leaf_139_i_clk core_0.dec_jump_cond_code\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7629__B _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ _2700_ _2701_ _2785_ _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6189__B1 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6728__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7925__A1 core_0.execute.rf.reg_outputs\[6\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5804_ _1793_ _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_186_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9572_ _0582_ clknet_4_9__leaf_i_clk core_0.execute.trap_flag vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6784_ _1930_ _1882_ _2717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_29_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5400__A2 _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8523_ _2403_ _4107_ _4108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5735_ core_0.execute.sreg_priv_control.o_d\[13\] _1700_ _1727_ _1697_ _1728_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_174_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8454_ _4046_ _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_161_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5666_ _1671_ _1672_ _1673_ _0126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8350__A1 core_0.execute.alu_mul_div.mul_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7153__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7364__B _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7405_ net270 _3243_ _3324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5164__A1 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4617_ core_0.execute.rf.reg_outputs\[6\]\[7\] net223 net312 core_0.execute.rf.reg_outputs\[2\]\[7\]
+ _0807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8385_ _3993_ _3995_ _3828_ _3997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6900__A2 _2785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4506__A4 _0675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5597_ _1591_ net40 _1369_ _1630_ _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_142_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4911__A1 core_0.fetch.prev_request_pc\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7336_ core_0.execute.alu_mul_div.i_mul core_0.execute.alu_mul_div.mul_res\[13\]
+ _3257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4911__B2 core_0.fetch.prev_request_pc\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4548_ core_0.execute.rf.reg_outputs\[10\]\[12\] _0695_ _0705_ core_0.execute.rf.reg_outputs\[9\]\[12\]
+ _0743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8102__A1 core_0.execute.rf.reg_outputs\[1\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8653__A2 _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7267_ _2124_ core_0.execute.alu_mul_div.mul_res\[11\] core_0.execute.alu_mul_div.i_div
+ _3190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4479_ net222 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
X_9006_ _0033_ clknet_leaf_135_i_clk core_0.dec_l_reg_sel\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6664__B2 _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6218_ core_0.execute.alu_mul_div.div_cur\[3\] _2075_ _2207_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7198_ _3121_ _3122_ _3123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4675__B1 net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ _1741_ _2138_ _1435_ _0144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5219__A2 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7464__I0 core_0.dec_rf_ie\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6967__A2 _2881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8169__A1 _3465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8964__I0 net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7258__C _2563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5927__B1 net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7392__A2 _2556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8341__A1 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7144__A2 _1925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_88_Right_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__A1 _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__B2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8892__A2 _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4902__A1 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6104__B1 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8644__A2 _4042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6655__A1 _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_196_Right_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_73_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4666__B1 net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Right_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9333__CLK clknet_leaf_155_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6958__A2 _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7080__A1 _2708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_240_3393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5091__B1 _1244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7207__I0 core_0.ew_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5630__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5918__B1 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8580__A1 _2918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Left_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5394__A1 core_0.decode.i_imm_pass\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5394__B2 core_0.decode.i_instr_l\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5520_ net57 _1556_ _1587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_146_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5146__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5451_ _1537_ _1540_ _1543_ _1545_ _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__5146__B2 _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8883__A2 _4383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6894__A1 core_0.execute.irq_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5697__A2 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6894__B2 core_0.execute.sreg_irq_flags.o_d\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8170_ net92 _3779_ _3797_ _3799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5382_ _1240_ _1281_ _1489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_239_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7121_ _1683_ _3047_ _3048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8635__A2 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_26_Left_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7052_ _1894_ _2979_ _2810_ _2980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_238_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4657__B1 _0686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6003_ core_0.execute.rf.reg_outputs\[1\]\[12\] _1779_ _1804_ core_0.execute.rf.reg_outputs\[11\]\[12\]
+ _1993_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_163_Right_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_241_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8399__A1 _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6247__C _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6949__A2 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7071__A1 core_0.execute.sreg_priv_control.o_d\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7954_ _3408_ _3672_ _3675_ _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_222_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5621__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6905_ _2709_ net216 _2836_ _2837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_166_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7885_ _3428_ _3628_ _3635_ _0383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9624_ _0634_ clknet_leaf_132_i_clk net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_176_2620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Left_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_147_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6836_ net78 _1411_ _2768_ core_0.execute.sreg_scratch.o_d\[1\] _2769_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_rebuffer52_I net279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7374__A2 _3293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5385__A1 _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9555_ _0565_ clknet_leaf_64_i_clk core_0.execute.sreg_irq_pc.o_d\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6767_ _2699_ _2700_ _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7873__I _3627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8506_ net84 _4040_ _4093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5718_ _1714_ _1716_ _0135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9486_ _0496_ clknet_leaf_21_i_clk net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_162_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7126__A2 _3040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6698_ _2635_ _2636_ _2637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_21_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5137__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8437_ _2230_ _4034_ _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ _1253_ _1660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_98_1688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6885__A1 _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5326__C _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8368_ _1542_ _1988_ _3980_ _3981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output166_I net166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7319_ _3209_ _2544_ _3240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_44_Left_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7822__B _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8299_ _1538_ _3915_ _3916_ _3917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_245_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_2760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6637__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8637__C _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_130_Right_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_244_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_125_2007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8653__B _4222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8372__C _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_2941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7269__B _3191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5612__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_wire215_I _0880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_107_1795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_218_3126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_6__f_i_clk_I clknet_3_3_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8562__A1 _4080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7365__A2 _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5376__A1 _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6876__A1 _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8828__B _4326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_229_3255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__C _2136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6628__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_229_3266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4639__B1 net347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_242_3411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_242_3422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5300__A1 net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_2276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7428__I0 core_0.ew_data\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5851__A2 net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput7 i_core_int_sreg[15] net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7053__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_2432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__A2 _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4951_ _1104_ _1113_ _1130_ _1131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_176_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7670_ core_0.execute.rf.reg_outputs\[13\]\[10\] _3504_ _3500_ _3511_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4882_ _0892_ net46 _1062_ _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_59_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8553__A1 _1175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6621_ net325 _2562_ _2563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_0_52_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5367__B2 _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9340_ _0350_ clknet_leaf_8_i_clk core_0.execute.rf.reg_outputs\[9\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6552_ _2453_ _2493_ _2494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5503_ _1058_ _1552_ _1578_ _0058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9271_ _0281_ clknet_leaf_149_i_clk core_0.execute.rf.reg_outputs\[14\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_232_Right_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_171_2561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6483_ net264 _1956_ _2425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_113_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8222_ core_0.execute.alu_mul_div.mul_res\[2\] _3846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6867__A1 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6867__B2 _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9379__CLK clknet_leaf_7_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5434_ _1267_ _1274_ _1271_ _1437_ _1530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_168_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8153_ net99 _3787_ _3785_ _3790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5365_ _1464_ _1477_ _0020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6619__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7104_ _2931_ _3030_ _2570_ _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_239_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_227_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8084_ core_0.execute.rf.reg_outputs\[2\]\[9\] _3743_ _3745_ _3750_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5296_ core_0.execute.prev_sys _0899_ _1417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__7292__A1 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6095__A2 _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ _2703_ _2963_ _2964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7292__B2 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_198_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5842__A2 net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7044__A1 _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8986_ core_0.dec_rf_ie\[4\] _1482_ _1462_ _1480_ _4461_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8192__C _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7595__A2 core_0.ew_data\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8792__A1 _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7937_ _3457_ _3652_ _3665_ _0405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5388__I _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7868_ core_0.execute.rf.reg_outputs\[8\]\[14\] _3605_ _3621_ _3625_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8544__A1 net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9607_ _0617_ clknet_leaf_51_i_clk core_0.execute.pc_high_buff_out\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6819_ _1880_ _2748_ _2752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5358__B2 _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7799_ _3584_ _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_46_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9538_ _0548_ clknet_leaf_73_i_clk net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_107_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9469_ _0479_ clknet_leaf_50_i_clk core_0.execute.rf.reg_outputs\[1\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4581__A2 _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_213_3067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6858__A1 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5530__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5833__A2 _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4892__I0 net62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7035__A1 _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_224_3196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7586__A2 _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5597__A1 _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5298__I core_0.dec_sreg_store vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_196_2859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7338__A2 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8535__A1 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5349__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7727__B _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6631__B _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6010__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_19_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_2305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5150_ _1267_ _1302_ _1303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7274__A1 _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6793__S _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ core_0.decode.i_instr_l\[4\] _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_236_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_224_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5824__A2 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8840_ core_0.execute.pc_high_buff_out\[5\] _4335_ _4364_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7026__B2 net12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7577__A2 _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8771_ _0765_ _4295_ _4309_ _4307_ _0595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5588__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9051__CLK clknet_leaf_92_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5983_ _0714_ _1962_ _1965_ _1972_ _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_59_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7722_ core_0.ew_reg_ie\[11\] _3395_ _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_47_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4934_ core_0.fetch.prev_request_pc\[3\] _1060_ _1063_ core_0.fetch.prev_request_pc\[2\]
+ _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_176_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8526__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7329__A2 _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8526__B2 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7637__B _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7653_ core_0.execute.rf.reg_outputs\[13\]\[2\] _3498_ _3500_ _3502_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4865_ _1017_ net53 _1045_ _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_90_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_12 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6604_ net237 _2546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _3456_ _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_145_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4796_ _0949_ _0970_ _0976_ _0977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9323_ _0333_ clknet_leaf_0_i_clk core_0.execute.rf.reg_outputs\[10\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6535_ _2143_ _2370_ _2477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8829__A2 _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4563__A2 _0682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5760__A1 _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9254_ _0264_ clknet_leaf_150_i_clk core_0.execute.rf.reg_outputs\[15\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6466_ _2413_ _0914_ _0186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_rebuffer15_I _0848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7501__A2 _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8205_ core_0.execute.alu_mul_div.mul_res\[0\] _3830_ _3831_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5417_ _1231_ _1297_ _1515_ _0034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput130 net130 o_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9185_ _0196_ clknet_leaf_47_i_clk net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput141 net141 o_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6397_ _1988_ _2371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XANTENNA_clkbuf_4_12__f_i_clk_I clknet_3_6_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput152 net152 o_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput163 net163 o_req_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_100_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput174 net174 o_req_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8136_ core_0.ew_reg_ie\[0\] _3394_ _3779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_227_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5348_ core_0.decode.i_instr_l\[8\] _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA_input42_I i_req_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput185 net185 sr_bus_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_195_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput196 net196 sr_bus_data_o[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_227_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7265__A1 _2480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6068__A2 _1791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8067_ _3408_ _3737_ _3740_ _0460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5279_ _0995_ _1005_ _1399_ _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_227_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7018_ _2501_ _2946_ core_0.decode.oc_alu_mode\[4\] _2947_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_3_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8765__A1 core_0.execute.sreg_scratch.o_d\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8969_ _1440_ _1230_ _1272_ _4452_ _0650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_78_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8517__A1 _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8650__C _4219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7039__S _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8222__I core_0.execute.alu_mul_div.mul_res\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwire213 _1911_ net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_18_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7740__A2 _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_20_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5751__A1 _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4554__A2 _0673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_239_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6700__B1 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_3225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6059__A2 _1801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5806__A2 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7008__A1 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4925__I core_0.fetch.prev_request_pc\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4490__A1 core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7559__A2 _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8756__A1 net243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8508__A1 _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8560__C _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_237_3354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5990__A1 core_0.execute.rf.reg_outputs\[6\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5990__B2 core_0.execute.rf.reg_outputs\[12\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4650_ core_0.execute.rf.reg_outputs\[11\]\[4\] _0680_ _0705_ core_0.execute.rf.reg_outputs\[9\]\[4\]
+ _0837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7731__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 i_core_int_sreg[3] net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput21 i_mem_data[0] net21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4545__A2 _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_2375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput32 i_mem_data[5] net32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4581_ core_0.execute.rf.reg_outputs\[15\]\[10\] _0702_ _0715_ _0774_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput43 i_req_data[14] net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_141_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5742__B2 _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput54 i_req_data[25] net54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6320_ core_0.execute.alu_mul_div.div_cur\[11\] _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput65 i_req_data[6] net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6251_ core_0.execute.alu_mul_div.div_cur\[2\] _2009_ _2238_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_122_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5202_ _0896_ _1146_ _1344_ _1345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_0_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6182_ core_0.execute.alu_mul_div.div_cur\[0\] _1875_ _2171_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_237_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _1231_ _1284_ _1287_ _0010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7920__B _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8735__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5064_ _0908_ net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_74_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4481__A1 _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8747__A1 _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8823_ core_0.execute.pc_high_out\[3\] _4342_ _4349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_36_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Left_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_8754_ _4293_ _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5966_ _1944_ _1955_ _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__7970__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7705_ core_0.execute.rf.reg_outputs\[12\]\[8\] _3526_ _3528_ _3532_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4917_ _1095_ _1096_ _1097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8685_ _1658_ _4245_ _4248_ _0570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_176_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5981__A1 core_0.execute.rf.reg_outputs\[1\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4784__A2 _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5981__B2 core_0.execute.rf.reg_outputs\[11\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5897_ core_0.decode.oc_alu_mode\[1\] core_0.decode.oc_alu_mode\[6\] core_0.decode.oc_alu_mode\[7\]
+ core_0.decode.oc_alu_mode\[4\] _1887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_164_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7636_ _3460_ _3477_ _3491_ _0278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4848_ _0893_ net52 _1028_ _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_62_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7722__A2 _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7567_ net27 _1347_ _3443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_172_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4536__A2 _0698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4779_ core_0.dec_l_reg_sel\[1\] core_0.dec_l_reg_sel\[0\] _0960_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_105_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5584__I1 core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9306_ _0316_ clknet_leaf_1_i_clk core_0.execute.rf.reg_outputs\[11\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6518_ _1846_ net213 _2460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_210_3037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7498_ _2709_ _2422_ _3383_ _0248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9237_ _0248_ clknet_leaf_44_i_clk core_0.ew_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6449_ _1180_ _2386_ _2407_ _0175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_219_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9168_ _0179_ clknet_leaf_104_i_clk core_0.execute.mem_stage_pc\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8119_ core_0.execute.rf.reg_outputs\[1\]\[8\] _3765_ _3756_ _3770_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_209_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7830__B _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9099_ _0124_ clknet_leaf_43_i_clk net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7789__A2 _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6446__B _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6461__A2 _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_221_3166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8661__B _1709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7410__A1 _2795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7961__A2 _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_193_2829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4775__A2 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7713__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8910__A1 _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__A2 net302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5724__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_3295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_2_i_clk clknet_4_2__leaf_i_clk clknet_leaf_2_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_131_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7740__B _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6452__A2 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7401__A1 _3073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5820_ _1789_ _1795_ _1800_ _1809_ _1810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_159_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7952__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5751_ _1736_ _1739_ _1740_ _1741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4702_ _0881_ _0882_ _0883_ _0884_ _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_8470_ _4047_ _4057_ _4061_ _4062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5682_ net186 _1687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_155_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8901__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7704__A2 _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7421_ _1684_ core_0.execute.sreg_irq_pc.o_d\[15\] _3340_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_13_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4633_ core_0.execute.rf.reg_outputs\[15\]\[6\] _0702_ _0715_ _0822_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7352_ _3262_ _3272_ core_0.dec_mem_access _3273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4564_ _0754_ _0755_ _0756_ _0757_ _0758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5191__A2 _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6303_ core_0.execute.alu_mul_div.div_cur\[8\] _2218_ _0999_ _2285_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7283_ core_0.ew_data\[11\] _3205_ _0199_ _3206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4495_ _0692_ _0693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_40_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9022_ _0049_ clknet_leaf_79_i_clk core_0.fetch.out_buffer_data_instr\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6234_ _2141_ _2174_ _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_168_2533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6140__A1 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6691__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6165_ _2144_ _2147_ _2150_ _2153_ _2154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5116_ _1234_ _1269_ _1270_ _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_176_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6096_ core_0.execute.rf.reg_outputs\[13\]\[3\] _0954_ _0955_ _0980_ _2086_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_240_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7640__A1 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5047_ core_0.fetch.prev_request_pc\[3\] _1148_ _1215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7491__I1 core_0.ew_reg_ie\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer82_I net309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8196__A2 _3821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6780__I core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8806_ _4322_ _1400_ _1414_ _4334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_79_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6998_ core_0.ew_data\[4\] _2642_ _2928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_2662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7943__A2 _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7097__B core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5954__A1 net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5949_ core_0.execute.rf.reg_outputs\[15\]\[10\] _0945_ _1821_ core_0.execute.rf.reg_outputs\[7\]\[10\]
+ _1938_ _1939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_8737_ core_0.execute.trap_flag _1418_ _4289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8668_ _4212_ core_0.execute.mem_stage_pc\[5\] _4201_ _4234_ _4235_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_164_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output196_I net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7619_ _3475_ _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_63_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4509__A2 _0675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5706__A1 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8599_ net201 _4165_ _4174_ _4175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclone68 _0682_ net296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_172_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_160_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5182__A2 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_177_Right_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_160_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8120__A2 _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6020__I _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output73_I net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4693__B2 core_0.execute.rf.reg_outputs\[10\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8423__A3 _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6434__A2 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__I _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_205_2972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8187__A2 _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__A2 _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_183_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4748__A2 _0928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_1993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_234_3324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9262__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_2334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5173__A2 _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_144_Right_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8111__A2 _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_150_i_clk clknet_4_0__leaf_i_clk clknet_leaf_150_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6122__A1 core_0.execute.rf.reg_outputs\[5\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6122__B2 core_0.execute.rf.reg_outputs\[3\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6673__A2 _2614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7870__A1 core_0.execute.rf.reg_outputs\[8\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_3453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_142_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6425__A2 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7970_ _3450_ _3672_ _3684_ _0419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7473__I1 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_2463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_163_2474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _2349_ _2755_ _2442_ _1885_ _2852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_233_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6852_ _1401_ _2767_ _2783_ _2784_ _2785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_9640_ _0650_ clknet_leaf_138_i_clk core_0.dec_jump_cond_code\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6189__A1 core_0.execute.alu_mul_div.div_cur\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6189__B2 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7925__A2 _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5803_ _0971_ _0943_ _0950_ _1793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_9571_ _0581_ clknet_leaf_45_i_clk net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_147_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4739__A2 _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5936__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6783_ _1857_ _1974_ _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_71_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8522_ net85 _4099_ _4107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5734_ _1726_ _1699_ _1727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_99_Left_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_103_i_clk clknet_4_13__leaf_i_clk clknet_leaf_103_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8453_ _1420_ _1735_ _4046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7689__A1 core_0.execute.rf.reg_outputs\[12\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5665_ _1545_ _1534_ _1673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8350__A2 _3830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7404_ _1883_ _2599_ _3322_ _2571_ _3323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_44_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4616_ _0802_ _0803_ _0804_ _0805_ _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8384_ _3993_ _3995_ _3996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5164__A2 _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_67_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5596_ _1591_ _1567_ _1630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_111_Right_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7335_ _1326_ _3242_ _3252_ _3255_ _3256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4911__A2 _1020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4547_ net90 _0742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_118_i_clk clknet_4_7__leaf_i_clk clknet_leaf_118_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8102__A2 _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6113__A1 _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7266_ _2713_ _3188_ _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4478_ _0660_ _0663_ core_0.dec_r_reg_sel\[1\] _0675_ _0676_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_111_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9005_ _0032_ clknet_leaf_135_i_clk core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6775__I core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6217_ core_0.execute.alu_mul_div.div_cur\[15\] net239 _2193_ _2205_ _2206_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_217_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7197_ core_0.execute.sreg_priv_control.o_d\[9\] _1693_ _2996_ net16 _2689_ _3122_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_51_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ _2130_ _2133_ _2137_ _2138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_225_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6079_ net99 _1771_ _2059_ _2068_ _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__6967__A3 _2896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8169__A2 _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output111_I net111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output209_I net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5227__I0 core_0.ew_data\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7377__B1 _3295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7916__A2 _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_246_Right_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8964__I1 core_0.decode.i_imm_pass\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5927__A1 core_0.execute.rf.reg_outputs\[5\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5927__B2 core_0.execute.rf.reg_outputs\[10\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5059__C _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__A2 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A2 _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6104__B2 core_0.execute.rf.reg_outputs\[1\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_82_i_clk clknet_4_14__leaf_i_clk clknet_leaf_82_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6655__A2 _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7852__A1 _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4666__A1 core_0.execute.rf.reg_outputs\[7\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6407__A2 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7604__B2 net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7080__A2 net289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_97_i_clk clknet_4_13__leaf_i_clk clknet_leaf_97_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_203_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_240_3394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5091__B2 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6353__C _2229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_213_Right_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5918__A1 core_0.execute.rf.reg_outputs\[4\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_20_i_clk clknet_4_6__leaf_i_clk clknet_leaf_20_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_129_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8580__A2 _2949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6591__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5394__A2 _1488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8332__A2 _3947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_35_i_clk clknet_4_8__leaf_i_clk clknet_leaf_35_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7184__C _3073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5450_ _1544_ _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_26_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5146__A2 _1297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__A1 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6894__A2 _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5381_ _1320_ _1324_ _1448_ _1487_ _1488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_151_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7120_ net84 _2995_ _3046_ _2893_ _3047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7051_ _2010_ _2801_ _2979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7843__A1 _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4657__A1 core_0.execute.rf.reg_outputs\[5\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6002_ core_0.execute.rf.reg_outputs\[6\]\[12\] net322 _1819_ core_0.execute.rf.reg_outputs\[12\]\[12\]
+ _1788_ core_0.execute.rf.reg_outputs\[3\]\[12\] _1992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_5_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4657__B2 core_0.execute.rf.reg_outputs\[14\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7446__I1 _3085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5004__I net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7071__A2 _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7953_ core_0.execute.rf.reg_outputs\[5\]\[1\] _3673_ _3663_ _3675_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5082__A1 core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ _2708_ _2835_ _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7884_ core_0.execute.rf.reg_outputs\[7\]\[4\] _3634_ _3621_ _3635_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_221_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8020__A1 _3469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9623_ _0633_ clknet_leaf_66_i_clk core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_176_2621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6835_ _1686_ net227 _2683_ _2768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_0_159_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6766_ _2673_ _2698_ _2700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9554_ _0564_ clknet_4_9__leaf_i_clk core_0.execute.sreg_irq_pc.o_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer45_I core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8505_ net84 _4091_ _4092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4593__B1 _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5717_ core_0.execute.sreg_priv_control.o_d\[7\] _1701_ _1715_ _1698_ _1716_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6697_ _2629_ _2630_ net210 _2622_ _2636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_17_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9485_ _0495_ clknet_leaf_23_i_clk net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_21_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8050__I _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5648_ _1658_ _1595_ _1086_ _0122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_33_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8436_ _4020_ _4031_ core_0.execute.alu_mul_div.div_res\[11\] _4034_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5137__A2 _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6334__A1 _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8367_ _1542_ _1999_ _3980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6885__A2 core_0.execute.alu_mul_div.mul_res\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5579_ _1242_ core_0.fetch.submitable _1620_ _0092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7318_ _2839_ _3238_ _3239_ _0212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8087__A1 _3456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8298_ _1538_ _3866_ _3916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7834__A1 core_0.ew_reg_ie\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6637__A2 _2578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_2761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7249_ _3171_ _2465_ _3172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_229_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__A1 net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4954__S _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8653__C _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7062__A2 core_0.execute.alu_mul_div.mul_res\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6454__B _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5849__I net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_202_2931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_202_2942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4820__A1 _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_107_1796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_218_3127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8562__A2 _3297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6325__A1 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_229_3256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7825__A1 _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4639__A1 core_0.execute.rf.reg_outputs\[6\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5836__B1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4639__B2 core_0.execute.rf.reg_outputs\[15\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_242_3412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5300__A2 net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9450__CLK clknet_leaf_136_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_2277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput8 i_core_int_sreg[1] net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8563__C _2136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7053__A2 _2487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_2433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5759__I _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4950_ core_0.fetch.prev_request_pc\[0\] _1054_ _1130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6800__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6083__C _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4811__A1 _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4881_ _0892_ _1061_ _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6620_ _2008_ _2561_ _1769_ _2562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_7_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5367__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__A1 _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6551_ net343 _2492_ _2493_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4575__B1 _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5502_ net47 _1554_ _1578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9270_ _0280_ clknet_leaf_151_i_clk core_0.execute.rf.reg_outputs\[14\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6482_ net264 _1956_ _2424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5427__C _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6316__A1 _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_171_2562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8221_ _3832_ _3844_ _3845_ _0509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5433_ _1232_ _1233_ _1240_ _1288_ _1529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__7923__B _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4878__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8069__A1 _3414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8152_ _3434_ _3780_ _3789_ _0496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_168_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5364_ core_0.dec_rf_ie\[10\] _1438_ _1472_ _1476_ _1477_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_239_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6539__B _2480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_227_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7103_ _1769_ _3029_ net267 _3030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_8083_ _3450_ _3737_ _3749_ _0467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5295_ _1397_ _1415_ _1416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_227_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7034_ _2897_ _2961_ _2963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6095__A3 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_182_2691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5055__A1 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8985_ _1497_ _4460_ _0658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_210_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7936_ core_0.execute.rf.reg_outputs\[6\]\[10\] _3657_ _3663_ _3665_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_210_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A1 core_0.ew_reg_ie\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4802__B2 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7867_ _3466_ _3607_ _3624_ _0376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6004__B1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9606_ _0616_ clknet_leaf_51_i_clk core_0.execute.pc_high_buff_out\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5358__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6818_ _1338_ _2341_ _1285_ _2751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7798_ _3584_ _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_9_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4566__B1 _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9537_ _0547_ clknet_leaf_77_i_clk net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_80_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6749_ _1690_ net177 _1409_ _2683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_162_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9468_ _0478_ clknet_leaf_25_i_clk core_0.execute.rf.reg_outputs\[1\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_104_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_213_3068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8419_ _2921_ _4023_ _2258_ _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4869__A1 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9399_ _0409_ clknet_leaf_148_i_clk core_0.execute.rf.reg_outputs\[6\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5530__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_131_2089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7807__A1 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9473__CLK clknet_leaf_37_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_218_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8480__A1 _1211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5294__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6963__I _2694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_109_1825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8232__A1 core_0.execute.alu_mul_div.cbit\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5046__A1 _1211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_244_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5597__A2 net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8535__A2 _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5349__A2 _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8471__A1 _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5080_ _1234_ _1236_ _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5285__A1 net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7026__A2 _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_204_Left_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4607__B _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8774__A2 _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5982_ _1813_ _1966_ _1967_ _1971_ _1972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8770_ core_0.execute.sreg_scratch.o_d\[11\] _4300_ _4309_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5588__A2 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4933_ core_0.fetch.prev_request_pc\[1\] _1043_ _1113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7721_ _3473_ _3521_ _3540_ _0314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7918__B _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8526__A2 _4048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4864_ _1017_ _1044_ _1045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6537__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7652_ _3409_ _3497_ _3501_ _0284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_13 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4548__B1 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6603_ _2544_ _2545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7583_ _3387_ core_0.ew_data\[10\] _3449_ net22 _3456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_28_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4795_ _0972_ _0973_ _0974_ _0975_ _0949_ _0976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5060__I1 _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6534_ _2468_ _2469_ _2472_ _2475_ _2476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_9322_ _0332_ clknet_leaf_1_i_clk core_0.execute.rf.reg_outputs\[10\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5760__A2 net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_213_Left_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7653__B _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6465_ _2413_ _0917_ _0185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9253_ _0263_ clknet_leaf_1_i_clk core_0.execute.rf.reg_outputs\[15\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5952__I _1941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8204_ _3829_ _3830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
X_5416_ core_0.dec_alu_carry_en _1286_ _1515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput120 net120 o_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9184_ _0195_ clknet_leaf_47_i_clk net134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7372__C _1768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput131 net131 o_mem_addr_high[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5512__A2 _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6396_ _1973_ _2370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
Xoutput142 net142 o_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_63_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput153 net153 o_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8135_ _3472_ _3760_ _3778_ _0490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput164 net164 o_req_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5347_ _1253_ _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput175 net175 o_req_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput186 net186 sr_bus_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput197 net294 sr_bus_data_o[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_184_2720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8462__A1 net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8066_ core_0.execute.rf.reg_outputs\[2\]\[1\] _3738_ _3730_ _3740_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5278_ core_0.decode.i_flush _1398_ _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input35_I i_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5901__B _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7017_ _2434_ _2903_ _2946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_3_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8765__A2 _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8968_ core_0.dec_jump_cond_code\[0\] _1250_ _4452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5579__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7828__B _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7919_ _3415_ _3651_ _3655_ _0397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8899_ _1253_ _2380_ _1228_ _0621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_104_1766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6528__A1 net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwire214 _2069_ net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_190_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5503__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6700__A1 core_0.execute.rf.reg_outputs\[7\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6700__B2 core_0.execute.rf.reg_outputs\[5\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_1895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_226_3226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8453__A1 _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5806__A3 _0951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8205__A1 core_0.execute.alu_mul_div.mul_res\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7008__A2 _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4490__A2 _0664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8756__A2 _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__A1 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7738__B _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_237_3355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5990__A2 net322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_62_Left_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_127_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput11 i_core_int_sreg[4] net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput22 i_mem_data[10] net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4580_ core_0.execute.rf.reg_outputs\[14\]\[10\] _0685_ _0699_ core_0.execute.rf.reg_outputs\[12\]\[10\]
+ _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_142_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_155_2376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5742__A2 _1700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput33 i_mem_data[6] net33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput44 i_req_data[16] net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput55 i_req_data[26] net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput66 i_req_data[7] net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7192__C _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6250_ _2219_ _2236_ _2237_ _2229_ _0146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_110_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8692__A1 _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5201_ _0896_ _1343_ _1344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6181_ core_0.execute.alu_mul_div.div_cur\[1\] _1895_ _2170_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_110_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5132_ _1285_ _1286_ _1287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8444__A1 _1680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Left_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_90_1589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5063_ _1086_ _1225_ _1227_ _1162_ net160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_165_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4481__A2 net298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8747__A2 _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8822_ _4316_ _4348_ _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6758__A1 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8751__C _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7648__B _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8753_ _0859_ _4294_ _4299_ _4287_ _0587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5965_ _1947_ _1949_ _1954_ _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_181_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4851__I _1031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7704_ _3447_ _3520_ _3531_ _0306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4916_ core_0.fetch.prev_request_pc\[8\] _1046_ _1049_ core_0.fetch.prev_request_pc\[9\]
+ _1096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_176_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8684_ _4212_ core_0.execute.mem_stage_pc\[8\] _4201_ _4247_ _4248_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5896_ core_0.decode.oc_alu_mode\[9\] core_0.decode.oc_alu_mode\[11\] core_0.decode.oc_alu_mode\[3\]
+ _1337_ _1886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_118_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_158_Right_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5981__A2 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7635_ core_0.execute.rf.reg_outputs\[14\]\[11\] _3482_ _3486_ _3491_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4847_ _0893_ _1027_ _1028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7183__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7566_ _3397_ _3441_ _3442_ _0257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_137_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6930__A1 _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4778_ _0957_ _0958_ _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_7_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6778__I _2710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9305_ _0315_ clknet_leaf_3_i_clk core_0.execute.rf.reg_outputs\[11\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6517_ _2432_ _2441_ _2455_ _2458_ _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_132_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_210_3027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_2790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4800__B _0980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5682__I net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7497_ _3382_ _2419_ _3383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_210_3038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8683__A1 _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9236_ _0247_ clknet_leaf_143_i_clk core_0.ew_reg_ie\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6448_ core_0.execute.mem_stage_pc\[11\] _2395_ _2404_ _2407_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_8_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6379_ _2344_ _2352_ _2140_ _2353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9167_ _0178_ clknet_leaf_102_i_clk core_0.execute.mem_stage_pc\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7238__A2 _3156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8118_ _3446_ _3759_ _3769_ _0482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_54_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9098_ _0123_ clknet_leaf_101_i_clk core_0.fetch.pc_reset_override vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_243_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8986__A2 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8049_ _3456_ _3716_ _3729_ _0453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6997__A1 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8738__A2 _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_221_3167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6749__A1 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8661__C _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7558__B _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_119_Left_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7410__A2 _3314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_210_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_125_Right_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8910__A2 _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6921__A1 _2349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6921__B2 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_3296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_128_Left_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8674__A1 _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5488__A1 net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8426__A1 _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6637__B _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8977__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6988__A1 _2759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8729__A2 _4283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_137_Left_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_159_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5412__A1 core_0.decode.i_instr_l\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5412__B2 core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5750_ _1704_ _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_146_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5963__A2 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4701_ core_0.execute.rf.reg_outputs\[9\]\[0\] _0705_ net257 core_0.execute.rf.reg_outputs\[8\]\[0\]
+ _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_17_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5681_ net185 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_60_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7420_ net77 _2995_ _3338_ _2893_ _3339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4632_ core_0.execute.rf.reg_outputs\[14\]\[6\] net310 net308 core_0.execute.rf.reg_outputs\[1\]\[6\]
+ _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_13_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6912__A1 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7351_ _3234_ _3269_ _3271_ _3272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4563_ core_0.execute.rf.reg_outputs\[7\]\[11\] _0682_ _0697_ core_0.execute.rf.reg_outputs\[3\]\[11\]
+ _0757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_114_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_146_Left_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4620__B _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6302_ _2220_ _2282_ _2283_ _2284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7282_ net305 _3204_ _2708_ _3205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4494_ net348 _0675_ _0671_ _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_92_1618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9021_ _0048_ clknet_leaf_78_i_clk core_0.fetch.out_buffer_data_instr\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_228_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7931__B _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6233_ _2170_ _2171_ _2222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_168_2523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_2534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6164_ _2151_ _2152_ _2153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_237_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8968__A2 _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5115_ core_0.decode.i_instr_l\[3\] core_0.decode.i_instr_l\[2\] _1270_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_225_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6095_ core_0.execute.rf.reg_outputs\[14\]\[3\] _0957_ _0958_ _0980_ _2085_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_209_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6979__A1 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_227_Right_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5046_ _1211_ _1165_ _1213_ _1214_ _1080_ net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__7640__A2 _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_63_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_212_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8805_ _4316_ _4333_ _0605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_138_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6997_ _2672_ net203 _2926_ _2927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_165_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_179_2663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8736_ _4288_ _0581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_220_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5948_ _1935_ _1936_ _1937_ _1938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5954__A2 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_101_1725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8667_ _4203_ _4077_ _4233_ _1661_ _4234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_35_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ _1519_ _1868_ _1869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_90_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7618_ _3421_ _3476_ _3481_ _0270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6903__A1 _2710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8598_ _3330_ _4165_ _4174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output189_I net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7549_ _3427_ _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8002__B _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_160_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8656__A1 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4957__S _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9219_ _0230_ clknet_leaf_82_i_clk net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_1854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8656__C _4205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8408__A1 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6457__B _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4693__A2 net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7631__A2 _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_2206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_205_2973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7288__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__A2 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_211_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A2 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_3325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7147__A1 core_0.decode.oc_alu_mode\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6920__B _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8895__A1 net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_2335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5028__S _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9557__CLK clknet_leaf_74_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7751__B _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6122__A2 _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7870__A2 _3605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_3454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5881__A1 _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7622__A2 _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_163_2464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5633__A1 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6920_ _1338_ _2349_ _1285_ _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_89_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6851_ _1401_ core_0.execute.sreg_irq_pc.o_d\[1\] _2784_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7386__A1 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6189__A2 _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _1791_ _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_147_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9570_ _0580_ clknet_leaf_62_i_clk core_0.execute.sreg_jtr_buff.o_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5936__A2 _1925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6782_ _1875_ _1973_ _2714_ _1897_ _2715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_92_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8521_ _4103_ _4106_ _4051_ _0548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5733_ net197 _1726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_17_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6830__B core_0.execute.alu_mul_div.i_div vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_154_Left_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8886__A1 _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8452_ _4039_ _4044_ _4045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7689__A2 _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5664_ _1001_ _1534_ _1672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_115_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7403_ net270 _2595_ _1883_ _3322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4615_ core_0.execute.rf.reg_outputs\[7\]\[7\] net297 _0697_ core_0.execute.rf.reg_outputs\[3\]\[7\]
+ _0805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8383_ _3994_ _3988_ _3995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5595_ core_0.decode.i_instr_l\[11\] _1628_ _1629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8638__A1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4546_ _0741_ net197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7334_ _3248_ _3253_ _3254_ _3255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_41_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7310__A1 _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7265_ _2480_ _3172_ _3187_ _3188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__6113__A2 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4477_ _0664_ _0675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_96_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9004_ _0031_ clknet_leaf_133_i_clk core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_111_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6216_ _2194_ _2195_ _2204_ _2205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_217_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7196_ core_0.execute.sreg_irq_pc.o_d\[9\] _3042_ _3044_ core_0.execute.sreg_scratch.o_d\[9\]
+ _3121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_216_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_51_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4675__A2 _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _0890_ _2134_ _2135_ _2136_ _2137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_163_Left_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_209_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8810__A1 _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7613__A2 _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6078_ _2060_ _2061_ _2062_ _2067_ _2068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_213_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5029_ net84 _1085_ _1201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_200_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7377__A1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7377__B2 _3296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5227__I1 core_0.ew_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output104_I net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_1_i_clk clknet_4_0__leaf_i_clk clknet_leaf_1_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5927__A2 net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8719_ core_0.execute.sreg_irq_pc.o_d\[14\] _4210_ _1431_ _4277_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7129__A1 core_0.ew_data\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8877__A1 core_0.execute.pc_high_buff_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_216_3099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__A2 _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8629__A1 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5560__B1 _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6104__A2 _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7852__A2 _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A2 _0683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5863__A1 net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7604__A2 core_0.ew_data\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8801__A1 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5615__A1 core_0.decode.i_imm_pass\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_240_3395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5091__A2 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5918__A2 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8868__A1 net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5551__B1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5380_ _1289_ _1298_ _1269_ _1487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7050_ _2010_ _2802_ _2977_ _2075_ _2978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_238_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7843__A2 _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6001_ _1989_ _1990_ _1991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A1 net287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4657__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7952_ _3401_ _3672_ _3674_ _0411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_179_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _2710_ _2821_ _2834_ _2835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7883_ _3627_ _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__8556__B1 net294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9622_ _0632_ clknet_leaf_132_i_clk core_0.dec_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6834_ _2694_ net78 _2767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8020__A2 _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_2622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9553_ _0563_ clknet_leaf_68_i_clk core_0.execute.sreg_irq_pc.o_d\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6765_ core_0.dec_sreg_load _2673_ _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_147_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8504_ net83 net82 _4076_ _4091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_174_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8859__A1 _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7375__C core_0.execute.alu_mul_div.i_div vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ net278 _1704_ _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_9484_ _0494_ clknet_leaf_17_i_clk net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6696_ _2627_ _2634_ _2635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_rebuffer38_I net264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8435_ _3153_ _4033_ _2258_ _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5647_ _1658_ _0896_ _1659_ _0121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_32_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8366_ _3966_ _3972_ _3979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5578_ _1073_ core_0.fetch.submitable _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_60_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input65_I i_req_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7317_ core_0.ew_data\[12\] _3168_ _3239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4529_ core_0.execute.rf.reg_outputs\[15\]\[14\] net347 _0705_ core_0.execute.rf.reg_outputs\[9\]\[14\]
+ _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8087__A2 _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8297_ _2362_ _2346_ _1544_ _3915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_187_2751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8492__C1 _2954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_2762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7248_ _3143_ _3134_ _3171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7834__A2 _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__A2 _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5845__A1 net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7179_ _2571_ net334 _3103_ _3104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_217_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9252__CLK clknet_leaf_3_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6270__A1 core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5073__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_202_2932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8547__B1 net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8011__A2 _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_218_3128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A1 core_0.execute.rf.reg_outputs\[7\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7770__A1 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4584__A1 net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7522__A1 _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8078__A2 _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8322__I0 core_0.execute.alu_mul_div.mul_res\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__A1 core_0.execute.rf.reg_outputs\[12\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_229_3257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7825__A2 _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4639__A2 _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5836__B2 core_0.execute.rf.reg_outputs\[7\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_242_3413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5300__A3 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_2278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_102_i_clk clknet_4_13__leaf_i_clk clknet_leaf_102_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput9 i_core_int_sreg[2] net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_188_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_160_2434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8860__B _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4811__A2 _0946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_117_i_clk clknet_4_7__leaf_i_clk clknet_leaf_117_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8002__A2 _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4880_ core_0.fetch.out_buffer_data_instr\[18\] _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6013__A1 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6550_ net218 _2492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_15_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5501_ _1061_ _1551_ _1577_ _0057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7108__A4 _3034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7513__A1 core_0.ew_reg_ie\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6481_ _2143_ _2370_ _2423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_171_2563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8220_ core_0.execute.alu_mul_div.mul_res\[1\] _3832_ _3845_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5432_ _1247_ _1279_ _1288_ _1528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_152_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5363_ core_0.decode.i_instr_l\[9\] _1465_ core_0.decode.i_instr_l\[7\] _1476_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__8069__A2 _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8151_ net98 _3787_ _3785_ _3789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _1883_ _2360_ _3028_ _3029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7816__A2 _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5294_ _1400_ _1414_ _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_8082_ core_0.execute.rf.reg_outputs\[2\]\[8\] _3743_ _3745_ _3749_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_168_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7033_ _2897_ _2961_ _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6095__A4 _0980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_182_2692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8984_ core_0.dec_rf_ie\[3\] _1482_ _1462_ _1478_ _4460_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_93_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5055__A2 _1220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7935_ _3454_ _3651_ _3664_ _0404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_210_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4802__A2 _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7866_ core_0.execute.rf.reg_outputs\[8\]\[13\] _3613_ _3621_ _3624_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6004__A1 core_0.execute.rf.reg_outputs\[5\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_9605_ _0615_ clknet_leaf_50_i_clk core_0.execute.pc_high_buff_out\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6004__B2 core_0.execute.rf.reg_outputs\[14\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6817_ _2480_ _2749_ _2750_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_175_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7752__A1 _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7797_ core_0.ew_reg_ie\[9\] _3395_ _3584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5685__I net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_81_i_clk clknet_4_14__leaf_i_clk clknet_leaf_81_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_163_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9536_ _0546_ clknet_leaf_76_i_clk net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_135_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6748_ core_0.execute.sreg_priv_control.o_d\[0\] _1405_ net227 _2680_ _2682_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_18_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9467_ _0477_ clknet_leaf_48_i_clk core_0.execute.rf.reg_outputs\[1\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6679_ _2618_ _2619_ _2620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_213_3069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8418_ _4015_ _4022_ _4023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9398_ _0408_ clknet_leaf_149_i_clk core_0.execute.rf.reg_outputs\[6\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_96_i_clk clknet_4_13__leaf_i_clk clknet_leaf_96_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4869__A2 _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output171_I net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8349_ _2366_ _3833_ _3963_ _3828_ _3964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_103_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5530__A3 _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7807__A2 _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6491__A1 _1745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__A2 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4764__I _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8232__A2 _3854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_224_3198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5046__A2 _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_100_Left_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_240_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_200_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7296__B _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_49_i_clk clknet_4_10__leaf_i_clk clknet_leaf_49_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5349__A3 core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6546__A2 _2487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7743__A1 _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8299__A2 _3915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6482__A1 net264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5285__A2 net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_10_Right_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_223_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4674__I net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_139_Right_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6234__A1 _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5981_ core_0.execute.rf.reg_outputs\[1\]\[14\] _1779_ _1804_ core_0.execute.rf.reg_outputs\[11\]\[14\]
+ _1970_ _1971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_151_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7720_ core_0.execute.rf.reg_outputs\[12\]\[15\] _3519_ _3539_ _3540_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4932_ core_0.fetch.prev_request_pc\[2\] _1063_ _1112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5993__B1 _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7651_ core_0.execute.rf.reg_outputs\[13\]\[1\] _3498_ _3500_ _3501_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4863_ core_0.fetch.out_buffer_data_instr\[24\] _1044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_170_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_157_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6537__A2 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7734__A1 core_0.execute.rf.reg_outputs\[11\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_14 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6602_ _2472_ _2543_ _2544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_157_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4548__B2 core_0.execute.rf.reg_outputs\[9\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7582_ _3397_ _3454_ _3455_ _0260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4794_ core_0.ew_reg_ie\[5\] _0963_ _0964_ core_0.ew_reg_ie\[6\] _0948_ core_0.ew_reg_ie\[4\]
+ _0975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_90_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9321_ _0331_ clknet_leaf_3_i_clk core_0.execute.rf.reg_outputs\[10\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6533_ _2473_ _2474_ _2475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__B _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8749__C _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9252_ _0262_ clknet_leaf_3_i_clk core_0.execute.rf.reg_outputs\[15\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6464_ _2413_ _0912_ _0184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_1649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8203_ _3828_ _3821_ _3829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput110 net110 o_instr_long_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5415_ _0971_ _1486_ _1514_ _1501_ _0033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_112_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9183_ _0194_ clknet_leaf_46_i_clk net133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput121 net121 o_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6395_ _1544_ _2368_ _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput132 net132 o_mem_addr_high[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_101_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput143 net143 o_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput154 net154 o_mem_long vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4720__A1 core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8134_ core_0.execute.rf.reg_outputs\[1\]\[15\] _3758_ _3771_ _3778_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput165 net165 o_req_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5346_ _1435_ _1463_ _0015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput176 net176 o_req_ppl_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_195_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput187 net187 sr_bus_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_227_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_2721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput198 net198 sr_bus_data_o[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8462__A2 _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8065_ _3401_ _3737_ _3739_ _0459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5277_ core_0.execute.hold_valid core_0.decode.o_submit _0923_ _1398_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_215_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6473__A1 core_0.dec_sys vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7016_ _2795_ _2936_ _2944_ _2945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_215_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input28_I i_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_133_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_106_Right_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6225__A1 _2165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8967_ _4451_ _0649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7973__A1 core_0.execute.rf.reg_outputs\[5\]\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7918_ core_0.execute.rf.reg_outputs\[6\]\[2\] _3652_ _3648_ _3655_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8898_ _1431_ _4411_ _0620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_194_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_1756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_2850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7849_ core_0.execute.rf.reg_outputs\[8\]\[5\] _3613_ _3609_ _3615_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6528__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8005__B _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwire215 _0880_ net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_136_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9519_ _0529_ clknet_leaf_118_i_clk core_0.execute.alu_mul_div.div_res\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7844__B _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_2108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_58_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output96_I net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8150__A1 _3427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6700__A2 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_226_3227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8453__A2 _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A1 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5267__A2 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8205__A2 _3830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7964__A1 _3434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4778__A1 _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_237_3356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7716__A1 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6519__A2 _1925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 i_core_int_sreg[5] net12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput23 i_mem_data[11] net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_155_2377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput34 i_mem_data[7] net34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8569__C _4046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput45 i_req_data[17] net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput56 i_req_data[27] net56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput67 i_req_data[8] net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8141__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_208_Right_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5200_ core_0.fetch.prev_req_branch_pred _1343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6180_ _2166_ _2167_ _2168_ _2169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5131_ _1250_ _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8444__A2 _4031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6455__A1 _1163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _1226_ _1086_ _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_236_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6207__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8821_ core_0.execute.pc_high_out\[2\] _4327_ _4347_ _4348_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7929__B _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7955__A1 core_0.execute.rf.reg_outputs\[5\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4769__A1 core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8752_ core_0.execute.sreg_scratch.o_d\[3\] _4295_ _4299_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5964_ _1950_ _1951_ _1952_ _1953_ _1954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_48_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7703_ core_0.execute.rf.reg_outputs\[12\]\[7\] _3526_ _3528_ _3531_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4915_ core_0.fetch.prev_request_pc\[10\] _1037_ _1049_ core_0.fetch.prev_request_pc\[9\]
+ _1095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8683_ _4203_ _4100_ _4246_ _1661_ _4247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5895_ core_0.decode.oc_alu_mode\[9\] _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_75_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7634_ _3457_ _3477_ _3490_ _0277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4846_ core_0.fetch.out_buffer_data_instr\[23\] _1027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_191_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8380__A1 _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__B _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ core_0.execute.rf.reg_outputs\[15\]\[6\] _3429_ _3422_ _3442_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4777_ core_0.dec_l_reg_sel\[0\] _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XANTENNA__6930__A2 _2733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9304_ _0314_ clknet_leaf_154_i_clk core_0.execute.rf.reg_outputs\[12\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6516_ _2456_ _2457_ _2458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_rebuffer20_I net247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7496_ _3381_ _3382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_210_3028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8132__A1 core_0.execute.rf.reg_outputs\[1\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_190_2791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5184__B _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9235_ _0246_ clknet_leaf_143_i_clk core_0.ew_reg_ie\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_70_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6447_ _1185_ _2386_ _2406_ _0174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6694__A1 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5497__A2 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9166_ _0177_ clknet_leaf_82_i_clk core_0.execute.mem_stage_pc\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6378_ _1544_ _2346_ _2351_ _2352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_246_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8117_ core_0.execute.rf.reg_outputs\[1\]\[7\] _3765_ _3756_ _3769_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5329_ _1239_ _1247_ _1259_ _1446_ _1447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8435__A2 _4033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9097_ _0122_ clknet_leaf_83_i_clk core_0.fetch.pc_flush_override vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_54_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8048_ core_0.execute.rf.reg_outputs\[3\]\[10\] _3722_ _3718_ _3729_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_215_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6997__A2 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_221_3168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8738__A3 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7946__A1 core_0.execute.rf.reg_outputs\[6\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6749__A2 net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8371__A1 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5185__A1 _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4932__A1 core_0.fetch.prev_request_pc\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8123__A1 _3453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_232_3297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4489__I core_0.execute.rf.reg_outputs\[4\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5488__A2 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_232_Left_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_219_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8426__A2 _1680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6988__A2 _2901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7749__B _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7937__A1 _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9486__CLK clknet_leaf_21_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_241_Left_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_33_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4700_ core_0.execute.rf.reg_outputs\[14\]\[0\] net262 net321 core_0.execute.rf.reg_outputs\[12\]\[0\]
+ _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_84_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5680_ _1684_ _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_151_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8362__A1 _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ core_0.execute.rf.reg_outputs\[12\]\[6\] _0699_ net286 core_0.execute.rf.reg_outputs\[13\]\[6\]
+ _0820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5176__A1 _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7350_ _2699_ _3270_ _3271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4562_ core_0.execute.rf.reg_outputs\[4\]\[11\] _0719_ _0709_ core_0.execute.rf.reg_outputs\[8\]\[11\]
+ _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8114__A1 _3434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6301_ _2185_ _2220_ _2283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7281_ _2711_ _3192_ _3203_ _3204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8665__A2 _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4493_ _0674_ _0681_ _0690_ _0691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_92_1619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6676__A1 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9020_ _0047_ clknet_leaf_78_i_clk core_0.fetch.out_buffer_data_instr\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6232_ _2141_ _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_168_2524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4687__B1 net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6163_ core_0.execute.alu_mul_div.div_cur\[12\] _1831_ _2152_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_209_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5114_ _1268_ _1245_ _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XPHY_EDGE_ROW_191_Right_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_176_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6094_ core_0.execute.rf.reg_outputs\[1\]\[3\] _0954_ _0955_ _0962_ _2084_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5045_ _1031_ _1146_ _1164_ _1214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_240_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8762__C _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6563__B _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7928__A1 _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8804_ core_0.execute.pc_high_out\[0\] _4327_ _4332_ _4333_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clone40_I _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6996_ _2672_ _2925_ _2926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_149_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_rebuffer68_I _1835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_2664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8735_ _1397_ _1415_ _1418_ net105 _1253_ _4288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_34_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5947_ core_0.execute.rf.reg_outputs\[2\]\[10\] _1797_ _1781_ core_0.execute.rf.reg_outputs\[10\]\[10\]
+ _1937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_177_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8666_ net82 _1699_ _1711_ _4205_ _4233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_192_2820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7156__A2 _3081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5878_ net177 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
Xclkbuf_4_7__f_i_clk clknet_3_3_0_i_clk clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7617_ core_0.execute.rf.reg_outputs\[14\]\[3\] _3477_ _3467_ _3481_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4829_ _0894_ _1009_ _1010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8597_ _4167_ _4172_ _4173_ _0557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5693__I _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__A2 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7548_ _3382_ core_0.ew_data\[4\] _3426_ _3427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__8105__A1 _3408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6116__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7479_ core_0.dec_rf_ie\[8\] core_0.ew_reg_ie\[8\] _3366_ _3373_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8656__A2 _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6667__A1 _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9218_ _0229_ clknet_leaf_80_i_clk net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4678__B1 net347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8408__A2 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9149_ _0161_ clknet_leaf_106_i_clk core_0.execute.hold_valid vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_228_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A1 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clone6_B _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8672__C _4219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__A2 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7919__A1 _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_205_2974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4772__I core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8592__A1 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4602__B1 _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_234_3315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_3326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7147__A2 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8344__A1 core_0.execute.alu_mul_div.mul_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5158__A1 _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8895__A2 _4383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_2336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6107__B1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5108__I _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6658__A1 _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4669__B1 net284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_3455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7458__I0 net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7083__A1 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_2465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5633__A2 _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6830__A1 _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8958__I0 net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _2773_ _2782_ _2783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_18_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5801_ _0957_ _0958_ _1790_ _1791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_159_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6781_ _1874_ _2371_ _2714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_8_Right_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8520_ _4047_ _4105_ _4106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5732_ _1714_ _1725_ _0140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_174_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8335__A1 _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8451_ _4041_ _4042_ _4043_ _4044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5663_ _1667_ _1670_ _1671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6897__A1 _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7402_ _1880_ _2556_ _3315_ _3320_ _3321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_5_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4614_ core_0.execute.rf.reg_outputs\[4\]\[7\] _0719_ net316 core_0.execute.rf.reg_outputs\[8\]\[7\]
+ _0804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8382_ core_0.execute.alu_mul_div.mul_res\[13\] _3986_ _3994_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5594_ _1368_ _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_53_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7333_ _3248_ _3253_ _1292_ _3254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7942__B _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4545_ _0730_ _0716_ _0735_ _0740_ _0741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_170_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7264_ _3186_ _3175_ _3187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_96_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ core_0.execute.rf.reg_outputs\[6\]\[15\] _0670_ _0673_ core_0.execute.rf.reg_outputs\[2\]\[15\]
+ _0674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9003_ _0030_ clknet_leaf_15_i_clk core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_96_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6215_ core_0.execute.alu_mul_div.div_cur\[14\] _2143_ _2149_ _2203_ _2204_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_96_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Right_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7195_ core_0.execute.alu_mul_div.div_cur\[9\] _2128_ _3117_ _3119_ _3120_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_244_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6146_ _1433_ _1735_ _2136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_51_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7074__A1 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8265__S _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6077_ _2063_ _2064_ _2065_ _2066_ _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5624__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6821__A1 _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _1199_ _1029_ _1158_ _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input10_I i_core_int_sreg[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5688__I _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__B _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8574__A1 net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7377__A2 _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6979_ _1751_ _2002_ _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XPHY_EDGE_ROW_48_Right_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8718_ _4212_ core_0.execute.mem_stage_pc\[14\] _4202_ _4275_ _4276_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7129__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8649_ core_0.dec_wfi _4219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__8877__A2 _4385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8013__B _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6888__A1 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5560__A1 core_0.fetch.prev_request_pc\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__B2 net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8667__C _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_57_Right_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7301__A2 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5312__A1 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_207_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7065__A1 _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A2 _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4716__B core_0.execute.irq_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_240_3396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_230_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_66_Right_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_230_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8317__A1 core_0.execute.alu_mul_div.mul_res\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8868__A2 _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6879__A1 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7540__A2 core_0.ew_data\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7762__B _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5551__A1 core_0.fetch.prev_request_pc\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5551__B2 net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_75_Right_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__A1 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6000_ core_0.execute.rf.reg_outputs\[13\]\[12\] _1792_ _1815_ core_0.execute.rf.reg_outputs\[9\]\[12\]
+ _1990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_226_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input2_I i_core_int_sreg[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7056__A1 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8253__B1 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__A2 _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6803__A1 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7951_ core_0.execute.rf.reg_outputs\[5\]\[0\] _3673_ _3663_ _3674_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Right_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_222_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6902_ _2699_ _2832_ _2833_ _2834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7882_ _3421_ _3628_ _3633_ _0382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8556__A1 _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8556__B2 _2134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9621_ _0631_ clknet_leaf_133_i_clk core_0.dec_used_operands\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6833_ core_0.execute.alu_mul_div.div_cur\[1\] _0997_ _2765_ _2766_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_176_2623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9552_ _0562_ clknet_leaf_67_i_clk core_0.execute.sreg_irq_pc.o_d\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _1402_ _2697_ _2135_ _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8308__A1 _3081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8503_ _4088_ _4090_ _4051_ _0546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_175_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5715_ _1249_ _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_134_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9483_ _0493_ clknet_leaf_15_i_clk net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__5790__A1 _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4593__A2 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _2621_ _2631_ _2634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_174_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8434_ _4018_ _4031_ _4033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5646_ core_0.decode.i_flush core_0.fetch.dbg_out core_0.fetch.flush_event_invalidate
+ _1659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_93_Right_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5542__A1 _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8365_ _3966_ _3863_ _3978_ _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5577_ _1235_ core_0.fetch.submitable _1619_ _0091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7316_ _2672_ net196 _3237_ _3238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_229_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4896__A3 _1071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4528_ core_0.execute.rf.reg_outputs\[3\]\[14\] net341 _0700_ core_0.execute.rf.reg_outputs\[12\]\[14\]
+ _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8296_ _1536_ _1680_ _3914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input58_I i_req_data[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7295__A1 _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8492__B1 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7247_ core_0.execute.alu_mul_div.div_res\[11\] _3170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__8492__C2 _4080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_2752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_244_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7178_ _2571_ _3102_ _3103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7047__A1 _2438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6129_ _2011_ _1898_ _2118_ _2119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8795__A1 core_0.dec_sreg_store vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7598__A2 _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A2 _0998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_2933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8547__A1 _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8547__B2 _2134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7847__B _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_107_1798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_218_3129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A2 _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_198_2892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_120_1954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7770__A2 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4584__A2 _0666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_136_2139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_128_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7522__A2 _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7286__A1 _2480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__A2 _1818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4497__I net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_229_3258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5836__A2 _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_242_3414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7038__A1 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5300__A4 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7601__I _3469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_2279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8786__A1 _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7589__A2 _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_2435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_182_Left_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_86_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8538__A1 _1185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7757__B _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7210__A1 _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5772__A1 _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4575__A2 _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5500_ net46 _1554_ _1577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ _2421_ _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_82_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8710__A1 _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7513__A2 _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_2564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5431_ _1519_ _1486_ _1527_ _1501_ _0036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_191_Left_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_1680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8150_ _3427_ _3780_ _3788_ _0495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5362_ _1464_ _1475_ _0019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7101_ _1899_ net214 _3028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8081_ _3446_ _3737_ _3748_ _0466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5293_ core_0.dec_jump_cond_code\[4\] _1413_ _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_227_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_0_i_clk clknet_4_0__leaf_i_clk clknet_leaf_0_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7032_ _1683_ core_0.execute.sreg_irq_pc.o_d\[5\] _2960_ _2961_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8226__B1 _3830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8777__A1 core_0.execute.sreg_scratch.o_d\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_2693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8983_ _1497_ _4459_ _0657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5031__I net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7934_ core_0.execute.rf.reg_outputs\[6\]\[9\] _3657_ _3663_ _3664_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8529__A1 net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7865_ _3463_ _3607_ _3623_ _0375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_194_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7201__A1 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6004__A2 _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9604_ _0614_ clknet_leaf_50_i_clk core_0.execute.pc_high_buff_out\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6816_ _2748_ _2447_ _2749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_203_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7796_ _3473_ _3564_ _3583_ _0346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_46_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7752__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9535_ _0545_ clknet_leaf_76_i_clk net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_175_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5763__A1 _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6747_ core_0.execute.sreg_irq_flags.o_d\[0\] _1686_ net227 _2680_ _2681_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_190_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6960__B1 _2768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9466_ _0476_ clknet_leaf_50_i_clk core_0.execute.rf.reg_outputs\[1\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_33_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6678_ core_0.execute.rf.reg_outputs\[7\]\[1\] _2611_ _2612_ core_0.execute.rf.reg_outputs\[5\]\[1\]
+ _2619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8701__A1 _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5629_ _1046_ _1628_ _1650_ _0112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8417_ _1667_ _1675_ _4022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9397_ _0407_ clknet_leaf_148_i_clk core_0.execute.rf.reg_outputs\[6\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4869__A3 _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8348_ _3960_ _3962_ _3963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_14_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output164_I net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8279_ core_0.execute.alu_mul_div.mul_res\[6\] _3898_ _3863_ _3899_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5818__A2 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6491__A2 _2039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8768__A1 core_0.execute.sreg_scratch.o_d\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_54_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6243__A2 _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7991__A2 _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7577__B _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_wire213_I _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer90 _1798_ net337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_185_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8940__A1 core_0.decode.i_imm_pass\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7743__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5754__A1 _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7259__A1 _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8456__B1 _2766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_236_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_208_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8471__A3 _4062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6482__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5285__A3 net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8759__A1 core_0.execute.sreg_scratch.o_d\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4891__S _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ _1968_ _1969_ _1970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7982__A2 _3671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4931_ _1109_ _1031_ _1110_ _1111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7650_ _1430_ _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__8231__I0 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4862_ _0892_ net45 _1042_ _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_28_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7195__B1 _3117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7734__A2 _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6601_ net266 _2366_ _2543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_170_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_15 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4548__A2 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7581_ core_0.execute.rf.reg_outputs\[15\]\[9\] _3429_ _3422_ _3455_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4793_ core_0.ew_reg_ie\[7\] _0966_ _0942_ _0974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6942__B1 _2870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9320_ _0330_ clknet_leaf_148_i_clk core_0.execute.rf.reg_outputs\[11\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6532_ net242 _2371_ _2470_ _2474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7498__A1 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9251_ _0261_ clknet_leaf_7_i_clk core_0.execute.rf.reg_outputs\[15\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6463_ _2413_ _0902_ _0183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9242__CLK clknet_leaf_2_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8111__B _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5227__S _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8202_ _1000_ _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_30_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5414_ core_0.decode.i_instr_l\[14\] _1509_ _1510_ core_0.decode.i_instr_l\[10\]
+ _1495_ _1514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_140_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput100 net100 dbg_r0[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9182_ _0193_ clknet_leaf_46_i_clk net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4705__C1 core_0.execute.rf.reg_outputs\[1\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput111 net111 o_instr_long_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_179_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6394_ _2354_ _2366_ _2367_ _2368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput122 net122 o_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput133 net133 o_mem_addr_high[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8133_ _3469_ _3760_ _3777_ _0489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput144 net144 o_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5345_ core_0.dec_rf_ie\[5\] _1438_ _1441_ _1462_ _1463_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_140_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput155 net155 o_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4720__A2 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput166 net166 o_req_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput177 net177 sr_bus_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_227_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput188 net188 sr_bus_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_clkbuf_4_5__f_i_clk_I clknet_3_2_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_2722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8064_ core_0.execute.rf.reg_outputs\[2\]\[0\] _3738_ _3730_ _3739_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput199 net231 sr_bus_data_o[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ _1396_ _1397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_49_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7015_ core_0.decode.oc_alu_mode\[6\] _2453_ _2938_ _2940_ _2943_ _2944_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6473__A2 _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__A1 net293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7422__A1 _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8966_ net183 core_0.decode.i_imm_pass\[15\] _1263_ _4451_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_39_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7973__A2 _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7917_ _3409_ _3651_ _3654_ _0396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4814__B _0994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5696__I _1700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8897_ core_0.execute.pc_high_buff_out\[7\] _4386_ _4410_ _4411_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_104_1757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7848_ _3428_ _3606_ _3614_ _0367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_195_2851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7725__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5736__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7779_ _3447_ _3563_ _3574_ _0338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_191_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9518_ _0528_ clknet_leaf_117_i_clk core_0.execute.alu_mul_div.div_res\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xwire227 _1408_ net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_163_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_101_i_clk clknet_4_13__leaf_i_clk clknet_leaf_101_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_163_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9449_ _0459_ clknet_leaf_136_i_clk core_0.execute.rf.reg_outputs\[2\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8021__B _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8150__A2 _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output89_I net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_116_i_clk clknet_4_7__leaf_i_clk clknet_leaf_116_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_115_1897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_226_3228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5380__B _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A2 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7661__A1 _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_2238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8691__B _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7964__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A2 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_237_3357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7716__A2 _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8913__A1 _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5727__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4935__C1 core_0.fetch.prev_request_pc\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 i_core_int_sreg[6] net13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_155_2367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput24 i_mem_data[12] net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_2378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput35 i_mem_data[8] net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput46 i_req_data[18] net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput57 i_req_data[28] net57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4950__A2 _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput68 i_req_data[9] net68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8141__A2 _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6230__I _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_172_Right_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6152__A1 _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_228_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5130_ core_0.decode.oc_alu_mode\[7\] _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_58_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6455__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7652__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_80_i_clk clknet_4_14__leaf_i_clk clknet_leaf_80_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5061_ net71 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7404__A1 _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6207__A2 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8820_ net216 _4328_ _4326_ _4346_ _4347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_0_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7955__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_95_i_clk clknet_4_13__leaf_i_clk clknet_leaf_95_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_36_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5963_ core_0.execute.rf.reg_outputs\[2\]\[11\] _1797_ _1781_ core_0.execute.rf.reg_outputs\[10\]\[11\]
+ _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4769__A2 core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8751_ net216 _4294_ _4298_ _4287_ _0586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8106__B _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4914_ _1092_ _1093_ _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7702_ _3441_ _3520_ _3530_ _0305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_220_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8682_ net85 _1699_ _1717_ _4205_ _4246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5894_ _1755_ net344 _1812_ _1884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_74_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8904__A1 _1257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7707__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _1017_ net58 _1025_ _1026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_35_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7633_ core_0.execute.rf.reg_outputs\[14\]\[10\] _3482_ _3486_ _3490_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5718__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7564_ _3440_ _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_172_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4776_ core_0.dec_l_reg_sel\[1\] _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_117_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9303_ _0313_ clknet_leaf_153_i_clk core_0.execute.rf.reg_outputs\[12\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6515_ _1846_ net213 _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_71_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7495_ core_0.ew_mem_access _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_160_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_210_3029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_2792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8132__A2 _3758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_33_i_clk clknet_4_8__leaf_i_clk clknet_leaf_33_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6446_ core_0.execute.mem_stage_pc\[10\] _2395_ _2404_ _2406_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9234_ _0245_ clknet_leaf_140_i_clk core_0.ew_reg_ie\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_rebuffer13_I net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7680__B _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6694__A2 _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9165_ _0176_ clknet_leaf_81_i_clk core_0.execute.mem_stage_pc\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7891__A1 core_0.execute.rf.reg_outputs\[7\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6377_ _1542_ net218 _2350_ core_0.execute.alu_mul_div.cbit\[1\] _2351_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7172__S _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8116_ _3440_ _3759_ _3768_ _0481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5328_ _1233_ _1313_ _1289_ _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9096_ _0121_ clknet_leaf_103_i_clk core_0.fetch.flush_event_invalidate vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input40_I i_req_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_i_clk clknet_4_10__leaf_i_clk clknet_leaf_48_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8047_ _3453_ _3715_ _3728_ _0452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6446__A2 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7643__A1 core_0.execute.rf.reg_outputs\[14\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5259_ core_0.execute.alu_flag_reg.o_d\[2\] _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_215_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_221_3169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8949_ _4442_ _0640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5709__A1 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7855__B _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__A1 _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5185__A2 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__A2 _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8123__A2 _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_232_3298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__I _2039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7882__A1 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4696__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_237_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6437__A2 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7634__A1 _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7485__I1 core_0.ew_reg_ie\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7937__A2 _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_11__f_i_clk_I clknet_3_5_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__A1 core_0.execute.rf.reg_outputs\[15\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_241_Right_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_146_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4630_ core_0.execute.rf.reg_outputs\[6\]\[6\] net223 net312 core_0.execute.rf.reg_outputs\[2\]\[6\]
+ _0819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_170_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ core_0.execute.rf.reg_outputs\[5\]\[11\] _0676_ _0679_ core_0.execute.rf.reg_outputs\[11\]\[11\]
+ _0755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8114__A2 _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _1547_ _2275_ _2281_ _2282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7280_ _2710_ _3201_ _3202_ _3203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6125__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4492_ core_0.execute.rf.reg_outputs\[7\]\[15\] net296 _0686_ core_0.execute.rf.reg_outputs\[14\]\[15\]
+ _0689_ _0690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_123_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8596__B _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6231_ _2215_ _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_110_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6676__A2 _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4687__A1 core_0.execute.rf.reg_outputs\[9\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_2525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ core_0.execute.alu_mul_div.div_cur\[12\] _1831_ _2151_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_176_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5113_ core_0.decode.i_instr_l\[5\] _1268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6428__A2 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7625__A1 _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6093_ core_0.execute.rf.reg_outputs\[2\]\[3\] net335 net317 core_0.execute.rf.reg_outputs\[6\]\[3\]
+ _2083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5044_ _1158_ _1212_ _1213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_109_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9430__CLK clknet_leaf_144_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5239__I0 core_0.ew_data\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7928__A2 _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8803_ _0890_ _4328_ _4327_ _4331_ _4332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_177_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5939__A1 net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6995_ _2897_ _2899_ _2924_ _2925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6061__B1 _1787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8734_ _4218_ _4283_ _4286_ _4287_ _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_179_2665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5946_ core_0.execute.rf.reg_outputs\[5\]\[10\] _1785_ _1802_ core_0.execute.rf.reg_outputs\[14\]\[10\]
+ _1936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_149_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9580__CLK clknet_leaf_21_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8665_ core_0.execute.sreg_irq_pc.o_d\[5\] _4210_ _4232_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5877_ _1768_ _1866_ _1867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_2821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8353__A2 _3947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4828_ core_0.fetch.out_buffer_data_instr\[0\] _1009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7616_ _3415_ _3476_ _3480_ _0269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8596_ core_0.execute.alu_flag_reg.o_d\[1\] _4167_ _3797_ _4173_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7547_ _3381_ _3424_ _3425_ _3426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4759_ _0936_ _0937_ _0938_ _0939_ _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_90_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8105__A2 _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6116__A1 core_0.execute.rf.reg_outputs\[1\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7478_ _3372_ _0239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9217_ _0228_ clknet_leaf_79_i_clk net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6667__A2 _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6429_ _1433_ _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_101_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4678__A1 core_0.execute.rf.reg_outputs\[5\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9148_ _0160_ clknet_leaf_117_i_clk core_0.execute.alu_mul_div.div_cur\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__8408__A3 _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7467__I1 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7616__A1 _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6419__A2 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9079_ _0104_ clknet_leaf_101_i_clk core_0.decode.i_imm_pass\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_215_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_215_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7919__A2 _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8041__A1 _3440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_205_2975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4602__A1 core_0.execute.rf.reg_outputs\[7\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4602__B2 core_0.execute.rf.reg_outputs\[3\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7585__B _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_234_3316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__A2 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_2337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6107__B2 core_0.execute.rf.reg_outputs\[9\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4669__B2 core_0.execute.rf.reg_outputs\[13\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_245_3456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7607__A1 _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7458__I1 _3297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_163_2466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6830__A2 core_0.execute.alu_mul_div.mul_res\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5060__S _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8032__A1 _3414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Left_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_159_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__B1 _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8583__A2 _2761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5800_ core_0.dec_l_reg_sel\[3\] core_0.dec_l_reg_sel\[2\] _1790_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6780_ core_0.execute.alu_mul_div.i_mul _2713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_186_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5731_ net196 _1697_ _1700_ core_0.execute.sreg_priv_control.o_d\[12\] _1725_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8450_ net78 _4041_ _4043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5662_ _1668_ _1669_ _1670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_29_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5149__A2 _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7401_ _3073_ _3319_ _3320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4613_ core_0.execute.rf.reg_outputs\[5\]\[7\] net222 _0679_ core_0.execute.rf.reg_outputs\[11\]\[7\]
+ _0803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6897__A2 _1411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8381_ core_0.execute.alu_mul_div.mul_res\[14\] _2375_ _3993_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_2595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5593_ _1627_ _0099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7332_ _2468_ _2472_ _2470_ _3253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4544_ _0736_ _0737_ _0738_ _0739_ _0740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XPHY_EDGE_ROW_68_Left_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7263_ _2859_ _3069_ _3182_ _1768_ _3185_ _3186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_229_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4475_ _0672_ _0673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5235__S _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7514__I _3396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9002_ _0029_ clknet_leaf_135_i_clk core_0.dec_r_reg_sel\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6214_ _2148_ _2152_ _2202_ _2203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_209_3020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7194_ _3118_ _1314_ core_0.execute.alu_mul_div.i_mod _3119_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_110_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6145_ _1402_ core_0.execute.sreg_irq_pc.o_d\[0\] _2135_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_51_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6076_ core_0.execute.rf.reg_outputs\[6\]\[6\] net219 _1787_ core_0.execute.rf.reg_outputs\[3\]\[6\]
+ _2066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_127_2041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5027_ _1150_ _1198_ _1199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_212_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_77_Left_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer80_I _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4832__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__C _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8574__A2 _4052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6978_ _2495_ _2906_ _2907_ core_0.decode.oc_alu_mode\[11\] _2908_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_49_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8717_ _4224_ _4141_ _4274_ _1662_ _4275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_0_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5929_ core_0.execute.rf.reg_outputs\[14\]\[8\] _1801_ net339 core_0.execute.rf.reg_outputs\[11\]\[8\]
+ _1919_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_165_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6337__A1 _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8648_ net201 _0900_ _4218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output194_I net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6888__A2 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_86_Left_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8579_ _3150_ _4156_ _4157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5560__A2 _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5312__A2 _1428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output71_I net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4520__B1 _0673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8683__C _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7065__A2 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_95_Left_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_215_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_124_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8014__A1 _3459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_3397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_196_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6576__A1 _2439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4587__B1 _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6879__A2 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5000__A1 core_0.fetch.prev_request_pc\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5551__A2 _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_49_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7828__A1 core_0.execute.rf.reg_outputs\[9\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6500__A1 _2074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5303__A2 net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_207_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8253__B2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5789__I _1778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6803__A2 _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7950_ _3671_ _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_89_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_206_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__A1 core_0.ew_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6901_ _2700_ _2785_ _2831_ _2833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_49_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7881_ core_0.execute.rf.reg_outputs\[7\]\[3\] _3629_ _3621_ _3633_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_194_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8556__A2 core_0.execute.sreg_irq_pc.o_d\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9620_ _0630_ clknet_leaf_133_i_clk core_0.dec_used_operands\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6832_ _2128_ _2764_ _2765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_15_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6567__A1 _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_176_2624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4578__B1 _0707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9551_ _0561_ clknet_leaf_58_i_clk core_0.execute.irq_en vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6763_ _2679_ _2686_ _2696_ _1226_ _2694_ _2697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_175_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8308__A2 _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8502_ _4047_ _4089_ _4090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5714_ _1608_ _1713_ _0134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6694_ _2422_ _2632_ _2633_ _0193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9482_ _0492_ clknet_leaf_22_i_clk net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__5790__A2 core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7953__B _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8433_ _3118_ _4032_ _2258_ _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5645_ _1249_ _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_131_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_215_3090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _1072_ core_0.fetch.submitable _1619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8364_ _3863_ _3977_ _3978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7315_ _3226_ _3236_ core_0.dec_mem_access _3237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4527_ core_0.execute.rf.reg_outputs\[1\]\[14\] net302 _0695_ core_0.execute.rf.reg_outputs\[10\]\[14\]
+ _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7819__A1 _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7244__I _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8295_ _3913_ _0515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_229_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8492__A1 _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7246_ _2839_ _3167_ _3169_ _0210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8492__B2 _2134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_2753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7177_ _1863_ _3101_ _3102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
X_6128_ _2076_ _2104_ _2117_ _2118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5058__A1 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8795__A2 _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8075__I _3647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6059_ core_0.execute.rf.reg_outputs\[14\]\[7\] _1801_ net339 core_0.execute.rf.reg_outputs\[11\]\[7\]
+ _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4805__A1 core_0.ew_reg_ie\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4805__B2 core_0.ew_reg_ie\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_202_2934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__B1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output207_I net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_198_2893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8678__C _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_50_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8483__A1 _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_229_3259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8694__B _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5297__A1 _1417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_242_3415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5049__A1 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_216_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_2436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6661__C _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_200_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5221__A1 core_0.ew_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8869__B _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5430_ _1495_ _1522_ _1523_ _1526_ _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_171_2565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6721__A1 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5361_ core_0.dec_rf_ie\[9\] _1438_ _1472_ _1474_ _1475_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_97_1681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7100_ _3022_ _3026_ _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8474__A1 _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8080_ core_0.execute.rf.reg_outputs\[2\]\[7\] _3743_ _3745_ _3748_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5292_ _1403_ _1412_ _1413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_77_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5288__A1 net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7031_ _1401_ _2959_ _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_227_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8226__A1 _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__B2 core_0.execute.alu_mul_div.mul_res\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8982_ core_0.dec_rf_ie\[2\] _1482_ _1462_ _1476_ _4459_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6788__A1 _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_2694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7933_ _3647_ _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__8529__A2 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7864_ core_0.execute.rf.reg_outputs\[8\]\[12\] _3613_ _3621_ _3623_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9603_ _0613_ clknet_leaf_50_i_clk core_0.execute.pc_high_buff_out\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _1896_ _2341_ _2748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_147_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7795_ core_0.execute.rf.reg_outputs\[10\]\[15\] _3562_ _3580_ _3583_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_46_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_186_Right_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9534_ _0544_ clknet_leaf_69_i_clk net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_46_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6746_ net184 _1868_ _1409_ _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_147_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5763__A2 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer43_I _0666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9465_ _0475_ clknet_leaf_61_i_clk core_0.execute.rf.reg_outputs\[1\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_162_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6677_ core_0.execute.rf.reg_outputs\[1\]\[1\] _2608_ _2609_ core_0.execute.rf.reg_outputs\[3\]\[1\]
+ _2618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_33_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8416_ _2230_ _4021_ _0528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5515__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6712__A1 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_4_0_i_clk clknet_0_i_clk clknet_3_4_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5628_ core_0.decode.i_imm_pass\[8\] _1645_ _1650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input70_I i_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9396_ _0406_ clknet_leaf_3_i_clk core_0.execute.rf.reg_outputs\[6\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4598__I _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8347_ _3945_ _3947_ _3961_ _3962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ _1608_ _1609_ _0083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8465__A1 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7268__A2 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8278_ net214 _3827_ _3897_ _3898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5279__A1 _0995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output157_I net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5818__A3 _1790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7229_ core_0.execute.alu_mul_div.div_res\[10\] _3153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_218_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8019__B _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8768__A2 _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5451__A1 _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer80 _0692_ net308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_95_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer91 _1803_ net338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_139_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8940__A2 _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_153_Right_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5754__A2 net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7593__B _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5892__I _1757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8456__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8456__B2 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8208__A1 _3828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5690__A1 _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8759__A2 _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7431__A2 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ core_0.fetch.prev_request_pc\[3\] _1060_ _1110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_188_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Left_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5993__A2 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8231__I1 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4861_ core_0.fetch.out_buffer_valid _1041_ _1042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7195__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6600_ _2539_ _2541_ _2542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_7_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_16 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7580_ _3453_ _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_172_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4792_ core_0.ew_reg_ie\[13\] _0963_ _0964_ core_0.ew_reg_ie\[14\] _0966_ core_0.ew_reg_ie\[15\]
+ _0973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XPHY_EDGE_ROW_120_Right_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5745__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6942__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6531_ net241 _2371_ _2473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_28_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7498__A2 _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8695__A1 _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9250_ _0260_ clknet_leaf_9_i_clk core_0.execute.rf.reg_outputs\[15\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6462_ _2413_ _0904_ _0182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_212_3060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8201_ _3802_ _1883_ _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__4705__B1 net318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5413_ _0947_ _1486_ _1513_ _1501_ _0032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput101 net101 dbg_r0[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_9181_ _0192_ clknet_leaf_44_i_clk net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_41_Left_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6393_ _2354_ _1999_ _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4705__C2 net302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput112 net112 o_instr_long_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput123 net123 o_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput134 net134 o_mem_addr_high[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8447__A1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8132_ core_0.execute.rf.reg_outputs\[1\]\[14\] _3758_ _3771_ _3777_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5344_ core_0.decode.i_instr_l\[10\] _1437_ _1461_ _1462_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xoutput145 net145 o_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_112_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput156 net156 o_mem_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_195_11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput167 net167 o_req_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5751__B _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput178 net178 sr_bus_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput189 net189 sr_bus_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_195_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8063_ _3736_ _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5275_ core_0.execute.sreg_jtr_buff.o_d\[0\] _0900_ _1396_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_195_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_2723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7014_ _1851_ _2941_ _2942_ _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7670__A2 _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__A2 _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6138__I core_0.execute.alu_mul_div.i_mod vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5042__I net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7678__B _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_50_Left_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8965_ _4450_ _0648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5433__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7916_ core_0.execute.rf.reg_outputs\[6\]\[1\] _3652_ _3648_ _3654_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_214_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8896_ net277 _4387_ _4385_ _4409_ _4410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_38_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_210_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7847_ core_0.execute.rf.reg_outputs\[8\]\[4\] _3613_ _3609_ _3614_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_195_2852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8922__A2 _1322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7778_ core_0.execute.rf.reg_outputs\[10\]\[7\] _3570_ _3568_ _3574_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6933__A1 _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9517_ _0527_ clknet_leaf_118_i_clk core_0.execute.alu_mul_div.div_res\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9067__CLK clknet_leaf_110_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ _2422_ _2663_ _2664_ _0197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_190_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9448_ _0458_ clknet_leaf_146_i_clk core_0.execute.rf.reg_outputs\[3\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_59_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9379_ _0389_ clknet_leaf_7_i_clk core_0.execute.rf.reg_outputs\[7\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_1887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_226_3229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7110__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7661__A2 _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_222_Right_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7413__A2 _3330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5424__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7177__A1 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_237_3358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8913__A2 _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5188__B1 _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6924__A1 _2795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6924__B2 _2480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4935__B1 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4935__C2 _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8212__B core_0.execute.alu_mul_div.cbit\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 i_core_int_sreg[7] net14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_155_2368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput25 i_mem_data[13] net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput36 i_mem_data[9] net36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8677__A1 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput47 i_req_data[19] net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput58 i_req_data[29] net58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput69 i_req_data_valid net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_150_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6152__A2 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4966__I _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7101__A1 _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ core_0.fetch.prev_request_pc\[0\] _1054_ _1158_ _1225_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_236_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7652__A2 _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_224_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5415__A1 _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8750_ core_0.execute.sreg_scratch.o_d\[2\] _4295_ _4298_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ core_0.execute.rf.reg_outputs\[5\]\[11\] _1785_ _1802_ core_0.execute.rf.reg_outputs\[14\]\[11\]
+ _1952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5966__A2 _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7701_ core_0.execute.rf.reg_outputs\[12\]\[6\] _3526_ _3528_ _3530_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4913_ core_0.fetch.prev_request_pc\[10\] _1037_ _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7168__A1 _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8681_ core_0.execute.sreg_irq_pc.o_d\[8\] _4209_ _4245_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5893_ _1882_ _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_75_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8904__A2 _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7632_ _3454_ _3476_ _3489_ _0276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4844_ _0892_ _1024_ _1025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7563_ _3382_ core_0.ew_data\[6\] _3439_ _3440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_43_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ _0954_ _0955_ _0956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8122__B _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9302_ _0312_ clknet_leaf_153_i_clk core_0.execute.rf.reg_outputs\[12\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8668__A1 _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6514_ net319 _1925_ _2456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_132_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7494_ _3380_ _0247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7961__B _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_190_2793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9233_ _0244_ clknet_leaf_140_i_clk core_0.ew_reg_ie\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_141_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6445_ _2403_ _2385_ _2405_ _0173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_141_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7340__A1 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8776__C _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_97_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9164_ _0175_ clknet_leaf_92_i_clk core_0.execute.mem_stage_pc\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7891__A2 _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6376_ _1541_ _2349_ _2350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8115_ core_0.execute.rf.reg_outputs\[1\]\[6\] _3765_ _3756_ _3768_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5327_ _1239_ _1443_ _1444_ _1445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_9095_ _0120_ clknet_leaf_81_i_clk core_0.fetch.dbg_out vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6296__C _2229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8046_ core_0.execute.rf.reg_outputs\[3\]\[9\] _3722_ _3718_ _3728_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7643__A2 _3475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5258_ _1373_ _1375_ _1377_ _1378_ _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_input33_I i_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ _1334_ _0003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_221_3159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8948_ net189 core_0.decode.i_imm_pass\[6\] _1264_ _4442_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_211_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7159__A1 _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8879_ _0902_ _4383_ _4397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6382__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8659__A1 _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_232_3299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7331__A1 _2939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7882__A2 _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4696__A2 _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8831__A1 core_0.execute.pc_high_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7634__A2 _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_202_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6070__A1 core_0.execute.rf.reg_outputs\[5\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_215_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__A2 _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_106_Left_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8898__A1 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6241__I _2229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4560_ core_0.execute.rf.reg_outputs\[10\]\[11\] _0694_ _0704_ core_0.execute.rf.reg_outputs\[9\]\[11\]
+ _0754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_119_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8877__B _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4491_ _0687_ net299 net275 net293 _0689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__6125__A2 _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6230_ _2218_ _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_228_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_168_2526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4687__A2 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_115_Left_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6161_ _2148_ _2149_ _2150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5112_ _1266_ _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__8822__A1 _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6092_ core_0.execute.rf.reg_outputs\[15\]\[3\] _0944_ _1784_ core_0.execute.rf.reg_outputs\[5\]\[3\]
+ _2082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7625__A2 _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5043_ _1109_ _1207_ _1212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_225_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_100_i_clk clknet_4_13__leaf_i_clk clknet_leaf_100_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7389__A1 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8117__B _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5239__I1 core_0.ew_data\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8802_ core_0.execute.pc_high_buff_out\[0\] _4329_ _4330_ _4324_ _4331_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6416__I _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5320__I _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6994_ _2710_ _2923_ _2924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5939__A2 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Left_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6061__B2 core_0.execute.rf.reg_outputs\[3\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8733_ _1249_ _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_125_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_2655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ core_0.execute.rf.reg_outputs\[1\]\[10\] _1779_ _1804_ core_0.execute.rf.reg_outputs\[11\]\[10\]
+ _1935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_179_2666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_115_i_clk clknet_4_7__leaf_i_clk clknet_leaf_115_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_177_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8631__I core_0.dec_wfi vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8664_ _1658_ _4228_ _4231_ _0566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_192_2811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5876_ _1760_ _1865_ _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_192_2822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7615_ core_0.execute.rf.reg_outputs\[14\]\[2\] _3477_ _3467_ _3480_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4827_ core_0.decode.input_valid _1007_ _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_8595_ net200 _4165_ _4171_ _4172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclone39 _1769_ _1829_ _1858_ _1862_ net267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_7_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7546_ net31 _1348_ _3425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4758_ core_0.ew_reg_ie\[10\] _0928_ _0931_ core_0.ew_reg_ie\[11\] _0930_ core_0.ew_reg_ie\[9\]
+ _0939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_172_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7691__B _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8279__S _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7313__A1 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7477_ core_0.dec_rf_ie\[7\] core_0.ew_reg_ie\[7\] _3366_ _3372_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6116__A2 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8510__B1 _3040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4689_ core_0.execute.rf.reg_outputs\[7\]\[1\] net296 net284 core_0.execute.rf.reg_outputs\[13\]\[1\]
+ _0873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9216_ _0227_ clknet_leaf_79_i_clk net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_133_Left_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6428_ _2393_ _2385_ _2394_ _0167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7864__A2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5875__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4678__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9147_ _0159_ clknet_leaf_98_i_clk core_0.execute.alu_mul_div.div_cur\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6359_ _2219_ _2332_ _2333_ _0159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_112_1857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8813__A1 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7616__A2 _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9078_ _0103_ clknet_leaf_114_i_clk core_0.decode.i_instr_l\[14\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_216_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5627__A1 _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5478__I1 net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8029_ core_0.execute.rf.reg_outputs\[3\]\[1\] _3716_ _3718_ _3719_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_215_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_141_2209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_205_2976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5230__I _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8041__A2 _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7866__B _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4602__A2 net297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_1986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_3317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer101_I core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7552__A1 _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_120_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_2338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7304__A1 _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6107__A2 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8501__B1 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_94_i_clk clknet_4_13__leaf_i_clk clknet_leaf_94_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7855__A2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5866__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4669__A2 net318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7607__A2 _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_3457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8804__A1 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5618__A1 _1060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_2467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_45_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8032__A2 _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5140__I _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_32_i_clk clknet_4_8__leaf_i_clk clknet_leaf_32_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_18_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6043__A1 core_0.execute.rf.reg_outputs\[15\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__B2 core_0.execute.rf.reg_outputs\[7\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7776__B _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ _1714_ _1724_ _0139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_47_i_clk clknet_4_10__leaf_i_clk clknet_leaf_47_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5661_ core_0.execute.alu_mul_div.cbit\[1\] _1669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__7067__I _2829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7400_ _1885_ _3316_ _3318_ _2146_ _3319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9128__CLK clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ core_0.execute.rf.reg_outputs\[10\]\[7\] net221 net220 core_0.execute.rf.reg_outputs\[9\]\[7\]
+ _0802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8380_ _3832_ _3991_ _3992_ _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_174_2596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5592_ _1136_ core_0.decode.i_instr_l\[10\] _1368_ _1627_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7331_ _2939_ _3069_ _3247_ _3251_ _3252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_142_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4543_ core_0.execute.rf.reg_outputs\[6\]\[13\] _0670_ _0710_ core_0.execute.rf.reg_outputs\[8\]\[13\]
+ _0739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8099__A2 _3394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8400__B _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7262_ _1885_ _2424_ _2465_ core_0.decode.oc_alu_mode\[6\] _3184_ _3185_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_96_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4474_ _0668_ net301 _0671_ _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_96_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9001_ _0028_ clknet_leaf_135_i_clk core_0.dec_r_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__5857__A1 net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6213_ _2151_ _2161_ _2201_ _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_40_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7193_ core_0.execute.alu_mul_div.div_res\[9\] _3118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_209_3021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ _2131_ _1685_ _2134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_110_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A1 _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8271__A2 _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6075_ core_0.execute.rf.reg_outputs\[9\]\[6\] net224 _1818_ core_0.execute.rf.reg_outputs\[12\]\[6\]
+ _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_127_2031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ core_0.fetch.prev_request_pc\[6\] _1149_ core_0.fetch.prev_request_pc\[7\]
+ _1198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_212_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__I0 core_0.de_jmp_pred vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4832__A2 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8023__A2 _3394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer73_I core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7231__B1 _3152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6977_ _2497_ _2906_ _2512_ _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_49_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8716_ net76 _1740_ _1730_ _4203_ _4274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_165_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5928_ core_0.execute.rf.reg_outputs\[15\]\[8\] _0944_ _1778_ core_0.execute.rf.reg_outputs\[1\]\[8\]
+ _1918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_165_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8647_ _0900_ _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5859_ _1846_ _1848_ _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_134_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5545__B1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8578_ _3188_ _4156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_161_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7529_ _3397_ _3409_ _3410_ _0252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output187_I net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7837__A2 _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5848__A1 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_235_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4520__A1 core_0.execute.rf.reg_outputs\[6\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8262__A2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4823__A2 net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_240_3387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8014__A2 _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_3398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__A1 _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7773__A1 _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__I core_0.decode.oc_alu_mode\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_183_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4587__A1 core_0.execute.rf.reg_outputs\[5\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7525__A1 _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__A2 _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_229_Left_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7828__A2 _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6500__A2 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5303__A3 net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4511__A1 _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8446__I _2136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8253__A2 _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_238_Left_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_234_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6264__A1 _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4814__A2 _0927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_167_Right_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6900_ _2700_ _2785_ _2831_ _2832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8005__A2 _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7880_ _3415_ _3628_ _3632_ _0381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6016__A1 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6831_ _2712_ core_0.execute.alu_mul_div.i_div _2762_ _2763_ _2764_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_187_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7764__A1 core_0.execute.rf.reg_outputs\[10\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6567__A2 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9550_ _0560_ clknet_leaf_134_i_clk core_0.execute.alu_flag_reg.o_d\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_176_2625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6762_ _2688_ _2689_ _2690_ _2695_ _2696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_119_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8501_ net288 _4048_ _2994_ _2133_ _3002_ _4089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_73_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5713_ net205 _1697_ _1700_ core_0.execute.sreg_priv_control.o_d\[6\] _1713_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_174_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9481_ _0491_ clknet_leaf_16_i_clk net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6693_ net132 _2616_ _2633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7516__A1 net21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8432_ _4016_ _4031_ _4032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5644_ _1079_ _1497_ _0896_ _1084_ _0120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_155_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_215_3091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8363_ _1999_ _3827_ _3974_ _3976_ _3977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8130__B _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5575_ _1143_ _1615_ _1618_ _0090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7314_ _3233_ _3235_ _3236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4526_ _0717_ _0718_ _0721_ _0722_ _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4750__A1 _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7819__A2 _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8294_ core_0.execute.alu_mul_div.mul_res\[7\] _3912_ _3863_ _3913_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_142_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7245_ core_0.ew_data\[10\] _3168_ _3169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_229_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_187_2754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7176_ _2730_ _2720_ _1329_ _3101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6127_ _2076_ _2116_ _1884_ _2117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_225_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5058__A2 _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6255__A1 _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6058_ core_0.execute.rf.reg_outputs\[15\]\[7\] _0944_ _1778_ core_0.execute.rf.reg_outputs\[1\]\[7\]
+ _2048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xclkbuf_3_0_0_i_clk clknet_0_i_clk clknet_3_0_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4805__A2 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5009_ _1180_ _1165_ _1184_ _1162_ net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XPHY_EDGE_ROW_134_Right_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_202_2935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7755__A1 core_0.execute.rf.reg_outputs\[11\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output102_I net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_198_2883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_198_2894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_1956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7507__A1 core_0.ew_reg_ie\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8180__A1 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8040__B _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6730__A2 _2660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5297__A2 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_242_3416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5049__A2 _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__A1 _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6797__A2 _1925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7994__A1 _3414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_2437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_101_Right_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8215__B core_0.execute.alu_mul_div.mul_res\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6549__A2 _2438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7746__A1 _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5221__A2 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4980__A1 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8171__A1 _3469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_171_2566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ core_0.decode.i_instr_l\[9\] core_0.decode.i_instr_l\[8\] _1440_ _1474_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_2_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8885__B _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_236_Right_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5291_ core_0.dec_sreg_store _1411_ _1412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_227_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6485__A1 net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5288__A2 net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7030_ net82 _2829_ _2958_ _2893_ _2959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8226__A2 _2740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9316__CLK clknet_leaf_3_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8981_ _1497_ _4458_ _0656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_124_2001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6788__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7985__A1 _3472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_2695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7932_ _3451_ _3651_ _3662_ _0403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4799__A1 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5460__A2 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7863_ _3460_ _3607_ _3622_ _0374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7737__A1 _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9602_ _0612_ clknet_leaf_60_i_clk core_0.execute.pc_high_out\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6814_ _2076_ _2115_ _2746_ _2747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_147_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7794_ _3470_ _3564_ _3582_ _0345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_3120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9533_ _0543_ clknet_leaf_69_i_clk net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_133_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6745_ _2674_ _2677_ _2678_ _2679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_107_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7456__S _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6960__A2 _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4971__A1 core_0.fetch.prev_request_pc\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9464_ _0474_ clknet_leaf_146_i_clk core_0.execute.rf.reg_outputs\[2\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6676_ _2422_ _2615_ _2617_ _0191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer36_I _1835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8162__A1 _3456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8415_ _4015_ _4020_ core_0.execute.alu_mul_div.div_res\[3\] _4021_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5627_ _1029_ _1628_ _1649_ _0111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9395_ _0405_ clknet_leaf_10_i_clk core_0.execute.rf.reg_outputs\[6\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4723__A1 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8346_ core_0.execute.alu_mul_div.mul_res\[10\] _3943_ _3961_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5558_ core_0.fetch.prev_request_pc\[11\] _1082_ _1083_ net162 _1609_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_115_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input63_I i_req_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ core_0.dec_r_reg_sel\[1\] _0675_ _0684_ _0707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__8465__A2 _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8277_ _3893_ _3895_ _3896_ _3897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_203_Right_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5489_ _1569_ _1551_ _1570_ _0052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7228_ _1290_ _3150_ _3151_ _1742_ _3152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_57_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7159_ _3083_ _3084_ _3085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__6228__A1 _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_109_1818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_2270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7976__A1 _3459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5987__B1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5451__A2 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7728__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer70 net271 net298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_197_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer81 _0685_ net309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_139_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer92 _1803_ net339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_95_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5739__B1 _1730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6400__A1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6951__A2 _2881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8689__C _4249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4962__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8153__A1 net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7900__A1 _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8456__A2 _4048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6467__A1 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9339__CLK clknet_leaf_155_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8208__A2 _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7967__A1 core_0.execute.rf.reg_outputs\[5\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5978__B1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__B1 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4860_ core_0.fetch.out_buffer_data_instr\[17\] _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_169_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8231__I2 _2115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8392__A1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7195__A2 _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7784__B _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4791_ core_0.ew_reg_ie\[12\] _0948_ _0971_ _0972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6942__A2 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _2470_ _2471_ _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_144_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8144__A1 _3414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_31_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6461_ _2413_ _0905_ _0181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8200_ core_0.execute.alu_mul_div.mul_res\[0\] _3825_ _3826_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5412_ core_0.decode.i_instr_l\[13\] _1509_ _1510_ core_0.decode.i_instr_l\[9\] _1495_
+ _1513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_140_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9180_ _0191_ clknet_leaf_46_i_clk core_0.ew_addr_high\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_212_3061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6392_ _2365_ _1962_ _1955_ _2366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xoutput102 net102 dbg_r0[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput113 net113 o_instr_long_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput124 net124 o_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8131_ _3465_ _3760_ _3776_ _0488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5343_ _1448_ _1453_ _1456_ _1460_ _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_88_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput135 net135 o_mem_addr_high[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8447__A2 _1737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput146 net146 o_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5524__S _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput157 net157 o_mem_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput168 net168 o_req_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_130_2071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput179 net179 sr_bus_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_195_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8062_ _3736_ _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5274_ core_0.de_jmp_pred _1394_ _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_184_2724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7013_ _2040_ _2755_ _2433_ core_0.decode.oc_alu_mode\[9\] _2942_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_227_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7958__A1 core_0.execute.rf.reg_outputs\[5\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8964_ net182 core_0.decode.i_imm_pass\[14\] _1263_ _4450_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_223_3190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clone56_I _0707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5433__A2 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_93_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7915_ _3402_ _3651_ _3653_ _0395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8895_ net114 _4383_ _4409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_214_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6154__I _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7846_ _3605_ _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_104_1759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7186__A2 _3069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_195_2853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5197__A1 _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7777_ _3441_ _3563_ _3573_ _0337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4989_ _1156_ _1167_ _1168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_191_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6728_ net136 _2642_ _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9516_ _0526_ clknet_leaf_118_i_clk core_0.execute.alu_mul_div.div_res\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xwire218 _2025_ net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__8135__A1 _3472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9447_ _0457_ clknet_leaf_145_i_clk core_0.execute.rf.reg_outputs\[3\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6659_ _2588_ _2598_ _2599_ _2600_ _2587_ _2601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_6_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9378_ _0388_ clknet_leaf_32_i_clk core_0.execute.rf.reg_outputs\[7\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_103_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8329_ _3944_ _3945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__8438__A2 _4031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6449__A1 _1180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_3219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5121__A1 _1244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6621__A1 net325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5424__A2 _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4632__B1 net308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8374__A1 core_0.execute.alu_mul_div.mul_res\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_237_3359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A1 core_0.decode.oc_alu_mode\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4935__B2 core_0.fetch.prev_request_pc\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8212__C core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput15 i_core_int_sreg[8] net15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_155_2369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput26 i_mem_data[14] net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput37 i_mem_exception net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8677__A2 _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput48 i_req_data[1] net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput59 i_req_data[2] net59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6688__A1 net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4699__B1 net284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5360__A1 core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7101__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_179_Left_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_224_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5663__A2 _1670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6683__B net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4982__I _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_115_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8454__I _4046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5415__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ core_0.execute.rf.reg_outputs\[1\]\[11\] _1779_ _1804_ core_0.execute.rf.reg_outputs\[11\]\[11\]
+ _1951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_177_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7700_ _3435_ _3520_ _3529_ _0304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4912_ core_0.fetch.prev_request_pc\[11\] _1057_ _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8680_ _1658_ _4241_ _4244_ _0569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_181_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5892_ _1757_ _1882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_87_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5179__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7631_ core_0.execute.rf.reg_outputs\[14\]\[9\] _3482_ _3486_ _3489_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4843_ core_0.fetch.out_buffer_data_instr\[29\] _1024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_188_Left_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7562_ _3381_ _3437_ _3438_ _3439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_74_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8117__A1 core_0.execute.rf.reg_outputs\[1\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ core_0.dec_l_reg_sel\[0\] _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_9301_ _0311_ clknet_leaf_153_i_clk core_0.execute.rf.reg_outputs\[12\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6513_ _2443_ _2451_ _2454_ _2440_ _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_71_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7493_ core_0.dec_rf_ie\[15\] core_0.ew_reg_ie\[15\] _2421_ _3380_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9232_ _0243_ clknet_leaf_142_i_clk core_0.ew_reg_ie\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_190_2794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6444_ core_0.execute.mem_stage_pc\[9\] _2395_ _2404_ _2405_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7340__A2 _3259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9163_ _0174_ clknet_leaf_82_i_clk core_0.execute.mem_stage_pc\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5351__A1 _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6375_ _2347_ _1962_ _2348_ _2349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_246_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8114_ _3434_ _3759_ _3767_ _0480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_228_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5326_ _1234_ _1258_ _1256_ _1236_ _1444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_197_Left_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_9094_ _0119_ clknet_leaf_91_i_clk core_0.decode.i_imm_pass\[15\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8045_ _3450_ _3715_ _3727_ _0451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5103__A1 _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5257_ _1376_ core_0.execute.alu_flag_reg.o_d\[1\] _1378_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8840__A2 _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6851__A1 _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7689__B _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5188_ core_0.decode.oc_alu_mode\[13\] _1251_ _1293_ _1333_ _1334_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input26_I i_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8947_ _1850_ _0038_ _4441_ _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4614__B1 net316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8878_ _4386_ _4395_ _4396_ _0615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8356__A1 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7829_ _3466_ _3586_ _3602_ _0360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8108__A1 core_0.execute.rf.reg_outputs\[1\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5590__A1 _1135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5228__I _1359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output94_I net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7331__A2 _3069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5342__A1 _1276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__C _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_12__f_i_clk clknet_3_6_0_i_clk clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6842__A1 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_201_Left_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8595__A1 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4605__B1 net286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6070__A2 net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_210_Left_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_182_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7570__A2 core_0.ew_data\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_231_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5581__A1 _1139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4490_ core_0.dec_r_reg_sel\[1\] _0664_ _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_12_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5333__A1 _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5884__A2 _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_2527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6160_ core_0.execute.alu_mul_div.div_cur\[13\] _1837_ _2149_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_110_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8893__B _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5111_ core_0.decode.i_instr_l\[6\] core_0.decode.i_instr_l\[4\] core_0.decode.i_instr_l\[5\]
+ _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_237_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6091_ core_0.execute.rf.reg_outputs\[10\]\[3\] _1780_ net338 core_0.execute.rf.reg_outputs\[11\]\[3\]
+ net330 core_0.execute.rf.reg_outputs\[4\]\[3\] _2081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_176_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5636__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5042_ net81 _1211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_224_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7389__A2 net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8801_ core_0.execute.pc_high_out\[0\] _4329_ _4330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6993_ core_0.execute.alu_mul_div.div_cur\[4\] core_0.execute.alu_mul_div.i_mod _2920_
+ _2922_ _2923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__6061__A2 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5944_ core_0.execute.rf.reg_outputs\[6\]\[10\] net322 _1819_ core_0.execute.rf.reg_outputs\[12\]\[10\]
+ _1788_ core_0.execute.rf.reg_outputs\[3\]\[10\] _1934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_8732_ core_0.execute.sreg_jtr_buff.o_d\[2\] _4217_ _4283_ _4286_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_2656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8338__A1 _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8663_ _4212_ core_0.execute.mem_stage_pc\[4\] _4202_ _4230_ _4231_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_164_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8889__A2 _4385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5875_ _1769_ _1812_ _1864_ _1865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_101_1729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_192_2812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7010__A1 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7614_ _3409_ _3476_ _3479_ _0268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4826_ _0925_ _1006_ _1007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_145_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8594_ net211 _4165_ _4171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclone29 _0709_ net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_90_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7545_ net24 _1347_ _3424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4757_ core_0.ew_reg_ie\[8\] _0665_ net271 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5572__A1 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7464__S _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7476_ _3371_ _0238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4780__C1 _0960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ core_0.execute.rf.reg_outputs\[5\]\[1\] _0677_ net347 core_0.execute.rf.reg_outputs\[15\]\[1\]
+ _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8510__A1 net277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8510__B2 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9215_ _0226_ clknet_leaf_77_i_clk net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6427_ core_0.execute.mem_stage_pc\[3\] _2386_ _2387_ _2394_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5875__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9146_ _0158_ clknet_leaf_97_i_clk core_0.execute.alu_mul_div.div_cur\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6358_ core_0.execute.alu_mul_div.div_cur\[15\] _2218_ _0999_ _2333_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_1858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5309_ _1371_ _1429_ _0923_ _0013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9077_ _0102_ clknet_leaf_100_i_clk core_0.decode.i_instr_l\[13\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__8813__A2 _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6289_ _2258_ _2272_ _0150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5627__A2 _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8028_ _3647_ _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8577__A1 _3293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_205_2977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4571__B _0764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_234_3318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7001__A1 _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7552__A2 _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5563__A1 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_2339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7304__A2 _3225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8501__A1 net288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8501__B2 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5315__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5866__A2 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_148_Right_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_245_3447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_245_3458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6718__S _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8804__A2 _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6945__C _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6815__A1 _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5618__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8218__B _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_234_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_2468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5421__I _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8568__A1 _4080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__B1 _1916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7240__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6043__A2 _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7791__A2 _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5577__B _1619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ core_0.execute.alu_mul_div.cbit\[0\] _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_139_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8740__A1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7543__A2 _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4611_ _0801_ net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__5554__A1 _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5591_ _1439_ core_0.fetch.submitable _1626_ _0098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_2597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7330_ _1885_ _2473_ _3248_ _1880_ _3250_ _3251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_13_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ core_0.execute.rf.reg_outputs\[7\]\[13\] net296 _0703_ core_0.execute.rf.reg_outputs\[15\]\[13\]
+ _0738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7261_ _1956_ _3072_ _3183_ net265 _3073_ _3184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__5306__A1 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ _0662_ _0660_ _0671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_111_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9000_ _0027_ clknet_leaf_133_i_clk core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_96_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4500__I _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6212_ _2162_ _2200_ _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7192_ _1743_ _3115_ _3116_ _0996_ _3117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_96_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_209_3022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_115_Right_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6143_ _2132_ _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_237_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6806__A1 _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A2 net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6074_ core_0.execute.rf.reg_outputs\[14\]\[6\] _1801_ _1803_ core_0.execute.rf.reg_outputs\[11\]\[6\]
+ _2064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_224_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8128__B _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5025_ _1086_ _1196_ _1197_ _1162_ net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_212_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8559__A1 net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7967__B _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7231__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6976_ _2845_ _2847_ _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_rebuffer66_I net197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7782__A2 _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8715_ _4272_ _4273_ _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5793__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5927_ core_0.execute.rf.reg_outputs\[5\]\[8\] net225 net226 core_0.execute.rf.reg_outputs\[10\]\[8\]
+ net336 core_0.execute.rf.reg_outputs\[2\]\[8\] _1917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_193_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5858_ _1754_ net207 _1847_ _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_152_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8646_ _1658_ _4211_ _4216_ _0563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_63_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5545__A1 core_0.fetch.prev_request_pc\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _0971_ _0943_ _0988_ _0989_ _0990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_91_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_17_Right_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5545__B2 net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8577_ _3293_ _3330_ _4155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5789_ _1778_ _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4753__C1 _0930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7528_ core_0.execute.rf.reg_outputs\[15\]\[1\] _3403_ _2404_ _3410_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7459_ _3362_ _0230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5848__A2 _1833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4520__A2 _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9129_ _0141_ clknet_leaf_104_i_clk core_0.execute.sreg_priv_control.o_d\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_228_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_26_Right_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8038__B _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__C2 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_215_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_9_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7877__B _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_3388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7222__A1 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7222__B2 core_0.decode.oc_alu_mode\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7773__A2 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5784__A1 core_0.execute.rf.reg_outputs\[7\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4587__A2 net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8722__A1 _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_217_Right_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__A4 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_114_i_clk clknet_4_7__leaf_i_clk clknet_leaf_114_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_207_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_152_Left_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_237_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_129_i_clk clknet_4_4__leaf_i_clk clknet_leaf_129_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_173_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7213__A1 _2528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6830_ _2124_ core_0.execute.alu_mul_div.mul_res\[1\] core_0.execute.alu_mul_div.i_div
+ _2763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7764__A2 _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5775__A1 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4578__A2 _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6761_ _2691_ _2692_ _2693_ _2694_ _2695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_176_2626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_53_Right_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8500_ _4039_ _4087_ _4088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5712_ _1608_ _1712_ _0133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _2628_ _2631_ _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_9480_ _0490_ clknet_leaf_144_i_clk core_0.execute.rf.reg_outputs\[1\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7516__A2 _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8713__A1 _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5790__A4 core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5643_ _1023_ _1628_ _1657_ _0119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8431_ _1537_ _2215_ _2216_ _4031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_33_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8362_ _3828_ _3975_ _3976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5574_ _1232_ _1616_ _1618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_215_3092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7313_ _2699_ _3234_ _3235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4525_ core_0.execute.rf.reg_outputs\[7\]\[14\] net296 _0686_ core_0.execute.rf.reg_outputs\[14\]\[14\]
+ _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8293_ _2054_ _3827_ _3911_ _3912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4750__A2 _0675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7244_ _2421_ _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__9395__CLK clknet_leaf_10_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Right_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_187_2755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7175_ _3099_ _2457_ _3100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7541__I _3420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6126_ _1899_ _2115_ _2116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6057_ core_0.execute.rf.reg_outputs\[5\]\[7\] net225 net226 core_0.execute.rf.reg_outputs\[10\]\[7\]
+ net336 core_0.execute.rf.reg_outputs\[2\]\[7\] _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__5061__I net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _1181_ _1146_ _1183_ _1164_ _1184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_213_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6007__A2 _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7204__A1 _2710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_202_2936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_71_Right_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7755__A2 _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8952__A1 core_0.decode.i_imm_pass\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_93_i_clk clknet_4_13__leaf_i_clk clknet_leaf_93_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_198_2884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5766__A1 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ core_0.execute.pc_high_buff_out\[4\] _2771_ _2775_ core_0.execute.pc_high_out\[4\]
+ _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5518__A1 net56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8629_ _0900_ _4200_ _4201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XANTENNA__6715__B1 _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8180__A2 _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6191__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5236__I _1363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_80_Right_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_88_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_31_i_clk clknet_4_8__leaf_i_clk clknet_leaf_31_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7691__A1 core_0.execute.rf.reg_outputs\[12\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_242_3417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_0__f_i_clk clknet_3_0_0_i_clk clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_46_i_clk clknet_4_10__leaf_i_clk clknet_leaf_46_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7443__A1 _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9118__CLK clknet_leaf_64_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7994__A2 _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_2427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_2438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7746__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8943__A1 _1687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5757__A1 _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9268__CLK clknet_leaf_7_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6706__B1 _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7626__I _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8171__A2 _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_171_2567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5290_ _1405_ net227 _1410_ _1411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_50_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6485__A2 net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5288__A3 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_160_Left_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4496__A1 _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7434__A1 net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6237__A2 _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6906__S _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8980_ core_0.dec_rf_ie\[1\] _1482_ _1462_ _1474_ _4458_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_207_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7985__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_2696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7931_ core_0.execute.rf.reg_outputs\[6\]\[8\] _3657_ _3648_ _3662_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5996__A1 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4799__A2 _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7862_ core_0.execute.rf.reg_outputs\[8\]\[11\] _3613_ _3621_ _3622_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8934__A1 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7737__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9601_ _0611_ clknet_leaf_50_i_clk core_0.execute.pc_high_out\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_77_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5748__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6813_ _2503_ _2504_ _2746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6945__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7793_ core_0.execute.rf.reg_outputs\[10\]\[14\] _3562_ _3580_ _3582_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_217_3121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9532_ _0542_ clknet_leaf_103_i_clk net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_18_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6744_ _1226_ _1405_ net227 _1410_ _2678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_147_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ core_0.ew_addr_high\[0\] _2616_ _2617_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9463_ _0473_ clknet_leaf_146_i_clk core_0.execute.rf.reg_outputs\[2\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4971__A2 core_0.fetch.prev_request_pc\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8141__B _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8162__A2 _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5626_ core_0.decode.i_imm_pass\[7\] _1645_ _1649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8414_ _2140_ _1670_ _4020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_135_2131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9394_ _0404_ clknet_leaf_26_i_clk core_0.execute.rf.reg_outputs\[6\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_rebuffer29_I _1798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7980__B _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4723__A2 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8345_ _3958_ _3959_ _3960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5557_ _1253_ _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_14_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4508_ core_0.execute.rf.reg_outputs\[15\]\[15\] _0703_ _0705_ core_0.execute.rf.reg_outputs\[9\]\[15\]
+ _0706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8276_ _3893_ _3895_ _3802_ _3896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5488_ net41 _1554_ _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input56_I i_req_data[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7227_ _1290_ core_0.execute.alu_mul_div.mul_res\[10\] _3151_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_228_3250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4487__A1 _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7158_ core_0.execute.alu_mul_div.div_cur\[8\] _0997_ _3084_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_70_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7425__A1 _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ core_0.execute.rf.reg_outputs\[13\]\[2\] _1792_ _1799_ core_0.execute.rf.reg_outputs\[6\]\[2\]
+ _2099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6228__A2 _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7089_ _2439_ _3014_ _3015_ _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_109_1819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_2260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7976__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5987__A1 core_0.execute.rf.reg_outputs\[8\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5987__B2 core_0.execute.rf.reg_outputs\[4\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9410__CLK clknet_leaf_37_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5451__A3 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer60 _0825_ net288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__7728__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer71 net298 net299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer82 net309 net310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_25_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer93 _1786_ net340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5739__A1 core_0.execute.sreg_priv_control.o_d\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5739__B2 _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8051__B _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8153__A2 _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7900__A2 _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7113__B1 _3037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6467__A2 _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7664__A1 core_0.execute.rf.reg_outputs\[13\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4478__A1 _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7416__A1 _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7967__A2 _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_1_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__B2 core_0.execute.rf.reg_outputs\[14\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8916__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4650__A1 core_0.execute.rf.reg_outputs\[11\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__B2 core_0.execute.rf.reg_outputs\[9\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8231__I3 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ core_0.dec_l_reg_sel\[3\] _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_28_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8144__A2 _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6260__I _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6460_ _2413_ _0908_ _0180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_31_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6155__A1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8896__B _4385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_111_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5411_ _0954_ _1486_ _1512_ _1501_ _0031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_212_3051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_212_3062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6391_ net89 _2365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5902__A1 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4705__A2 _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5902__B2 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput103 net103 o_c_data_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8130_ core_0.execute.rf.reg_outputs\[1\]\[13\] _3765_ _3771_ _3776_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput114 net114 o_instr_long_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5342_ _1276_ _1457_ _1459_ _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xoutput125 net125 o_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput136 net136 o_mem_addr_high[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput147 net147 o_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_140_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput158 net158 o_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8061_ core_0.ew_reg_ie\[2\] _3394_ _3736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7655__A1 core_0.execute.rf.reg_outputs\[13\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6458__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput169 net169 o_req_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5273_ _1372_ _1385_ _1393_ _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_130_2072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_184_2725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7012_ _1337_ _2040_ core_0.decode.oc_alu_mode\[7\] _2941_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_195_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5418__B1 _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_207_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7958__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5969__A1 _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8963_ _4449_ _0647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_223_3191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7914_ core_0.execute.rf.reg_outputs\[6\]\[0\] _3652_ _3648_ _3653_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5433__A3 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8894_ _4386_ _4407_ _4408_ _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_195_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8907__A1 core_0.dec_sys vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7975__B _3677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7845_ _3421_ _3606_ _3612_ _0366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_194_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7467__S _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_195_2854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6394__A1 _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7776_ core_0.execute.rf.reg_outputs\[10\]\[6\] _3570_ _3568_ _3573_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4988_ _1158_ _1166_ _1167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9515_ _0525_ clknet_leaf_117_i_clk core_0.execute.alu_mul_div.div_res\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6727_ _2660_ _2662_ _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_19_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8135__A2 _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6146__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9446_ _0456_ clknet_leaf_145_i_clk core_0.execute.rf.reg_outputs\[3\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6658_ _1875_ _2588_ _2600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_59_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6697__A2 _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7894__A1 _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5609_ _1591_ net43 _1369_ _1639_ _1640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_9377_ _0387_ clknet_leaf_39_i_clk core_0.execute.rf.reg_outputs\[7\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6589_ _2523_ _2530_ _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8328_ core_0.execute.alu_mul_div.mul_res\[10\] _3943_ _3944_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_103_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output162_I net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6449__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8259_ _3878_ _3879_ _3880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_218_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8071__A1 _3420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8046__B _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4632__A1 core_0.execute.rf.reg_outputs\[14\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4632__B2 core_0.execute.rf.reg_outputs\[1\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_201_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_wire211_I _2606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5188__A2 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__A2 _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8126__A2 _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput16 i_core_int_sreg[9] net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput27 i_mem_data[15] net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__9306__CLK clknet_leaf_1_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput38 i_req_data[0] net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_24_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput49 i_req_data[20] net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7885__A1 _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4699__A1 core_0.execute.rf.reg_outputs\[7\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5360__A2 core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7637__A1 core_0.execute.rf.reg_outputs\[14\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_2499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__B1 _1778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5960_ core_0.execute.rf.reg_outputs\[15\]\[11\] _0945_ _1821_ core_0.execute.rf.reg_outputs\[7\]\[11\]
+ _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_149_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4623__A1 net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7795__B _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4911_ core_0.fetch.prev_request_pc\[12\] _1020_ _1057_ core_0.fetch.prev_request_pc\[11\]
+ _1091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_5891_ _1880_ _1876_ _1881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8365__A2 _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7630_ _3451_ _3476_ _3488_ _0275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4842_ _0892_ net61 _1022_ _1023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_114_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7561_ net33 _1348_ _3438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4773_ _0953_ _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_117_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8117__A2 _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9300_ _0310_ clknet_leaf_6_i_clk core_0.execute.rf.reg_outputs\[12\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6128__A1 _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6512_ _2434_ _2452_ _2453_ _2454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_160_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7492_ _3379_ _0246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9231_ _0242_ clknet_leaf_142_i_clk core_0.ew_reg_ie\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7876__A1 _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6443_ _1430_ _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_113_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_2795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6374_ _2080_ _2089_ _2348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9162_ _0173_ clknet_leaf_70_i_clk core_0.execute.mem_stage_pc\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8113_ core_0.execute.rf.reg_outputs\[1\]\[5\] _3765_ _3756_ _3767_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5325_ _1244_ _1442_ _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7628__A1 _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7479__I1 core_0.ew_reg_ie\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9093_ _0118_ clknet_leaf_91_i_clk core_0.decode.i_imm_pass\[14\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8044_ core_0.execute.rf.reg_outputs\[3\]\[8\] _3722_ _3718_ _3727_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_54_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5256_ _1376_ _1374_ _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6300__A1 _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6851__A2 core_0.execute.sreg_irq_pc.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5187_ _1236_ _1256_ _1258_ _1295_ _1316_ _1333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4862__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_rebuffer96_I _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8053__A1 core_0.execute.rf.reg_outputs\[3\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_2230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input19_I i_mc_core_int vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7800__A1 core_0.execute.rf.reg_outputs\[9\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8946_ core_0.decode.i_imm_pass\[5\] _1264_ _4441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4614__B2 core_0.execute.rf.reg_outputs\[8\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8877_ core_0.execute.pc_high_buff_out\[2\] _4385_ _3797_ _4396_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_195_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7828_ core_0.execute.rf.reg_outputs\[9\]\[13\] _3591_ _3595_ _3602_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_65_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7759_ core_0.ew_reg_ie\[10\] _3395_ _3562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_81_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8108__A2 _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_129_Right_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5590__A2 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9429_ _0439_ clknet_leaf_144_i_clk core_0.execute.rf.reg_outputs\[4\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9479__CLK clknet_leaf_144_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7867__A1 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7724__I _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output87_I net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8292__A1 _3901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6842__A2 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8044__A1 core_0.execute.rf.reg_outputs\[3\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4605__B2 core_0.execute.rf.reg_outputs\[13\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8347__A2 _3947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_4__f_i_clk_I clknet_3_2_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6358__A1 core_0.execute.alu_mul_div.div_cur\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__A1 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5581__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5863__B _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7858__A1 _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4541__B1 _0693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_2528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5110_ _1253_ _1254_ _1229_ _1256_ _1265_ _0009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_176_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8283__A1 _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6090_ _1770_ _2077_ _2078_ _2079_ _2080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5041_ _1206_ _1165_ _1209_ _1210_ _1080_ net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_85_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Left_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6833__A2 _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4844__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6046__B1 net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8800_ _0901_ _1415_ _4329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_220_3150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6992_ _2921_ core_0.execute.alu_mul_div.i_div core_0.execute.alu_mul_div.i_mod _2922_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8731_ _4214_ _4283_ _4285_ _1501_ _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_220_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5943_ _1931_ _1932_ _1933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_149_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_179_2657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8662_ _4224_ _4070_ _4229_ _1662_ _4230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_87_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5874_ _1863_ _1864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_146_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_192_2813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7613_ core_0.execute.rf.reg_outputs\[14\]\[1\] _3477_ _3467_ _3479_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_38_Left_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4825_ _0926_ _0995_ _1005_ _1006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5021__A1 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8593_ _4169_ _4170_ _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9621__CLK clknet_leaf_133_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7544_ _3397_ _3421_ _3423_ _0254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_173_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4756_ core_0.ew_reg_ie\[12\] _0665_ _0930_ core_0.ew_reg_ie\[13\] _0931_ core_0.ew_reg_ie\[15\]
+ _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__5572__A2 _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7475_ core_0.dec_rf_ie\[6\] core_0.ew_reg_ie\[6\] _3366_ _3371_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4687_ core_0.execute.rf.reg_outputs\[9\]\[1\] _0705_ net257 core_0.execute.rf.reg_outputs\[8\]\[1\]
+ _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4780__C2 core_0.ew_reg_ie\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8510__A2 _4048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9214_ _0225_ clknet_leaf_77_i_clk net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_231_3290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6426_ net80 _2393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_141_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9145_ _0157_ clknet_leaf_98_i_clk core_0.execute.alu_mul_div.div_cur\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5064__I _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6357_ _2331_ _2142_ _2246_ _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8274__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5308_ core_0.dec_jump_cond_code\[4\] _1395_ _1428_ _1413_ _1429_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XPHY_EDGE_ROW_47_Left_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_9076_ _0101_ clknet_leaf_114_i_clk core_0.decode.i_instr_l\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6288_ core_0.execute.alu_mul_div.div_cur\[6\] _2219_ _2271_ _2272_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_227_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5088__A1 core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8027_ _3401_ _3715_ _3717_ _0443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5239_ core_0.ew_data\[7\] core_0.ew_data\[15\] _1349_ _1365_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_242_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8026__A1 core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_242_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8577__A2 _3330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_205_2967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_205_2978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_196_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__B1 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8929_ _4428_ _4430_ _4431_ _4432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__A1 core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7719__I _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_195_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_123_1988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_234_3319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5012__A1 _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5563__A2 _1611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_5_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8501__A2 _4048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5315__A2 core_0.execute.sreg_priv_control.o_d\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5866__A3 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_219_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_245_3448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7403__B _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6815__A2 _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8017__A1 core_0.execute.rf.reg_outputs\[4\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_163_2469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8568__A2 _3335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6579__B2 _1923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5858__B _1847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5003__A1 _1175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8740__A2 _1418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4610_ net101 net324 _0800_ _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_127_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5590_ _1135_ _1369_ _1626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_25_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6751__A1 core_0.execute.sreg_scratch.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_174_2598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4541_ core_0.execute.rf.reg_outputs\[2\]\[13\] _0673_ _0693_ core_0.execute.rf.reg_outputs\[1\]\[13\]
+ _0737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7260_ _1337_ _2366_ core_0.decode.oc_alu_mode\[7\] _3183_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6503__A1 _1753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4472_ _0669_ _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_13_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6211_ core_0.execute.alu_mul_div.div_cur\[10\] _1833_ _2199_ _2200_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_150_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7191_ _2124_ core_0.execute.alu_mul_div.mul_res\[9\] _3116_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_209_3023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _2131_ _1403_ _2132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6073_ core_0.execute.rf.reg_outputs\[15\]\[6\] _0944_ _1778_ core_0.execute.rf.reg_outputs\[1\]\[6\]
+ _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6806__A2 _2115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4817__A1 _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9174__CLK clknet_leaf_42_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5024_ net85 _1085_ _1197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_127_2033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8008__A1 _3450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8559__A2 _4052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_205_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7231__A2 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6975_ core_0.decode.oc_alu_mode\[4\] _2903_ _2904_ _2905_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_76_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8714_ core_0.execute.sreg_irq_pc.o_d\[13\] _4210_ _1431_ _4273_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6443__I _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5926_ core_0.execute.rf.reg_outputs\[7\]\[8\] _1821_ _1915_ _1916_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_165_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6990__A1 _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer59_I _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8645_ _4212_ core_0.execute.mem_stage_pc\[1\] _4202_ _4215_ _4216_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_192_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5857_ net313 _1688_ _1847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_35_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7475__S _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8731__A2 _4283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4808_ core_0.ew_reg_ie\[4\] _0963_ _0964_ core_0.ew_reg_ie\[5\] _0966_ core_0.ew_reg_ie\[6\]
+ _0989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__5545__A2 _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8576_ _3079_ _3115_ _3220_ _3256_ _4154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_145_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6742__A1 net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5788_ _0957_ _0958_ _0951_ _1778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_138_2173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__I core_0.fetch.dbg_out vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7527_ _3408_ _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4753__B1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4739_ core_0.execute.prev_pc_high\[5\] _0917_ _0914_ core_0.execute.prev_pc_high\[6\]
+ _0919_ _0920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_133_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8495__A1 _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7458_ net119 _3297_ _2415_ _3362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_160_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5848__A3 _1835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ core_0.de_jmp_pred core_0.decode.i_jmp_pred_pass _1264_ _2381_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_4_10__f_i_clk_I clknet_3_5_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7389_ _2672_ net198 _3308_ _3309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8247__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9128_ _0140_ clknet_4_12__leaf_i_clk core_0.execute.sreg_priv_control.o_d\[12\]
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9059_ _0085_ clknet_leaf_92_i_clk core_0.fetch.prev_request_pc\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4808__A1 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__B2 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_max_cap219_I _1798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_240_3389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7222__A2 _2155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_64_Left_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_84_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8970__A2 _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6981__A1 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5784__A2 _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7893__B _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_181_Right_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_73_Left_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8238__A1 core_0.execute.alu_mul_div.mul_res\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8789__A2 _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8944__S _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6760_ core_0.dec_sreg_jal_over _2694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_176_2627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5711_ core_0.execute.sreg_priv_control.o_d\[5\] _1701_ _1711_ _1698_ _1712_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_174_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6691_ _2629_ _2630_ _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer9_I net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8430_ _2230_ _4030_ _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5642_ core_0.decode.i_imm_pass\[15\] _1368_ _1657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5527__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4735__B1 net111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8361_ _3958_ _3967_ _3973_ _3975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _1011_ _1615_ _1617_ _0089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_215_3093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7312_ _3201_ _3232_ _3234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8477__A1 _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4524_ core_0.execute.rf.reg_outputs\[4\]\[14\] net318 _0716_ _0721_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8292_ _3901_ _3909_ _3910_ _3911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7243_ _2709_ _3165_ _3166_ _3167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8229__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_2756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5160__B1 _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7174_ _3057_ _2456_ _2461_ _3099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8139__B _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6125_ net94 _1813_ _2109_ _2114_ _2115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__7452__A2 _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6056_ _1771_ _2043_ _2044_ _2045_ _2046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_198_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5007_ _1145_ _1153_ _1182_ _1183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_212_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_106_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_206_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_240_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7204__A2 _3120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_2937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5215__A1 core_0.ew_data\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8952__A2 _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6958_ core_0.execute.sreg_irq_flags.o_d\[4\] _2777_ _2774_ core_0.execute.sreg_irq_pc.o_d\[4\]
+ _2888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__A2 _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_198_2885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5909_ _1882_ _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_48_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_1947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6889_ core_0.execute.alu_mul_div.div_cur\[2\] _1317_ _2818_ _2820_ _2821_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__7507__A3 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8628_ _1419_ _1433_ _3042_ _4200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_8_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5518__A2 _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6715__A1 core_0.execute.rf.reg_outputs\[1\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6715__B2 core_0.execute.rf.reg_outputs\[3\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output192_I net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8559_ net75 _4052_ _4140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_20_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6191__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7140__A1 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7691__A2 _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_242_3418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7443__A2 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8640__A1 core_0.execute.sreg_irq_pc.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5454__A1 _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_243_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_160_2428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5057__I1 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8943__A2 _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6954__A1 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5757__A2 net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8512__B _4051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7907__I _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6706__A1 core_0.execute.rf.reg_outputs\[1\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6706__B2 core_0.execute.rf.reg_outputs\[3\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6182__A2 _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_171_2568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5288__A4 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7682__A2 _3496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4496__A2 _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7434__A2 _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7930_ _3447_ _3651_ _3661_ _0402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_182_2697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7861_ _3512_ _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_89_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5048__I1 _1060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9600_ _0610_ clknet_leaf_49_i_clk core_0.execute.pc_high_out\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6812_ _2006_ _2729_ _2744_ _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_148_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5748__A2 _1737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6945__A1 core_0.execute.sreg_long_ptr_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7792_ _3466_ _3564_ _3581_ _0344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6945__B2 net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9531_ _0541_ clknet_leaf_74_i_clk net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_217_3111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _2675_ _1686_ _1689_ _2676_ _2677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_TAPCELL_ROW_217_3122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9462_ _0472_ clknet_leaf_146_i_clk core_0.execute.rf.reg_outputs\[2\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6674_ _2421_ _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_73_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8413_ _2819_ _4019_ _2258_ _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5625_ _1039_ _1615_ _1648_ _0110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9393_ _0403_ clknet_leaf_33_i_clk core_0.execute.rf.reg_outputs\[6\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7370__A1 _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6173__A2 _1835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8344_ core_0.execute.alu_mul_div.mul_res\[11\] _3957_ _3959_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_131_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5556_ _1597_ _1607_ _0082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_32_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4507_ net220 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__7122__A1 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8275_ core_0.execute.alu_mul_div.mul_res\[6\] _3894_ _3895_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5487_ core_0.fetch.out_buffer_data_instr\[12\] _1569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_218_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7226_ _3133_ _3135_ _3138_ _3149_ _3150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__8870__A1 _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5684__A1 _1687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I i_req_data[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_3251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7157_ core_0.execute.alu_mul_div.div_res\[8\] _1314_ _3080_ _3082_ core_0.execute.alu_mul_div.i_mod
+ _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_67_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7425__A2 _3335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6108_ core_0.execute.rf.reg_outputs\[10\]\[2\] _1781_ _1794_ core_0.execute.rf.reg_outputs\[8\]\[2\]
+ _2098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7088_ _2439_ _3014_ _1292_ _3015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_146_2261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6039_ core_0.execute.rf.reg_outputs\[13\]\[5\] _1791_ _1815_ core_0.execute.rf.reg_outputs\[9\]\[5\]
+ _2029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_241_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5987__A2 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5451__A4 _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer50 _0813_ net278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_200_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer61 net288 net289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_output205_I net279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8925__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer72 _0664_ net300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer83 _2528_ net311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_25_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6936__A1 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5739__A2 _1700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_239_3380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_113_i_clk clknet_4_7__leaf_i_clk clknet_leaf_113_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_36_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8689__A1 _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5247__I _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_128_i_clk clknet_4_4__leaf_i_clk clknet_leaf_128_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5911__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7664__A2 _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5675__A1 _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4478__A2 _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8613__A1 _3188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7416__A2 _3333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A1 _1294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5978__A2 _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_231_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4650__A2 _0680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_5_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6927__A1 _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9385__CLK clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5157__I core_0.decode.oc_alu_mode\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6155__A2 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5410_ core_0.decode.i_instr_l\[12\] _1509_ _1510_ core_0.decode.i_instr_l\[8\] _1495_
+ _1512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_212_3052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6390_ _1544_ _2357_ _2363_ _2364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6697__B net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5902__A2 _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput104 net104 o_c_instr_long vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_140_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput115 net115 o_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5341_ _1331_ _1458_ _1240_ _1459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_140_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput126 net126 o_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput137 net137 o_mem_addr_high[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput148 net148 o_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput159 net159 o_req_active vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8060_ _3472_ _3716_ _3735_ _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7655__A2 _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_92_i_clk clknet_4_15__leaf_i_clk clknet_leaf_92_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5272_ core_0.dec_jump_cond_code\[2\] _1386_ _1377_ _1389_ _1392_ _1393_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_TAPCELL_ROW_130_2073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_2715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7011_ _1759_ _2939_ _2810_ _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_227_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_2726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Left_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8604__A1 _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8962_ net181 core_0.decode.i_imm_pass\[13\] _1263_ _4449_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8080__A2 _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6091__A1 core_0.execute.rf.reg_outputs\[10\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_223_3192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7913_ _3650_ _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6091__B2 core_0.execute.rf.reg_outputs\[11\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8893_ core_0.execute.pc_high_buff_out\[6\] _4385_ _1430_ _4408_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_210_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8907__A2 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4641__A2 net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7844_ core_0.execute.rf.reg_outputs\[8\]\[3\] _3607_ _3609_ _3612_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_i_clk clknet_4_8__leaf_i_clk clknet_leaf_30_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_195_2855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7775_ _3435_ _3563_ _3572_ _0336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4987_ core_0.fetch.prev_request_pc\[14\] _1155_ _1166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6394__A2 _2366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7591__B2 net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9514_ _0524_ clknet_leaf_41_i_clk core_0.execute.next_ready_delayed vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6726_ _2655_ _2661_ _2662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_190_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer41_I net268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7991__B _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_45_i_clk clknet_4_10__leaf_i_clk clknet_leaf_45_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_9445_ _0455_ clknet_leaf_145_i_clk core_0.execute.rf.reg_outputs\[3\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6146__A2 _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6657_ _1829_ _1858_ _1862_ _2599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__5067__I _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7343__A1 net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7483__S _3366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5608_ _1591_ _1573_ _1639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9376_ _0386_ clknet_leaf_39_i_clk core_0.execute.rf.reg_outputs\[7\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7894__A2 _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6588_ _2522_ _2529_ _2530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8327_ _1679_ _1539_ _2344_ _3942_ _3943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_239_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5539_ core_0.fetch.prev_request_pc\[2\] _1595_ _1084_ net168 _1599_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8258_ _3835_ _3836_ _3879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9258__CLK clknet_leaf_1_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7209_ _2459_ _2463_ _2532_ _3133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8189_ _1674_ _1831_ _1837_ _2372_ _2140_ _3815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_245_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5409__A1 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8071__A2 _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A1 _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7582__A1 _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput17 i_disable net17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6137__A2 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput28 i_mem_data[1] net28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput39 i_req_data[10] net39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_220_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5345__B1 _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7885__A2 _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__A1 core_0.decode.oc_alu_mode\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4699__A2 net296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6310__B _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5360__A3 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8834__A1 _4324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7637__A2 _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__A1 _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A1 core_0.execute.rf.reg_outputs\[15\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7270__B1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__B2 core_0.execute.rf.reg_outputs\[1\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4623__A2 net324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4910_ _1088_ _1016_ _1089_ _1090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5890_ core_0.decode.oc_alu_mode\[6\] _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_87_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4841_ core_0.fetch.out_buffer_valid _1021_ _1022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7573__A1 _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6376__A2 _2349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ net26 _1347_ _3437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4772_ core_0.dec_l_reg_sel\[1\] _0953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_23_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6511_ _1745_ _2040_ _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7491_ core_0.dec_rf_ie\[14\] core_0.ew_reg_ie\[14\] _2421_ _3379_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7325__A1 _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8700__B _1723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9230_ _0241_ clknet_leaf_142_i_clk core_0.ew_reg_ie\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_141_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6442_ net86 _2403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_132_2102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7876__A2 _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_2796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5887__A1 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9161_ _0172_ clknet_leaf_75_i_clk core_0.execute.mem_stage_pc\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6373_ net96 _2347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__9400__CLK clknet_leaf_145_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8112_ _3427_ _3759_ _3766_ _0479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8825__A1 core_0.execute.pc_high_buff_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5324_ core_0.decode.i_instr_l\[3\] core_0.decode.i_instr_l\[2\] _1273_ _1442_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7628__A2 _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9092_ _0117_ clknet_leaf_95_i_clk core_0.decode.i_imm_pass\[13\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5639__A1 _1026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6836__B1 _2768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8043_ _3446_ _3715_ _3726_ _0450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_54_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5255_ core_0.dec_jump_cond_code\[1\] _1376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_225_3210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5186_ _1330_ _1332_ _0002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4862__A2 net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8053__A2 _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_2231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_rebuffer89_I _1796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6064__A1 net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6064__B2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7800__A2 _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8945_ _4440_ _0638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5811__A1 _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4614__A2 _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8876_ net201 _4387_ _4394_ _4395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7013__B1 _2433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7827_ _3463_ _3586_ _3601_ _0359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6367__A2 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_175_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_236_3350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7758_ _3473_ _3543_ _3561_ _0330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_191_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _2636_ _2640_ _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7316__A1 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7689_ core_0.execute.rf.reg_outputs\[12\]\[1\] _3521_ _3513_ _3523_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_123_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9428_ _0438_ clknet_leaf_14_i_clk core_0.execute.rf.reg_outputs\[4\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_117_1919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_2360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7867__A2 _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9359_ _0369_ clknet_leaf_29_i_clk core_0.execute.rf.reg_outputs\[8\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6130__B _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8816__A1 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__B1 _2758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6842__A3 _2687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8057__B _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8044__A2 _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_1_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6055__A1 core_0.execute.rf.reg_outputs\[13\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_154_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A2 net309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7555__A1 _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6358__A2 _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_166_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5566__B1 _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7858__A2 _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_79_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4541__B2 core_0.execute.rf.reg_outputs\[1\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_168_2529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8283__A2 _2487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7650__I _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6294__A1 _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ _1033_ _1146_ _1164_ _1210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_224_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_225_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__B2 core_0.execute.rf.reg_outputs\[10\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_195_Right_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6991_ core_0.execute.alu_mul_div.div_res\[4\] _2921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_220_3151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7794__A1 _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8730_ core_0.execute.sreg_jtr_buff.o_d\[1\] _4217_ _4283_ _4285_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5942_ core_0.execute.rf.reg_outputs\[13\]\[10\] _1792_ _1815_ core_0.execute.rf.reg_outputs\[9\]\[10\]
+ _1932_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_220_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_2658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8661_ net81 _1699_ _1709_ _4205_ _4229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_75_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5873_ _1769_ _1829_ _1858_ _1862_ _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_75_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7612_ _3402_ _3476_ _3478_ _0267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_192_2814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4824_ core_0.dec_wfi core_0.execute.alu_mul_div.comp _1001_ _1004_ _1005_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_185_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8592_ core_0.execute.alu_flag_reg.o_d\[0\] _4167_ _1431_ _4170_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7543_ core_0.execute.rf.reg_outputs\[15\]\[3\] _3403_ _3422_ _3423_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4755_ core_0.ew_reg_ie\[14\] _0928_ _0663_ _0936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4780__A1 core_0.ew_reg_ie\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7474_ _3370_ _0237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7849__A2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4780__B2 core_0.ew_reg_ie\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4686_ _0870_ net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_126_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9213_ _0224_ clknet_leaf_77_i_clk net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_160_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_231_3280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6425_ _2391_ _2385_ _2392_ _0166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9144_ _0156_ clknet_leaf_98_i_clk core_0.execute.alu_mul_div.div_cur\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6356_ _2325_ _2330_ _2141_ _2331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5307_ net105 _1416_ _1427_ _0922_ _1428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_9075_ _0100_ clknet_leaf_101_i_clk core_0.decode.i_instr_l\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6287_ _2246_ _2269_ _2270_ _2217_ _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5088__A2 core_0.decode.i_instr_l\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8026_ core_0.execute.rf.reg_outputs\[3\]\[0\] _3716_ _3704_ _3717_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5238_ _1364_ net143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_215_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input31_I i_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6824__A3 _2756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8026__A2 _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5169_ _1230_ _1316_ _1289_ _1318_ _0000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6037__A1 net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7234__B1 _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_205_2968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7785__A1 _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_162_Right_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8982__B1 _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output118_I net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4599__A1 core_0.execute.rf.reg_outputs\[10\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8928_ core_0.dec_used_operands\[1\] _1495_ _4431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_211_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5260__A2 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7537__A1 net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8859_ _4328_ _4380_ _4381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9446__CLK clknet_leaf_145_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_10_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4771__A1 core_0.ew_reg_ie\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5315__A3 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_80_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5720__B1 _1717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_3449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_218_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6086__I _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8017__A2 _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A1 core_0.execute.rf.reg_outputs\[14\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__B1 _3142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7776__A1 core_0.execute.rf.reg_outputs\[10\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__A2 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5539__B1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5003__A2 _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6751__A2 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_2599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4540_ core_0.execute.rf.reg_outputs\[14\]\[13\] _0686_ _0700_ core_0.execute.rf.reg_outputs\[12\]\[13\]
+ _0736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ _0660_ _0663_ _0668_ _0664_ _0669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_111_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6503__A2 _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7700__A1 _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6210_ _2157_ _2196_ _2197_ _2198_ _2199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_229_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5711__B1 _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7190_ _1292_ _3100_ _3111_ _3114_ _3115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6141_ _1419_ _2131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_209_3024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6267__A1 _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ core_0.execute.rf.reg_outputs\[10\]\[6\] net226 _2062_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4817__A2 _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ _1195_ _1046_ _1158_ _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8008__A2 _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_205_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7767__A1 _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_221_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _2902_ _2495_ _2904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_221_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5242__A2 core_0.ew_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8713_ _4212_ core_0.execute.mem_stage_pc\[13\] _4202_ _4271_ _4272_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_76_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ _1771_ _1913_ _1914_ _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_48_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6990__A2 _2918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8644_ _4203_ _4042_ _4213_ _4214_ _1661_ _4215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5856_ net314 net208 _1845_ _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_152_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8192__A1 _1674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8192__B2 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4807_ core_0.ew_reg_ie\[7\] _0948_ _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8575_ _4053_ _4152_ _4153_ _1702_ _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_28_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5787_ core_0.execute.rf.reg_outputs\[4\]\[0\] _1776_ _1777_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_2163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6742__A2 net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7526_ _3382_ core_0.ew_data\[1\] _3407_ _3408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__4753__A1 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4738_ core_0.execute.prev_pc_high\[5\] _0917_ _0918_ _0919_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_102_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_2330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7457_ _3361_ _0229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4669_ core_0.execute.rf.reg_outputs\[4\]\[3\] net318 net284 core_0.execute.rf.reg_outputs\[13\]\[3\]
+ _0855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5075__I core_0.decode.i_instr_l\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7491__S _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6408_ _1714_ _2380_ _0161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7388_ _2672_ _3307_ _3308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5848__A4 _1837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_231_Right_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_9127_ _0139_ clknet_leaf_70_i_clk core_0.execute.sreg_priv_control.o_d\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6339_ _2219_ _2315_ _2316_ _0156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6258__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_9058_ _0084_ clknet_leaf_89_i_clk core_0.fetch.prev_request_pc\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_73_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4808__A2 _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8009_ core_0.execute.rf.reg_outputs\[4\]\[9\] _3700_ _3704_ _3707_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_215_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_212_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7758__A1 _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_27_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8183__A1 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8070__B _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7930__A1 _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5941__B1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6497__A1 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8238__A2 _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6249__A1 core_0.execute.alu_mul_div.div_cur\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcore0_228 o_mem_addr_high[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_206_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4680__B1 net341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8960__S _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_207_Left_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4492__C _0689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_2628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5710_ net251 _1704_ _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4983__A1 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6690_ core_0.execute.rf.reg_outputs\[7\]\[2\] _2611_ _2612_ core_0.execute.rf.reg_outputs\[5\]\[2\]
+ _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_17_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8174__A1 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4999__I _1020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5641_ _1656_ _0118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7921__A1 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8360_ _3958_ _3967_ _3973_ _3974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5572_ _1241_ _1616_ _1617_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7311_ _3201_ _3232_ _3233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_215_3094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5109__B _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4523_ _0719_ _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
X_8291_ _3901_ _3909_ _3802_ _3910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_216_Left_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_170_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__A1 _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7242_ _2708_ net307 _3166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_229_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5160__A1 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7173_ _3098_ _0208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8229__A2 core_0.execute.alu_mul_div.cbit\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_2757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_238_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6124_ _2110_ _2111_ _2112_ _2113_ _2114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_237_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6055_ core_0.execute.rf.reg_outputs\[13\]\[7\] _1791_ net333 core_0.execute.rf.reg_outputs\[4\]\[7\]
+ _2045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5999__B1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5006_ core_0.fetch.prev_request_pc\[11\] _1152_ _1182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_198_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5463__A2 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4683__B _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8155__B _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_225_Left_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_rebuffer71_I net298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_202_2938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5215__A2 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6412__A1 core_0.execute.sreg_data_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7460__I0 net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6957_ _2839_ _2886_ _2887_ _0203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_198_2886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4974__A1 core_0.fetch.prev_request_pc\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5908_ _1897_ _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_9_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6888_ _2819_ _1314_ core_0.execute.alu_mul_div.i_mod _2820_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8165__A1 net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8627_ _4198_ _1696_ _1702_ _4199_ _0561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5839_ _1828_ _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XANTENNA__6403__B _2217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6715__A2 _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8960__I0 net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A1 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8558_ _4138_ _4139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_20_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_234_Left_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_161_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output185_I net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7509_ core_0.ew_reg_ie\[12\] core_0.ew_reg_ie\[13\] core_0.ew_reg_ie\[14\] core_0.ew_reg_ie\[15\]
+ _3392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_161_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8489_ net82 _1738_ _4078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_75_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5533__I _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_229_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_242_3419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8640__A2 _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_243_Left_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_204_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_2429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6364__I net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6403__A1 _2206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6954__A2 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8156__A1 _3446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6706__A2 _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9164__CLK clknet_leaf_92_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5914__B1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5914__C2 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_171_2569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5142__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5443__I core_0.execute.alu_mul_div.cbit\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9062__D core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__A3 _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6983__B core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_219_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6642__A1 _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_2698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4653__B1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7860_ _3457_ _3607_ _3620_ _0373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8395__A1 _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6811_ _2075_ _2736_ _2743_ _2744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7791_ core_0.execute.rf.reg_outputs\[10\]\[13\] _3570_ _3580_ _3581_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6945__A2 _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9530_ _0540_ clknet_leaf_120_i_clk core_0.execute.alu_mul_div.div_res\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6742_ net184 net177 _1421_ _2676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_217_3112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8147__A1 _3420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9507__CLK clknet_leaf_122_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9461_ _0471_ clknet_leaf_137_i_clk core_0.execute.rf.reg_outputs\[2\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6673_ _2607_ _2614_ _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__9237__D _0248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5624_ core_0.decode.i_imm_pass\[6\] _1645_ _1648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8412_ _4015_ _4018_ _4019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9392_ _0402_ clknet_leaf_33_i_clk core_0.execute.rf.reg_outputs\[6\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_135_2133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8343_ core_0.execute.alu_mul_div.mul_res\[11\] _3957_ _3958_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5555_ core_0.fetch.prev_request_pc\[10\] _1082_ _1083_ net161 _1607_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_41_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6877__C _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4506_ _0661_ _0662_ core_0.dec_r_reg_sel\[1\] _0675_ _0704_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_8274_ _1535_ _2353_ _3894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5486_ _1567_ _1551_ _1568_ _0051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7122__A2 core_0.execute.sreg_irq_pc.o_d\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7225_ _2804_ _3069_ _3142_ _1768_ _3148_ _3149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__5133__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_228_3252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6881__A1 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6881__B2 _1865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7156_ _1743_ _3081_ core_0.execute.alu_mul_div.i_div _3082_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7989__B _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Left_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_238_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6107_ core_0.execute.rf.reg_outputs\[2\]\[2\] _1797_ _1815_ core_0.execute.rf.reg_outputs\[9\]\[2\]
+ _2097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_70_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8622__A2 _4194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7087_ _2430_ _2974_ _3014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6633__A1 _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5436__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6038_ core_0.execute.rf.reg_outputs\[8\]\[5\] net345 net332 core_0.execute.rf.reg_outputs\[4\]\[5\]
+ _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_197_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4644__B1 net318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer40 net206 net268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8386__A1 _2370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer51 net205 net279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_68_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer62 _0684_ net290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_240_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__C _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer73 core_0.dec_l_reg_sel\[1\] net328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_139_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer84 _0672_ net312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6936__A2 _2859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7989_ core_0.execute.rf.reg_outputs\[4\]\[0\] _3695_ _3689_ _3696_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer95 _1841_ net342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA_output100_I net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4947__A1 core_0.fetch.prev_request_pc\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_239_3381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5528__I _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_2391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7113__A2 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5124__A1 core_0.decode.i_instr_l\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8861__A2 _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5675__A2 _1680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4478__A3 core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7899__B _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8613__A2 _3150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6624__A1 _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A2 _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7411__C _3329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8377__A1 _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8129__A1 _3462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_99_1703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5363__A1 core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_212_3053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_149_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5340_ _1294_ _1298_ _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput105 net105 o_c_instr_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_149_Left_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput116 net116 o_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput127 net127 o_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput138 net138 o_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput149 net149 o_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5271_ core_0.dec_jump_cond_code\[3\] _1391_ _1392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8852__A2 _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7010_ _2009_ _2719_ _2939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_184_2716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7602__B _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8604__A2 _3311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6615__A1 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5418__A2 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8961_ _4448_ _0646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_1810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4626__B1 _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4517__I net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_223_3193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7912_ _3650_ _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_222_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8892_ net280 _4387_ _4406_ _4407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8368__A1 _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7843_ _3415_ _3606_ _3611_ _0365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8433__B _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4986_ _1164_ _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7774_ core_0.execute.rf.reg_outputs\[10\]\[5\] _3570_ _3568_ _3572_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_195_2856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7591__A2 core_0.ew_data\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9513_ _0523_ clknet_leaf_122_i_clk core_0.execute.alu_mul_div.mul_res\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6725_ _2627_ _2654_ _2661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5348__I core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6656_ _1883_ _1864_ _2595_ _2597_ _2598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_9444_ _0454_ clknet_leaf_13_i_clk core_0.execute.rf.reg_outputs\[3\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_rebuffer34_I _1848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7343__A2 _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8540__A1 _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6888__B core_0.execute.alu_mul_div.i_mod vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5607_ core_0.decode.i_instr_l\[14\] _1616_ _1638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5354__A1 _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9375_ _0385_ clknet_leaf_40_i_clk core_0.execute.rf.reg_outputs\[7\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_5_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6587_ _2456_ _2525_ _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_59_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _1597_ _1598_ _0073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8326_ _1538_ _2364_ _3941_ _1679_ _3942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_input61_I i_req_data[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6400__C _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8257_ _1669_ _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_100_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _1550_ _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__8843__A2 _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5083__I _1239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7208_ _3132_ _0209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6854__A1 core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5657__A2 _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5016__C _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8188_ _1543_ _2143_ _3813_ _1545_ _3814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7139_ _2500_ _2515_ _2519_ _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5409__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4617__B1 net312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8359__A1 core_0.execute.alu_mul_div.mul_res\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6909__A2 _2740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7031__A1 _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_2420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7582__A2 _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput18 i_irq net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8531__A1 _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput29 i_mem_data[2] net29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5345__B2 _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_150_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__A2 core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7098__A1 _2054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7098__B2 net287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__A2 _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6845__A1 _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_176_Right_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_236_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_229_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8598__A1 _3330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_205_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_232_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7270__A1 core_0.execute.sreg_priv_control.o_d\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__A2 _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7270__B2 net3 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_232_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_220_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_75_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7022__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4840_ core_0.fetch.out_buffer_data_instr\[31\] _1021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_75_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7573__A2 _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8770__A1 core_0.execute.sreg_scratch.o_d\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4771_ core_0.ew_reg_ie\[9\] _0950_ _0951_ _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6510_ _1749_ net218 _2452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7490_ _3378_ _0245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8522__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6441_ _2401_ _2385_ _2402_ _0172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5336__A1 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_157_Left_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_2797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9160_ _0171_ clknet_leaf_75_i_clk core_0.execute.mem_stage_pc\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6372_ _1541_ net214 _2345_ _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8111_ core_0.execute.rf.reg_outputs\[1\]\[4\] _3765_ _3756_ _3766_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7089__A1 _2439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5323_ _1439_ core_0.decode.i_instr_l\[8\] _1440_ _1441_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_100_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9091_ _0116_ clknet_leaf_95_i_clk core_0.decode.i_imm_pass\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_228_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8825__A2 _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8042_ core_0.execute.rf.reg_outputs\[3\]\[7\] _3722_ _3718_ _3726_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5639__A2 _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6836__A1 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5254_ _1374_ core_0.execute.alu_flag_reg.o_d\[0\] _1375_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_114_1880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6836__B2 core_0.execute.sreg_scratch.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_143_Right_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_227_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_225_3211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_112_i_clk clknet_4_6__leaf_i_clk clknet_leaf_112_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_139_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5185_ _0038_ _1247_ _1331_ _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_EDGE_ROW_166_Left_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_208_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7261__A1 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6064__A2 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8944_ net187 core_0.decode.i_imm_pass\[4\] _1264_ _4440_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_155_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_127_i_clk clknet_4_4__leaf_i_clk clknet_leaf_127_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5811__A2 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8875_ _0904_ _4383_ _4394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8163__B _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7013__A1 _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8210__B1 _1783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7013__B2 core_0.decode.oc_alu_mode\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7826_ core_0.execute.rf.reg_outputs\[9\]\[12\] _3591_ _3595_ _3601_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8761__A1 core_0.execute.sreg_scratch.o_d\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_236_3340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5575__A1 _1143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _1105_ _1109_ _1147_ _1148_ _1149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7757_ core_0.execute.rf.reg_outputs\[11\]\[15\] _3541_ _3554_ _3561_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6708_ _2644_ _2645_ _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_191_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_175_Left_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_191_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7316__A2 net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7688_ _3402_ _3520_ _3522_ _0299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8389__I core_0.execute.alu_mul_div.mul_res\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__A1 _1239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9427_ _0437_ clknet_leaf_16_i_clk core_0.execute.rf.reg_outputs\[4\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _1769_ _2580_ net267 _2581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_117_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_2361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9358_ _0368_ clknet_leaf_27_i_clk core_0.execute.rf.reg_outputs\[8\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8309_ core_0.execute.alu_mul_div.mul_res\[8\] _3918_ _3926_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_219_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8816__A2 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4550__A2 _0680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9289_ _0299_ clknet_leaf_5_i_clk core_0.execute.rf.reg_outputs\[12\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_219_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__A1 _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6827__B2 _2759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_110_Right_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_245_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_184_Left_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_245_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_165_2490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6055__A2 _1791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8073__B _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_91_i_clk clknet_4_15__leaf_i_clk clknet_leaf_91_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8752__A1 core_0.execute.sreg_scratch.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5566__A1 core_0.fetch.prev_request_pc\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_193_Left_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5566__B2 net166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6763__B1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8504__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_245_Right_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4541__A2 _0673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6818__A1 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_236_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_224_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_44_i_clk clknet_4_10__leaf_i_clk clknet_leaf_44_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7243__A1 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6046__A2 net336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6990_ _2124_ _2918_ _2919_ _0996_ _2920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__7794__A2 _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_220_3152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_232_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5941_ core_0.execute.rf.reg_outputs\[8\]\[10\] _1794_ _1776_ core_0.execute.rf.reg_outputs\[4\]\[10\]
+ _1931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_220_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_2659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8660_ core_0.execute.sreg_irq_pc.o_d\[4\] _4210_ _4228_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5872_ _1859_ _1860_ _1861_ _1862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_34_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8743__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _1002_ net20 _1003_ _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_29_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7611_ core_0.execute.rf.reg_outputs\[14\]\[0\] _3477_ _3467_ _3478_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_192_2815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9248__CLK clknet_leaf_37_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8711__B _1727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8591_ _4154_ _4164_ _4168_ _4169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7542_ _1430_ _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_16_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4754_ _0929_ _0932_ _0933_ _0934_ _0935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_133_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_212_Right_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5309__A1 _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7473_ core_0.dec_rf_ie\[5\] core_0.ew_reg_ie\[5\] _3366_ _3370_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4685_ net95 net323 _0864_ _0869_ _0870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_43_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9212_ _0223_ clknet_leaf_77_i_clk net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6424_ core_0.execute.mem_stage_pc\[2\] _2386_ _2387_ _2392_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_231_3281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9143_ _0155_ clknet_leaf_98_i_clk core_0.execute.alu_mul_div.div_cur\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6355_ _2147_ _2329_ _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4532__A2 _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6809__A1 _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5306_ net105 _1426_ _1427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9074_ _0099_ clknet_leaf_106_i_clk core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6286_ core_0.execute.alu_mul_div.div_cur\[5\] _2224_ _2270_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_227_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5237_ core_0.ew_data\[6\] core_0.ew_data\[14\] _1349_ _1364_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8025_ _3714_ _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_215_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_242_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5168_ _1317_ _1250_ _1318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input24_I i_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7489__S _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6037__A2 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7234__B2 core_0.execute.sreg_scratch.o_d\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5099_ core_0.decode.i_instr_l\[6\] _1238_ core_0.decode.i_instr_l\[5\] _1255_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_67_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_205_2969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7785__A2 _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8982__B2 _1476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8927_ _1494_ _4423_ _4430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5796__A1 _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4599__A2 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6993__B1 _2920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8858_ core_0.execute.pc_high_buff_out\[7\] _4329_ _4379_ _4380_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5548__A1 _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7809_ core_0.execute.rf.reg_outputs\[9\]\[4\] _3591_ _3580_ _3592_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8789_ core_0.execute.sreg_irq_flags.o_d\[3\] _4217_ _4320_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4756__C1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4771__A2 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__I _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output92_I net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_23_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6512__A3 _2453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5720__A1 core_0.execute.sreg_priv_control.o_d\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5472__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__B2 _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8068__B _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7225__A1 _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__A2 _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8582__I _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7225__B2 _1768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7776__A2 _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8973__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6316__B _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7528__A2 _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5539__A1 core_0.fetch.prev_request_pc\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5539__B2 net168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6751__A3 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8958__S _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__I core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4470_ core_0.dec_r_reg_sel\[1\] _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_52_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7700__A2 _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5711__B2 _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6140_ _1317_ _2127_ _2129_ _2130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_209_3025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_51_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ core_0.execute.rf.reg_outputs\[2\]\[6\] net336 _2061_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5181__I _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5022_ core_0.fetch.prev_request_pc\[8\] _1150_ _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_127_2035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7767__A2 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6973_ _2902_ _2495_ _2903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8712_ _4224_ _4135_ _4270_ _1662_ _4271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_178_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ core_0.execute.rf.reg_outputs\[13\]\[8\] _1791_ net333 core_0.execute.rf.reg_outputs\[4\]\[8\]
+ _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8716__A1 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8643_ _1705_ _4214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _1518_ net192 _1845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__7836__I _3605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8192__A2 net306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_233_3310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4806_ _0985_ _0986_ _0942_ _0947_ _0987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8574_ net77 _4052_ _4153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_173_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5786_ _1775_ _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_118_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7525_ _3381_ _3405_ _3406_ _3407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4737_ core_0.execute.prev_pc_high\[4\] _0912_ _0918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4753__A2 _0928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5950__A1 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5356__I core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_2320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7456_ net118 _3261_ _2415_ _3361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4668_ core_0.execute.rf.reg_outputs\[5\]\[3\] _0677_ _0703_ core_0.execute.rf.reg_outputs\[15\]\[3\]
+ _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_102_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6407_ _0926_ _1371_ _2380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5702__A1 core_0.execute.sreg_data_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7387_ _2703_ _3297_ _3304_ _3306_ _3307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7571__I _3446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4599_ core_0.execute.rf.reg_outputs\[10\]\[8\] net221 net220 core_0.execute.rf.reg_outputs\[9\]\[8\]
+ _0790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5702__B2 _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9126_ _0138_ clknet_leaf_108_i_clk core_0.execute.sreg_priv_control.o_d\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6338_ core_0.execute.alu_mul_div.div_cur\[12\] _2218_ _0999_ _2316_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6258__A2 _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9057_ _0083_ clknet_leaf_86_i_clk core_0.fetch.prev_request_pc\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_73_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6269_ _2141_ _2215_ _2255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_215_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8008_ _3450_ _3694_ _3706_ _0435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_231_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_2460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7758__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__A1 _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6430__A2 _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8707__A1 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5467__S _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7930__A2 _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4744__A2 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6497__A2 _2054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_112_Left_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7694__A1 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6249__A2 _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_237_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_13_Right_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_173_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7749__A2 _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4680__B2 core_0.execute.rf.reg_outputs\[3\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Left_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6421__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_176_2629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5640_ _1016_ core_0.decode.i_imm_pass\[14\] _1368_ _1656_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7921__A2 _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Right_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5571_ _1368_ _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4735__A2 _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7310_ _1684_ core_0.execute.sreg_irq_pc.o_d\[12\] _3231_ _3232_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_26_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ net293 _0663_ _0688_ _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XPHY_EDGE_ROW_130_Left_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_143_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_215_3095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ core_0.execute.alu_mul_div.mul_res\[7\] _3908_ _3909_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_40_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7241_ _2711_ _3155_ _3162_ _3164_ _3165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_151_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5904__I net325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7172_ core_0.ew_data\[8\] _3097_ _0199_ _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7324__C _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5160__A2 _1309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_2758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7437__A1 _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6123_ core_0.execute.rf.reg_outputs\[13\]\[1\] _1792_ _1804_ core_0.execute.rf.reg_outputs\[11\]\[1\]
+ _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6054_ core_0.execute.rf.reg_outputs\[8\]\[7\] net346 _2044_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_225_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Right_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_147_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5999__B2 core_0.execute.rf.reg_outputs\[4\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5005_ _1057_ _1181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_225_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8937__A1 _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4671__A1 core_0.execute.rf.reg_outputs\[11\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9586__CLK clknet_leaf_110_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_202_2939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6412__A2 _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7460__I1 _3335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6956_ core_0.ew_data\[3\] _2642_ _2887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_198_2887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5907_ _1859_ net256 _1861_ _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_48_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6887_ core_0.execute.alu_mul_div.div_res\[2\] _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_120_1949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8165__A2 _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6470__I _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8626_ _1696_ _4055_ _4199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_40_Right_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5838_ net93 _1813_ _1817_ _1827_ _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_64_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4726__A2 net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8557_ _1736_ _4135_ _4136_ _4137_ _4138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_173_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_161_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5769_ _1518_ net217 _1758_ _1759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_20_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7508_ core_0.ew_reg_ie\[8\] core_0.ew_reg_ie\[9\] core_0.ew_reg_ie\[10\] core_0.ew_reg_ie\[11\]
+ _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_115_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8488_ _1206_ _4076_ _4077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_32_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output178_I net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7439_ _2616_ _2923_ _3352_ _0220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5814__I _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9109_ _0012_ clknet_leaf_112_i_clk core_0.decode.oc_alu_mode\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_216_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6100__A1 net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7600__B2 net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_223_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8156__A2 _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6380__I _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9309__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7903__A2 _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5914__A1 core_0.execute.rf.reg_outputs\[9\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_2559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7116__B1 _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7667__A1 _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8100__I _3758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5142__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4496__A4 _0664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_2699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8919__A1 _1488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4653__A1 core_0.execute.rf.reg_outputs\[10\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_145_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6810_ _2011_ _1898_ _2742_ _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7790_ _3512_ _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_202_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6741_ core_0.execute.sreg_irq_pc.o_d\[0\] _2675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_217_3113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6504__B _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8147__A2 _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9460_ _0470_ clknet_leaf_14_i_clk core_0.execute.rf.reg_outputs\[2\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6158__A1 core_0.execute.alu_mul_div.div_cur\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6672_ _2610_ _2613_ _2614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8411_ _2140_ _2354_ _1545_ _4018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_128_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5623_ _1034_ _1615_ _1647_ _0109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9391_ _0401_ clknet_leaf_33_i_clk core_0.execute.rf.reg_outputs\[6\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_135_2134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8342_ _1536_ _3855_ _3956_ _3957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5554_ _1597_ _1606_ _0081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7658__A1 core_0.execute.rf.reg_outputs\[13\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4505_ _0702_ _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5485_ net40 _1554_ _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8273_ _3877_ _3888_ _3892_ _3893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_41_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7224_ _1338_ _3143_ _2464_ core_0.decode.oc_alu_mode\[6\] _3147_ _3148_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_111_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6330__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_228_3253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7155_ core_0.execute.alu_mul_div.mul_res\[8\] _3081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_226_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6106_ _2092_ _2093_ _2094_ _2095_ _2096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_70_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8083__A1 _3450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7086_ _2489_ _3011_ _3012_ _3013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_241_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7830__A1 core_0.execute.rf.reg_outputs\[9\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6633__A2 _2574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6037_ net98 _1771_ _2027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_146_2263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4644__A1 core_0.execute.rf.reg_outputs\[5\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_241_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer30 _1843_ net258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer41 net268 net269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_240_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8386__A2 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer52 net279 net280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer63 _0684_ net291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_139_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer74 core_0.dec_l_reg_sel\[1\] net329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_7988_ _3693_ _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_25_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer85 net331 net332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_194_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer96 _1748_ net343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4947__A2 _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6939_ _1290_ _2868_ _2869_ _1742_ _2870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_95_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_3382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5809__I _1798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4713__I _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8609_ _1431_ _4182_ _4183_ _4184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_174_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9589_ _0599_ clknet_leaf_108_i_clk core_0.execute.sreg_scratch.o_d\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_2392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_157_Right_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7649__A1 _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__B1 _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5124__A2 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4478__A4 _0675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5480__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4883__A1 _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8074__A1 _3427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8076__B _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7821__A1 _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_15__f_i_clk clknet_3_7_0_i_clk clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_231_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5832__B1 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_232_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6388__A1 _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8129__A2 _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7888__A1 _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6978__C core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5363__A2 _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_124_Right_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_212_3054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput106 net106 o_icache_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8966__S _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput117 net117 o_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput128 net128 o_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_71_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput139 net139 o_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5270_ _1377_ _1390_ core_0.dec_jump_cond_code\[2\] _1391_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8999__CLK clknet_leaf_133_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_2717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8065__A1 _3401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__B1 _1787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6615__A2 _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7812__A1 _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8960_ net180 core_0.decode.i_imm_pass\[12\] _1263_ _4448_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4626__A1 core_0.execute.rf.reg_outputs\[5\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7911_ core_0.ew_reg_ie\[6\] _3395_ _3650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_223_3183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_223_3194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8891_ _0914_ _4383_ _4406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8714__B _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8368__A2 _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7842_ core_0.execute.rf.reg_outputs\[8\]\[2\] _3607_ _3609_ _3611_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7773_ _3428_ _3563_ _3571_ _0335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4985_ core_0.fetch.pc_flush_override core_0.decode.i_flush _1164_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XANTENNA__5051__A1 core_0.fetch.prev_request_pc\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_195_2857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4533__I _0729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9512_ _0522_ clknet_leaf_119_i_clk core_0.execute.alu_mul_div.mul_res\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6724_ _2658_ _2659_ _2660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_175_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9443_ _0453_ clknet_leaf_45_i_clk core_0.execute.rf.reg_outputs\[3\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7879__A1 core_0.execute.rf.reg_outputs\[7\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6655_ _1329_ _1988_ _2596_ _1883_ _2597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_128_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6000__B1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5606_ _1635_ _1637_ _0102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9374_ _0384_ clknet_leaf_40_i_clk core_0.execute.rf.reg_outputs\[7\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_30_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6586_ _2500_ _2515_ _2519_ _2527_ _2528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA_rebuffer27_I net254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7065__B _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8325_ _1538_ _2352_ _3941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4562__B1 _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5537_ core_0.fetch.prev_request_pc\[1\] _1595_ _1084_ net167 _1598_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_169_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8256_ _3865_ _3870_ _3876_ _3877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5468_ _1558_ _0043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input54_I i_req_data[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9004__CLK clknet_leaf_133_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_245_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7207_ core_0.ew_data\[9\] _3131_ _0199_ _3132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_218_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8187_ _1543_ _2146_ _3813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4865__A1 _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5399_ _1247_ _1442_ _1339_ _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8056__A1 _3465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7138_ _3061_ _3062_ _3063_ _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_226_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_214_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4708__I _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6606__A2 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7803__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ net13 _2996_ _2768_ core_0.execute.sreg_scratch.o_d\[6\] _2689_ _2997_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_213_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5290__A1 _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_226_Right_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6909__A3 _2737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_159_2421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6790__A1 _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 i_mc_core_int net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5345__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4553__B1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5896__A3 core_0.decode.oc_alu_mode\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_229_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__A3 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6845__A2 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7703__B _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4856__A1 _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8047__A1 _3453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6058__B1 _1778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_205_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5805__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_232_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7270__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_18_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7022__A2 core_0.execute.alu_mul_div.mul_res\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5033__A1 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5449__I core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8770__A2 _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6781__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ core_0.dec_l_reg_sel\[3\] core_0.dec_l_reg_sel\[2\] _0951_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_173_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4792__C2 core_0.ew_reg_ie\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6440_ core_0.execute.mem_stage_pc\[8\] _2395_ _2387_ _2402_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5336__A2 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_2787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_2798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6371_ _1541_ _2040_ _2345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8110_ _3758_ _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_140_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8286__A1 _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5322_ core_0.decode.i_instr_l\[7\] _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_2_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9090_ _0115_ clknet_leaf_96_i_clk core_0.decode.i_imm_pass\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8709__B _4201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8041_ _3440_ _3715_ _3725_ _0449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_228_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7613__B _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6836__A2 _1411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5253_ core_0.dec_jump_cond_code\[0\] _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4847__A1 _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8038__A1 core_0.execute.rf.reg_outputs\[3\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_225_3212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5184_ _1234_ _1258_ _1243_ _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_236_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_2233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7261__A2 _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8943_ _1687_ _0038_ _4439_ _0637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7839__I _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5811__A3 _1790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8874_ _4386_ _4392_ _4393_ _0614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_195_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8210__A1 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7825_ _3460_ _3586_ _3600_ _0358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8210__B2 _1810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5024__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8761__A2 _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_236_3341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7756_ _3470_ _3543_ _3560_ _0329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6772__A1 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4968_ core_0.fetch.prev_request_pc\[2\] core_0.fetch.prev_request_pc\[1\] core_0.fetch.prev_request_pc\[0\]
+ _1148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_93_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6707_ core_0.execute.rf.reg_outputs\[7\]\[4\] _2611_ _2612_ core_0.execute.rf.reg_outputs\[5\]\[4\]
+ _2645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_191_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7687_ core_0.execute.rf.reg_outputs\[12\]\[0\] _3521_ _3513_ _3522_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4899_ core_0.fetch.pc_reset_override _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_163_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9426_ _0436_ clknet_leaf_22_i_clk core_0.execute.rf.reg_outputs\[4\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_190_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6638_ _2103_ _2116_ _2580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5327__A2 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_2362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4535__B1 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5308__B _1428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9357_ _0367_ clknet_leaf_29_i_clk core_0.execute.rf.reg_outputs\[8\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5094__I _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6569_ _2508_ _2509_ _2510_ _2511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8308_ _3081_ _3863_ _3925_ _0516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8277__A1 _3893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9288_ _0298_ clknet_leaf_153_i_clk core_0.execute.rf.reg_outputs\[13\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output160_I net160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8239_ _3832_ _3860_ _3861_ _0511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5822__I _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4838__A1 _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8029__A1 core_0.execute.rf.reg_outputs\[3\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_165_2491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5799__C1 _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8201__A1 _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Right_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8752__A2 _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5566__A2 _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6763__B2 _2694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8504__A2 net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6515__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_78_Right_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6818__A2 _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4829__A1 _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_220_3153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5940_ _1929_ _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_220_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_87_Right_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5871_ net212 _1855_ _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_87_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5006__A1 core_0.fetch.prev_request_pc\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7610_ _3475_ _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__8743__A2 _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4822_ core_0.ew_mem_access core_0.ew_submit _1003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8590_ _0890_ _4165_ _4167_ _4168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6754__A1 core_0.execute.pc_high_buff_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_192_2816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8711__C _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7541_ _3420_ _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_141_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4753_ core_0.ew_reg_ie\[2\] _0928_ _0931_ core_0.ew_reg_ie\[3\] _0930_ core_0.ew_reg_ie\[1\]
+ _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_83_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7472_ _3369_ _0236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6506__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4684_ _0865_ _0866_ _0867_ _0868_ _0869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_71_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6357__I1 _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9211_ _0222_ clknet_leaf_54_i_clk net126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6423_ net79 _2391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_231_3282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_96_Right_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8259__A1 _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9142_ _0154_ clknet_leaf_98_i_clk core_0.execute.alu_mul_div.div_cur\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6354_ _2144_ _2324_ _2194_ _2329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6738__I core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ _1397_ _1418_ _1422_ _1425_ _1426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_9073_ _0098_ clknet_leaf_128_i_clk core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_11_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6285_ _2261_ _2268_ _2141_ _2269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_227_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8024_ _3714_ _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5236_ _1363_ net142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6690__B1 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ core_0.execute.alu_mul_div.i_mod _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_208_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7234__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8431__A1 _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5098_ core_0.decode.oc_alu_mode\[6\] _1254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__5245__A1 _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input17_I i_disable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8982__A2 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8926_ _1497_ _4429_ _0630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_196_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5796__A2 _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8857_ _4329_ _4378_ _4379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8734__A2 _4283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7808_ _3584_ _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_149_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8788_ _4316_ _4319_ _0602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_149_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4756__B1 _0930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7739_ _3441_ _3542_ _3551_ _0321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4756__C2 core_0.ew_reg_ie\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_25_Left_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8498__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5038__B core_0.fetch.prev_request_pc\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9409_ _0419_ clknet_leaf_36_i_clk core_0.execute.rf.reg_outputs\[5\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4508__B1 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7170__A1 core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output85_I net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5720__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_2520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_34_Left_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4692__C1 core_0.execute.rf.reg_outputs\[1\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_3__f_i_clk clknet_3_1_0_i_clk clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_233_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7225__A2 _3069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8422__A1 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__A3 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8084__B _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8973__A2 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6984__A1 _2492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5787__A2 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6984__B2 core_0.decode.oc_alu_mode\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8812__B _4326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__A1 net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5539__A2 _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_100_1711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_194_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_43_Left_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5944__C1 _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_111_i_clk clknet_4_7__leaf_i_clk clknet_leaf_111_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8489__A1 net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7161__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5711__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_209_3015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_209_3026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_111_1840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8661__A1 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6070_ core_0.execute.rf.reg_outputs\[5\]\[6\] net225 _2060_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input9_I i_core_int_sreg[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5021_ _1086_ _1193_ _1194_ _1162_ net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_224_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8413__A1 _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_232_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6972_ _2443_ _2451_ _2902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_232_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6975__A1 core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8711_ net75 _1740_ _1727_ _4203_ _4270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_178_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5923_ core_0.execute.rf.reg_outputs\[8\]\[8\] net346 _1913_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8716__A2 _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8642_ net78 _1740_ _4205_ _4213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6727__A1 _2660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5854_ net287 net259 _1844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_158_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4805_ core_0.ew_reg_ie\[8\] _0950_ _0956_ core_0.ew_reg_ie\[9\] _0986_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_118_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_233_3311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8573_ _4147_ _4148_ _4151_ _4152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5785_ _0942_ _0947_ _0950_ _1775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_134_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7524_ net28 _1349_ _3406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4736_ core_0.execute.pc_high_out\[5\] _0901_ _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_90_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7455_ _3360_ _0228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_151_2321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4667_ _0849_ _0850_ _0851_ _0852_ _0853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_4_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6406_ _0999_ _2378_ _2379_ _0160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7386_ _2699_ _3305_ _3306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5702__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _0789_ net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_9125_ _0137_ clknet_leaf_68_i_clk core_0.execute.sreg_priv_control.o_d\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_228_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6337_ _2220_ _2313_ _2314_ _2315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5372__I _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_3__f_i_clk_I clknet_3_1_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9056_ _0082_ clknet_leaf_86_i_clk core_0.fetch.prev_request_pc\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_177_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8652__A1 _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_90_i_clk clknet_4_15__leaf_i_clk clknet_leaf_90_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6268_ _2218_ _2253_ _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_244_3440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8007_ core_0.execute.rf.reg_outputs\[4\]\[8\] _3700_ _3704_ _3706_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5219_ core_0.ew_data\[5\] net156 _1355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6199_ _2167_ _2187_ _2188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_215_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8404__A1 _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output123_I net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_2461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__A1 _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__A2 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__C _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8909_ _4416_ _4417_ _0625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_184_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8707__A2 _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7391__A1 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6194__A2 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5941__A2 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_43_i_clk clknet_4_10__leaf_i_clk clknet_leaf_43_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_35_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8891__A1 _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7694__A2 _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58_i_clk clknet_4_11__leaf_i_clk clknet_leaf_58_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_246_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9238__CLK clknet_leaf_133_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7711__B _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5209__A1 core_0.ew_data\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4680__A2 _0680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8946__A2 _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6957__A1 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9388__CLK clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_2619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5457__I _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7382__A1 _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6185__A2 _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ _1368_ _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_5_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4521_ core_0.execute.rf.reg_outputs\[5\]\[14\] _0677_ net303 core_0.execute.rf.reg_outputs\[11\]\[14\]
+ _0718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_215_3096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7134__A1 _2074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7672__I _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_141_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7240_ _2711_ _3163_ _3164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8882__A1 _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_229_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6893__B1 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7171_ _2672_ _3095_ _3096_ _3097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_238_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__A3 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_2759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ core_0.execute.rf.reg_outputs\[5\]\[1\] _1785_ _1788_ core_0.execute.rf.reg_outputs\[3\]\[1\]
+ _2112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7437__A2 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8634__A1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6053_ core_0.execute.rf.reg_outputs\[7\]\[7\] _1773_ _2043_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5999__A2 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5004_ net73 _1180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_147_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8937__A2 _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4671__A2 net303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7070__B1 _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6955_ _2709_ _2884_ _2885_ _2886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_66_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5906_ _1895_ _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_76_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_138_Right_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_198_2888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6886_ _1290_ _2816_ _2817_ _0996_ _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_119_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer57_I _0707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8625_ core_0.execute.irq_en _4198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5837_ _1813_ _1820_ _1826_ _1827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_146_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8556_ _1685_ core_0.execute.sreg_irq_pc.o_d\[13\] net294 _2134_ _2136_ _4137_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_174_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5768_ _1517_ net186 _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7507_ core_0.ew_reg_ie\[0\] core_0.ew_reg_ie\[1\] core_0.ew_reg_ie\[2\] core_0.ew_reg_ie\[3\]
+ _3390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4719_ net104 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_44_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7125__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8487_ _1211_ _2393_ _4058_ _4076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5699_ _1703_ _0129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7438_ net124 _3168_ _3352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8873__A1 core_0.execute.pc_high_buff_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7676__A2 _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5687__A1 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7369_ net249 _2590_ _2588_ _3289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9108_ _0011_ clknet_leaf_113_i_clk core_0.execute.alu_mul_div.i_mul vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5035__C _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8627__B _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5439__A1 core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9039_ _0066_ clknet_leaf_88_i_clk core_0.fetch.out_buffer_data_instr\[27\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6100__A2 _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_max_cap217_I _0859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6147__B _2135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6939__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7600__A2 core_0.ew_data\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5478__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5611__A1 core_0.decode.i_imm_pass\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_105_Right_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_156_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7364__A1 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6167__A2 _2155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5914__A2 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7116__A1 core_0.execute.sreg_irq_pc.o_d\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8864__A1 _4383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7667__A2 _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8616__A1 _2918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8092__A2 _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4653__A2 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ core_0.execute.alu_flag_reg.o_d\[0\] _1686_ net227 _1410_ _2674_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_106_1783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_3114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6671_ core_0.execute.rf.reg_outputs\[7\]\[0\] _2611_ _2612_ core_0.execute.rf.reg_outputs\[5\]\[0\]
+ _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7355__A1 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6158__A2 _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8410_ _2712_ _4017_ _2258_ _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_183_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer7_I _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ core_0.decode.i_imm_pass\[5\] _1645_ _1647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9390_ _0400_ clknet_leaf_35_i_clk core_0.execute.rf.reg_outputs\[6\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8341_ _1539_ _3905_ _3955_ _1536_ _3956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_5553_ core_0.fetch.prev_request_pc\[9\] _1082_ _1083_ net175 _1606_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7107__A1 _1768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__S _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4504_ _0678_ net290 _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_8272_ core_0.execute.alu_mul_div.mul_res\[5\] _3887_ _3892_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7658__A2 _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5484_ core_0.fetch.out_buffer_data_instr\[11\] _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_130_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7223_ _3146_ _3147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6330__A2 _1833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_3243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8607__A1 _0859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7154_ _2713_ _3079_ _3080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_228_3254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6105_ core_0.execute.rf.reg_outputs\[3\]\[2\] _1788_ _1804_ core_0.execute.rf.reg_outputs\[11\]\[2\]
+ _2095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_70_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7085_ _2489_ _3011_ core_0.decode.oc_alu_mode\[11\] _3012_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8083__A2 _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_207_Right_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6094__A1 core_0.execute.rf.reg_outputs\[1\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7291__B1 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6036_ _1874_ net218 _2026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_226_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7830__A2 _3584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4644__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5841__A1 net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer20 net247 net248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer31 _1843_ net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_179_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer42 _0666_ net323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
Xrebuffer53 _2844_ net281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xrebuffer64 _0684_ net292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_194_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7594__A1 _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7987_ _3693_ _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_178_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer75 _1775_ net330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__8791__B1 _4217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer86 net331 net333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_193_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer97 _1756_ net344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_193_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6938_ _1743_ core_0.execute.alu_mul_div.mul_res\[3\] _2869_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_239_3383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6869_ _1896_ _1976_ _2801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_76_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5097__I _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8608_ core_0.execute.alu_flag_reg.o_d\[3\] _4167_ _4183_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7897__A2 _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9588_ _0598_ clknet_leaf_107_i_clk core_0.execute.sreg_scratch.o_d\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_2393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output190_I net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8539_ _1180_ _4121_ _4122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6430__B _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5825__I net340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__A2 _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4883__A2 _1057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_218_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8074__A2 _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7821__A2 _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5832__A1 core_0.execute.rf.reg_outputs\[1\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__B2 core_0.execute.rf.reg_outputs\[11\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8092__B _3745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6388__A2 _1925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4904__I _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6391__I net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8820__B _4326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7888__A2 _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5899__A1 core_0.decode.oc_alu_mode\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5363__A3 core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_212_3055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4571__A1 net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8837__A1 _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput107 net107 o_instr_long_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_51_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_14_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput118 net118 o_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6848__B1 _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput129 net129 o_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7950__I _3671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_130_2076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_2718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8065__A2 _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6076__B2 core_0.execute.rf.reg_outputs\[3\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7812__A2 _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4626__A2 net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7910_ _3473_ _3629_ _3649_ _0394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8890_ _4386_ _4404_ _4405_ _0618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_223_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_223_3184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7841_ _3409_ _3606_ _3610_ _0364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7772_ core_0.execute.rf.reg_outputs\[10\]\[4\] _3570_ _3568_ _3571_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4984_ net76 _1163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_74_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_195_2847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6723_ core_0.execute.rf.reg_outputs\[7\]\[6\] _2611_ _2612_ core_0.execute.rf.reg_outputs\[5\]\[6\]
+ _2659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_195_2858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9511_ _0521_ clknet_leaf_124_i_clk core_0.execute.alu_mul_div.mul_res\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_46_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7328__A1 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8730__B _4283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9442_ _0452_ clknet_leaf_45_i_clk core_0.execute.rf.reg_outputs\[3\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_128_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6654_ _1864_ _2596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7879__A2 _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6000__B2 core_0.execute.rf.reg_outputs\[9\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7346__B _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5605_ _1591_ net42 _1369_ _1636_ _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_9373_ _0383_ clknet_leaf_38_i_clk core_0.execute.rf.reg_outputs\[7\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_171_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6585_ _2526_ _2524_ _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_119_1941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5645__I _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6551__A2 _2492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8324_ _1942_ _3940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8828__A1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ _1253_ _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_131_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6839__B1 _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8255_ _3862_ _3869_ _3876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5467_ core_0.fetch.out_buffer_data_instr\[3\] net62 _1556_ _1558_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6303__A2 _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7206_ _2709_ _0789_ _3130_ _3131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8186_ _3811_ _3812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5398_ _0661_ _1486_ _1500_ _1501_ _0029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input47_I i_req_data[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7137_ _1763_ _1767_ _3063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__8056__A2 _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__I _2418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6067__A1 core_0.execute.rf.reg_outputs\[8\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7068_ _2780_ _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7803__A2 _3585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4617__A2 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6019_ _2008_ _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_2_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5290__A2 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_190_Right_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7567__A1 net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9449__CLK clknet_leaf_136_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output203_I net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_2422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6790__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8819__A1 _4324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4553__A1 core_0.execute.rf.reg_outputs\[14\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4553__B2 core_0.execute.rf.reg_outputs\[12\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5896__A4 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8866__I _4383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4856__A2 net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8047__A2 _3715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6058__A1 core_0.execute.rf.reg_outputs\[15\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6058__B2 core_0.execute.rf.reg_outputs\[1\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4835__S _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7558__A1 core_0.execute.rf.reg_outputs\[15\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_103_1753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6781__A2 _2371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4792__A1 core_0.ew_reg_ie\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4792__B2 core_0.ew_reg_ie\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7730__A1 _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_190_2788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6370_ _1669_ _2342_ _2343_ _2344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__5592__I0 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5321_ core_0.decode.i_instr_l\[9\] _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_23_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8040_ core_0.execute.rf.reg_outputs\[3\]\[6\] _3722_ _3718_ _3725_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5252_ core_0.dec_jump_cond_code\[1\] core_0.dec_jump_cond_code\[0\] core_0.execute.alu_flag_reg.o_d\[2\]
+ _1373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_121_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8038__A2 _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_225_3213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5183_ _1263_ _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_223_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__A1 core_0.ew_reg_ie\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8942_ core_0.decode.i_imm_pass\[3\] _1264_ _4439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_2234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8873_ core_0.execute.pc_high_buff_out\[1\] _4386_ _3797_ _4393_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8210__A2 _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7824_ core_0.execute.rf.reg_outputs\[9\]\[11\] _3591_ _3595_ _3600_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5024__A2 _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4967_ core_0.fetch.prev_request_pc\[3\] _1147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7755_ core_0.execute.rf.reg_outputs\[11\]\[14\] _3541_ _3554_ _3560_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_236_3342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6772__A2 net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6706_ core_0.execute.rf.reg_outputs\[1\]\[4\] _2608_ _2609_ core_0.execute.rf.reg_outputs\[3\]\[4\]
+ _2644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4783__A1 _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7686_ _3519_ _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4898_ core_0.fetch.dbg_out _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6637_ _1769_ _2578_ _1863_ _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_9425_ _0435_ clknet_leaf_23_i_clk core_0.execute.rf.reg_outputs\[4\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7721__A1 _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_2363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4535__B2 core_0.execute.rf.reg_outputs\[9\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6568_ _1759_ _2349_ _2510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XPHY_EDGE_ROW_89_Left_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_9356_ _0366_ clknet_leaf_9_i_clk core_0.execute.rf.reg_outputs\[8\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5519_ _1055_ _1552_ _1586_ _0066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8686__I _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8307_ _3863_ _3924_ _3925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7804__B _3580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9287_ _0297_ clknet_leaf_152_i_clk core_0.execute.rf.reg_outputs\[13\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6499_ _2437_ _2440_ _2441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_219_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6288__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9121__CLK clknet_leaf_64_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8238_ core_0.execute.alu_mul_div.mul_res\[3\] _3832_ _3861_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_7_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8029__A2 _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4719__I net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8169_ _3465_ _3781_ _3798_ _0504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_245_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_226_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_2492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5799__B1 net340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_98_Left_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_241_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5799__C2 core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6460__A1 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6870__S _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8201__A2 _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5015__A2 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8504__A3 _4076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__A2 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7712__A1 _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__A1 _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7779__A1 _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8440__A2 _4031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6451__A1 _1175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__A2 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_220_3154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5870_ _1328_ net254 _1860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4821_ net155 _1002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_201_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8743__A3 _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7951__A1 core_0.execute.rf.reg_outputs\[5\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6754__A2 net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_192_2817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7540_ _3382_ core_0.ew_data\[3\] _3419_ _3420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_200_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4752_ core_0.ew_reg_ie\[0\] _0665_ net271 _0933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5962__B1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7471_ core_0.dec_rf_ie\[4\] core_0.ew_reg_ie\[4\] _3366_ _3369_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4683_ core_0.execute.rf.reg_outputs\[14\]\[2\] net262 _0716_ _0868_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6506__A2 _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9210_ _0221_ clknet_leaf_55_i_clk net125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6422_ _2389_ _2385_ _2390_ _0165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_1900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_231_3283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9141_ _0153_ clknet_leaf_99_i_clk core_0.execute.alu_mul_div.div_cur\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_12_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__A1 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6353_ _2142_ _2256_ _2328_ _2229_ _0158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7624__B _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5304_ _1423_ _1424_ _1425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9072_ _0097_ clknet_leaf_128_i_clk core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_122_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6284_ _2188_ _2267_ _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8023_ core_0.ew_reg_ie\[3\] _3394_ _3714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
X_5235_ core_0.ew_data\[5\] core_0.ew_data\[13\] _1349_ _1363_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_227_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_243_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6690__A1 core_0.execute.rf.reg_outputs\[7\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6690__B2 core_0.execute.rf.reg_outputs\[5\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5166_ core_0.decode.i_instr_l\[5\] _1245_ _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_236_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8431__A2 _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5097_ _1249_ _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_223_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5245__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8925_ core_0.dec_used_operands\[0\] _1229_ _4423_ _4428_ _4429_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_clkbuf_leaf_136_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6993__A2 core_0.execute.alu_mul_div.i_mod vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8856_ core_0.execute.pc_high_out\[7\] _4377_ _4378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_149_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7807_ _3421_ _3585_ _3590_ _0350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8787_ core_0.execute.sreg_irq_flags.o_d\[2\] _4217_ core_0.execute.sreg_irq_flags.i_d\[2\]
+ _4319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_176_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5999_ core_0.execute.rf.reg_outputs\[8\]\[12\] _1794_ _1776_ core_0.execute.rf.reg_outputs\[4\]\[12\]
+ _1989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7942__A1 core_0.execute.rf.reg_outputs\[6\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4756__A1 core_0.ew_reg_ie\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4756__B2 core_0.ew_reg_ie\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7738_ core_0.execute.rf.reg_outputs\[11\]\[6\] _3548_ _3539_ _3551_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8498__A2 _4040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7669_ _3454_ _3497_ _3510_ _0292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_191_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9408_ _0418_ clknet_leaf_37_i_clk core_0.execute.rf.reg_outputs\[5\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_61_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4508__B2 core_0.execute.rf.reg_outputs\[9\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7170__A2 net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9339_ _0349_ clknet_leaf_155_i_clk core_0.execute.rf.reg_outputs\[9\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output78_I net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_2521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8670__A2 _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6681__A1 _2614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4692__B1 net318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4692__C2 _0693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A4 _0980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A1 _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8973__A3 _1272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7709__B _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_2650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6736__A2 _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4747__A1 _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5944__B1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__C2 core_0.execute.rf.reg_outputs\[3\]\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8489__A2 _1738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7161__A2 _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5172__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7163__C _2689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_209_3016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8661__A2 _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6121__B1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ net86 _1085_ _1194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_225_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_119_Right_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_136_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5411__C _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _2900_ _2901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_88_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_2960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8710_ _1658_ _4265_ _4269_ _0574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_177_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _1899_ net213 _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8177__A1 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8722__C _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ net313 net205 _1842_ _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_8641_ _1661_ _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_220_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9537__D _0547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7924__A1 _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4804_ core_0.ew_reg_ie\[10\] _0959_ _0960_ core_0.ew_reg_ie\[11\] _0985_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_63_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_1981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_233_3312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8572_ _4039_ _4150_ _4151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5784_ core_0.execute.rf.reg_outputs\[7\]\[0\] _1773_ _1774_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_16_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6242__C _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7523_ net36 _1347_ _3405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4735_ core_0.execute.prev_pc_high\[7\] _0911_ net111 _0913_ _0915_ _0916_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_43_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7454_ net117 _3225_ _2415_ _3360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ core_0.execute.rf.reg_outputs\[7\]\[3\] _0683_ net257 core_0.execute.rf.reg_outputs\[8\]\[3\]
+ _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_151_2322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6405_ _0999_ _1829_ _2379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7385_ _3270_ _3303_ _3305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4597_ net102 _0666_ _0788_ _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_3_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_62_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6336_ _2299_ _2220_ _2314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9124_ _0136_ clknet_leaf_108_i_clk core_0.execute.sreg_priv_control.o_d\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6685__S _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9055_ _0081_ clknet_leaf_86_i_clk core_0.fetch.prev_request_pc\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6267_ _2246_ _2251_ _2252_ _2253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_244_3441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6663__A1 _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5218_ _1354_ net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8006_ _3446_ _3694_ _3705_ _0434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_209_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ core_0.execute.alu_mul_div.div_cur\[6\] _1843_ _2187_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_149_2295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_208_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5149_ _1234_ _1243_ _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_98_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_162_2451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_2462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4977__A1 core_0.fetch.prev_request_pc\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8908_ _0038_ _1240_ _1275_ _4417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_196_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8168__A1 net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8839_ core_0.execute.pc_high_out\[5\] _4362_ _4363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7915__A1 _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_173_2591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8340__A1 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8891__A2 _4383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_219_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6103__B1 _1776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4665__B1 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5209__A2 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6406__A1 _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__C _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__A1 core_0.fetch.prev_request_pc\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8159__A1 net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6709__A2 _2640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7906__A1 _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8954__I0 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5917__B1 _1794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5393__A1 _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4520_ core_0.execute.rf.reg_outputs\[6\]\[14\] _0670_ _0673_ core_0.execute.rf.reg_outputs\[2\]\[14\]
+ _0717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_81_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_215_3097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5145__A1 _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_229_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6893__A1 core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7170_ core_0.dec_mem_access net207 _3096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6893__B2 net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6121_ core_0.execute.rf.reg_outputs\[14\]\[1\] _1802_ _1776_ core_0.execute.rf.reg_outputs\[4\]\[1\]
+ _2111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__8634__A2 _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8717__C _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6052_ _2026_ _2041_ _2042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_7_Right_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_225_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4656__B1 _0710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5003_ _1175_ _1165_ _1179_ _1162_ net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_178_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone78_A1 net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _2709_ net217 _2885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5620__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5905_ _1753_ _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_198_2889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _2124_ core_0.execute.alu_mul_div.mul_res\[2\] _2817_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8024__I _3714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8624_ _4196_ _4197_ _0560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_174_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5836_ core_0.execute.rf.reg_outputs\[15\]\[15\] _0945_ _1821_ core_0.execute.rf.reg_outputs\[7\]\[15\]
+ _1825_ _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_63_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone22_I _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8570__A1 _1163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5384__A1 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8555_ _4080_ _3261_ _4136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5767_ _1755_ _1756_ _1757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__5584__S _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7506_ core_0.ew_reg_ie\[4\] core_0.ew_reg_ie\[5\] core_0.ew_reg_ie\[6\] core_0.ew_reg_ie\[7\]
+ _3389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4718_ core_0.execute.prev_sys _0899_ _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_20_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8486_ _4073_ _4075_ _4051_ _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5698_ net193 _1698_ _1701_ core_0.execute.sreg_priv_control.o_d\[0\] _1702_ _1703_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_17_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6479__I _2418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7437_ _2616_ _2873_ _3351_ _0219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4649_ net251 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_75_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8873__A2 _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5687__A2 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7368_ _2587_ net272 _2987_ _3288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_203_Left_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9107_ _0010_ clknet_leaf_131_i_clk core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_229_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6319_ _2297_ _2298_ _0154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7299_ _2124_ core_0.execute.alu_mul_div.mul_res\[12\] _3221_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5439__A2 _1001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9038_ _0065_ clknet_leaf_88_i_clk core_0.fetch.out_buffer_data_instr\[26\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_216_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_110_i_clk clknet_4_6__leaf_i_clk clknet_leaf_110_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6147__C _2136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6939__A2 _2868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5986__C _1897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_125_i_clk clknet_4_5__leaf_i_clk clknet_leaf_125_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5611__A2 _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_223_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7364__A2 _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8561__A1 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__B2 _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7116__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A1 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6875__A1 _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8616__A2 _2949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6627__A1 _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4638__B1 net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6338__B _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4637__I _0825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5850__A2 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7052__A1 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_10_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_201_2930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__A2 _1634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_3115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6670_ _0947_ _0957_ _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_46_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8552__A1 net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5621_ _1032_ _1615_ _1646_ _0108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5366__A1 core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5552_ _1597_ _1605_ _0080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8340_ _1539_ _3954_ _3955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_135_2136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7107__A2 _2563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ core_0.execute.rf.reg_outputs\[3\]\[15\] _0698_ _0700_ core_0.execute.rf.reg_outputs\[12\]\[15\]
+ _0701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_53_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8271_ _3875_ _3832_ _3891_ _0513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5118__A1 core_0.decode.i_instr_l\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5483_ _1566_ _0050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7222_ _1285_ _2155_ _3144_ core_0.decode.oc_alu_mode\[9\] _3145_ _3146_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_41_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7153_ _3059_ _3064_ _3078_ _3079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_TAPCELL_ROW_228_3244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6618__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6104_ core_0.execute.rf.reg_outputs\[15\]\[2\] _0945_ _1779_ core_0.execute.rf.reg_outputs\[1\]\[2\]
+ _2094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XPHY_EDGE_ROW_171_Right_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7084_ _2517_ _2970_ _3011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_241_3400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4547__I net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6094__A2 _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6035_ net97 _1771_ _2015_ _2024_ _2025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__7291__B2 _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5841__A2 net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_61_Left_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xrebuffer10 _1853_ net238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_42_i_clk clknet_4_10__leaf_i_clk clknet_leaf_42_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xrebuffer21 _2598_ net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_240_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer32 net259 net260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_240_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xrebuffer43 _0666_ net324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xrebuffer54 _2814_ net282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7986_ core_0.ew_reg_ie\[4\] _3394_ _3693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
Xrebuffer65 _0688_ net326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__8791__A1 core_0.execute.irq_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7594__A2 _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer76 net195 net304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__8791__B2 core_0.execute.sreg_irq_flags.o_d\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer87 _3030_ net334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_1
XFILLER_0_77_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6937_ _2759_ net281 _2855_ _2867_ _2868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xrebuffer98 _1793_ net345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_1
XFILLER_0_49_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_3384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_57_i_clk clknet_4_11__leaf_i_clk clknet_leaf_57_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6868_ _1309_ _2791_ _2797_ _2011_ _2799_ _2800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_193_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8543__A1 _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8607_ _0859_ _4165_ _4177_ _4181_ _4167_ _4182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_81_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9228__CLK clknet_leaf_144_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5819_ core_0.execute.rf.reg_outputs\[14\]\[0\] _1802_ _1804_ core_0.execute.rf.reg_outputs\[11\]\[0\]
+ _1808_ _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_9587_ _0597_ clknet_leaf_107_i_clk core_0.execute.sreg_scratch.o_d\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6799_ _1882_ _2040_ _2732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_2394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8538_ _1185_ _4113_ _4121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_45_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_70_Left_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output183_I net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_170_2550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8846__A2 core_0.execute.pc_high_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8469_ _1738_ _4060_ _4047_ _4061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4580__A2 _0685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__A1 core_0.ew_data\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5046__C _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4883__A3 _1060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7261__C _3073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_216_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5832__A2 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4891__I0 net59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7768__I _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_2690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8782__A1 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7585__A2 _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5596__A1 _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7337__A2 _3256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_109_Left_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7717__B _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_212_3056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4571__A2 _0666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput108 net108 o_instr_long_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6848__A1 core_0.execute.sreg_data_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput119 net119 o_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6848__B2 net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_2719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_118_Left_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput90 net90 dbg_r0[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_208_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7273__A1 net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6076__A2 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7273__B2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_1813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_223_3185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7025__A1 _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7840_ core_0.execute.rf.reg_outputs\[8\]\[1\] _3607_ _3609_ _3610_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_203_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8773__A1 core_0.execute.sreg_scratch.o_d\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5587__A1 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7771_ _3562_ _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_148_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4983_ _1086_ _1160_ _1161_ _1162_ net166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_19_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9510_ _0520_ clknet_leaf_123_i_clk core_0.execute.alu_mul_div.mul_res\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6722_ core_0.execute.rf.reg_outputs\[1\]\[6\] _2608_ _2609_ core_0.execute.rf.reg_outputs\[3\]\[6\]
+ _2658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_195_2848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_127_Left_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8525__A1 _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7328__A2 _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9441_ _0451_ clknet_leaf_45_i_clk core_0.execute.rf.reg_outputs\[3\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5339__A1 _1257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7627__B _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6653_ _1329_ _1973_ _2595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6000__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5604_ _1591_ _1571_ _1636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9372_ _0382_ clknet_leaf_9_i_clk core_0.execute.rf.reg_outputs\[7\]\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_116_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_240_Right_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6584_ _2525_ _2456_ _2526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_30_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6250__C _2229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_1942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8323_ _3939_ _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5535_ _1594_ _1596_ _1435_ _0072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4562__A2 _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8828__A2 _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6839__A1 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6839__B2 core_0.execute.pc_high_buff_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5466_ _1557_ _0042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8254_ core_0.execute.alu_mul_div.mul_res\[5\] _3875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_112_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7205_ _2708_ _3129_ _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_136_Left_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5397_ _1249_ _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5661__I core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8185_ _3806_ _3807_ _3809_ _3810_ _1536_ _3811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_112_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7136_ _2010_ _1894_ _2561_ _1865_ _3062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_226_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7067_ _2829_ _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_213_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ net314 net201 _2007_ _2008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_2_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7588__I _3459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7016__A1 _2795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5290__A3 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8764__A1 _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_145_Left_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5578__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7969_ core_0.execute.rf.reg_outputs\[5\]\[8\] _3679_ _3677_ _3684_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9050__CLK clknet_leaf_92_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_2423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8516__A1 _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9639_ _0649_ clknet_leaf_95_i_clk net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_80_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_220_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4553__A2 _0686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5502__A1 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5571__I _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6058__A2 _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5805__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7558__A2 _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_103_1743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8507__A1 _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9543__CLK clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4792__A2 _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__B _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7730__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer1 _0713_ net229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_190_2789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5592__I1 core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5320_ _1437_ _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_106_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5251_ core_0.dec_jump_cond_code\[3\] _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_121_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_1883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _1329_ _1251_ _1330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_225_3214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7246__A1 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6049__A2 _2038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8294__I0 core_0.execute.alu_mul_div.mul_res\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7797__A2 _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8941_ _1405_ _0038_ _4438_ _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_143_2224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8872_ net200 _4387_ _4391_ _4392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4480__A1 net301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8746__A1 core_0.execute.sreg_scratch.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7823_ _3457_ _3586_ _3599_ _0357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7754_ _3466_ _3543_ _3559_ _0328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4966_ _1145_ _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_46_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_236_3343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6705_ _2422_ _2641_ _2643_ _0194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7685_ _3519_ _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4783__A2 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _0895_ _0896_ _1008_ _1077_ _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_74_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9424_ _0434_ clknet_leaf_24_i_clk core_0.execute.rf.reg_outputs\[4\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6636_ _2026_ _2091_ _2578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7721__A2 _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_2364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4535__A2 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9355_ _0365_ clknet_leaf_0_i_clk core_0.execute.rf.reg_outputs\[8\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5732__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6567_ _1751_ _2102_ _2509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5592__S _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8306_ _1925_ _3827_ _3923_ _3924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_132_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5518_ net56 _1556_ _1586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9286_ _0296_ clknet_leaf_152_i_clk core_0.execute.rf.reg_outputs\[13\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6498_ _2438_ _2439_ _2440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6288__A2 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__B _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8237_ _2349_ _3833_ _3859_ _3860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_7_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5449_ core_0.execute.alu_mul_div.cbit\[1\] _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_218_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8168_ net91 _3787_ _3797_ _3798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_196_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7237__A1 _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9416__CLK clknet_leaf_136_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7820__B _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7119_ _3041_ _3043_ _3045_ _3046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8099_ core_0.ew_reg_ie\[1\] _3394_ _3758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7788__A2 _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8985__A1 _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8635__C _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5799__A1 core_0.execute.rf.reg_outputs\[5\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_2493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5799__B2 core_0.execute.rf.reg_outputs\[9\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_153_Left_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6460__A2 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8207__I _3830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4471__A1 _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8737__A1 core_0.execute.trap_flag vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_57_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8651__B _1661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7267__B core_0.execute.alu_mul_div.i_div vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5971__A1 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4470__I core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7712__A2 _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5723__A1 core_0.execute.sreg_priv_control.o_d\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5723__B2 _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6397__I _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7228__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_245_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7779__A2 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6451__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_220_3155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7400__A1 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7400__B2 _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4820_ _0999_ _1000_ _1001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_32_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_192_2818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7951__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6754__A3 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4751_ core_0.ew_reg_ie\[4\] _0665_ _0930_ core_0.ew_reg_ie\[5\] _0931_ core_0.ew_reg_ie\[7\]
+ _0932_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_64_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5962__A1 core_0.execute.rf.reg_outputs\[5\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4765__A2 core_0.execute.sreg_long_ptr_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7470_ _3368_ _0235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4682_ core_0.execute.rf.reg_outputs\[10\]\[2\] _0695_ net257 core_0.execute.rf.reg_outputs\[8\]\[2\]
+ _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5409__C _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8900__A1 _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7703__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7905__B _3636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6421_ core_0.execute.mem_stage_pc\[1\] _2386_ _2387_ _2390_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_40_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5714__A1 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_231_3284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9140_ _0152_ clknet_leaf_99_i_clk core_0.execute.alu_mul_div.div_cur\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6352_ core_0.execute.alu_mul_div.div_cur\[13\] _2246_ _2326_ _2327_ _2256_ _2328_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_24_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5303_ net192 net179 net178 net181 _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_9071_ _0096_ clknet_leaf_128_i_clk core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6283_ _2266_ _2260_ _2190_ _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8022_ _3472_ _3695_ _3713_ _0442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5234_ _1362_ net141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_215_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6690__A2 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5165_ _1233_ _1230_ _1313_ _1315_ _0008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_243_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4983__C _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9589__CLK clknet_leaf_108_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _1231_ _1248_ _1252_ _0004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6256__B _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8924_ _1229_ _1335_ _4427_ _4428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclone6 net314 net246 _1845_ net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_196_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__A4 _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8855_ core_0.execute.pc_high_out\[6\] core_0.execute.pc_high_out\[5\] core_0.execute.pc_high_out\[4\]
+ _4349_ _4377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_182_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8195__A2 core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7806_ core_0.execute.rf.reg_outputs\[9\]\[3\] _3586_ _3580_ _3590_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8786_ _4316_ _4318_ _0601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5998_ _0730_ _1962_ _1987_ _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__7942__A2 _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5953__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7737_ _3435_ _3542_ _3550_ _0320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4949_ _1107_ _1108_ _1111_ _1114_ _1129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_35_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7668_ core_0.execute.rf.reg_outputs\[13\]\[9\] _3504_ _3500_ _3510_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9407_ _0417_ clknet_leaf_36_i_clk core_0.execute.rf.reg_outputs\[5\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6619_ _1895_ _1882_ _2561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4508__A2 _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5705__A1 core_0.execute.sreg_long_ptr_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5705__B2 _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7599_ _3403_ _3466_ _3468_ _0264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9338_ _0348_ clknet_leaf_155_i_clk core_0.execute.rf.reg_outputs\[9\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9269_ _0279_ clknet_leaf_151_i_clk core_0.execute.rf.reg_outputs\[14\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_2511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_2522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6130__A1 _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A2 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7630__A1 _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7481__I1 core_0.ew_reg_ie\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_195_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_2651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A2 net301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7725__B _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7697__A1 _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7449__A1 _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5245__B _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_209_3017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_2780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7621__A1 _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6970_ _2567_ _2583_ _2856_ _1865_ _2900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_45_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_2961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5921_ net102 _1772_ _1903_ _1910_ _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_76_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7686__I _3519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8291__B _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8177__A2 _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8640_ core_0.execute.sreg_irq_pc.o_d\[1\] _4210_ _4211_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ _1517_ net189 _1842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_146_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7924__A2 _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4803_ _0962_ _0982_ _0983_ _0984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_152_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4738__A2 _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5935__A1 net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8571_ _2411_ _4149_ _4150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5783_ _0942_ _0947_ _0960_ _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_233_3313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7522_ _3397_ _3402_ _3404_ _0251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4734_ core_0.execute.prev_pc_high\[7\] _0911_ _0914_ core_0.execute.prev_pc_high\[6\]
+ _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_173_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7688__A1 _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7635__B _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7453_ _2616_ _3192_ _3359_ _0227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ core_0.execute.rf.reg_outputs\[2\]\[3\] net250 _0705_ core_0.execute.rf.reg_outputs\[9\]\[3\]
+ _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__9261__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_151_2323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6404_ core_0.execute.alu_mul_div.div_cur\[0\] _2218_ _2375_ _2377_ _2378_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_3_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7384_ _3270_ _3303_ _3304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4596_ _0782_ _0787_ _0788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_101_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9123_ _0135_ clknet_leaf_109_i_clk core_0.execute.sreg_priv_control.o_d\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6335_ _1547_ _2303_ _2312_ _2313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4910__A2 _1016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9054_ _0080_ clknet_leaf_85_i_clk core_0.fetch.prev_request_pc\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__6112__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6266_ core_0.execute.alu_mul_div.div_cur\[3\] _2224_ _2252_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8005_ core_0.execute.rf.reg_outputs\[4\]\[7\] _3700_ _3704_ _3705_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_244_3442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5217_ core_0.ew_data\[4\] net156 _1354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6663__A2 _1866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7860__A1 _3457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6197_ _2185_ net342 _2186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8185__C _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5148_ _1247_ _1275_ _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input22_I i_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7612__A1 _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_2452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5079_ core_0.decode.i_instr_l\[3\] _1235_ _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_193_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8907_ core_0.dec_sys _1251_ _4416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_211_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7596__I _3465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8168__A2 _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8838_ core_0.execute.pc_high_out\[4\] _4349_ _4362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7915__A2 _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4729__A2 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5926__A1 core_0.execute.rf.reg_outputs\[7\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8769_ _0777_ _4295_ _4308_ _4307_ _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_19_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7679__A1 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_185_Right_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_173_2592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output90_I net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__A1 _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7851__A1 core_0.execute.rf.reg_outputs\[8\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4665__B2 core_0.execute.rf.reg_outputs\[9\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7603__A1 _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7454__I1 _3225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4968__A2 core_0.fetch.prev_request_pc\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8159__A2 _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7906__A2 _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6343__C _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8954__I1 core_0.decode.i_imm_pass\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5393__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_215_3087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_215_3098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_152_Right_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6342__A1 _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6893__A2 _2770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8095__A1 _3469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6120_ core_0.execute.rf.reg_outputs\[9\]\[1\] _1815_ _1781_ core_0.execute.rf.reg_outputs\[10\]\[1\]
+ _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_193_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6051_ _1874_ _2040_ _2041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_56_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__B2 core_0.execute.rf.reg_outputs\[8\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5002_ _1176_ _1146_ _1178_ _1164_ _1179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA_clone78_A2 net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_221_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7070__A2 _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _2711_ _2873_ _2883_ _2884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9627__CLK clknet_leaf_110_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5904_ net325 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_9_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6884_ _2812_ _2815_ _2816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_159_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8623_ core_0.execute.alu_flag_reg.o_d\[4\] _4167_ _1431_ _4197_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5835_ _1822_ _1823_ _1824_ _1825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_91_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8570__A2 _4133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8554_ _4133_ _4134_ _4135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5766_ net87 _0667_ _0885_ _0889_ _1518_ _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_91_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7505_ _3387_ core_0.ew_submit _3388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_115_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4717_ _0897_ _0898_ _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8485_ _4047_ _4074_ _4075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5697_ _0891_ _0900_ _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_20_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7436_ net123 _3168_ _3351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4648_ net98 _0667_ _0830_ _0835_ _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_130_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout1 _1754_ net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_102_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7367_ _2979_ _3069_ _3286_ _3287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_97_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4579_ core_0.execute.rf.reg_outputs\[6\]\[10\] net223 _0692_ core_0.execute.rf.reg_outputs\[1\]\[10\]
+ _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4895__A1 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9106_ _0009_ clknet_leaf_111_i_clk core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6318_ core_0.execute.alu_mul_div.div_cur\[10\] _2219_ _0999_ _2298_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7298_ _3208_ _3211_ _3215_ _3219_ _3220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_9037_ _0064_ clknet_leaf_87_i_clk core_0.fetch.out_buffer_data_instr\[25\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7833__A1 _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6249_ core_0.execute.alu_mul_div.div_cur\[2\] _2218_ _2237_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_228_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6444__B _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__I _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4743__I core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8010__A1 _3453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_2610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_223_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8561__A2 _4133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__A2 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8077__A1 _3434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_186_2750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6627__A2 _1757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7052__A2 _2979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5063__A1 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_2920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_221_Right_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_175_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8001__A1 _3434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_3116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8552__A2 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5620_ core_0.decode.i_imm_pass\[4\] _1645_ _1646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5366__A2 _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4574__B1 _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5551_ core_0.fetch.prev_request_pc\[8\] _1595_ _1084_ net174 _1605_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_135_2137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4502_ _0699_ _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_13_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8270_ _2040_ _3833_ _3890_ _3830_ _3891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6315__A1 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ core_0.fetch.out_buffer_data_instr\[10\] net39 _1559_ _1566_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8855__A3 core_0.execute.pc_high_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7221_ _1942_ _3072_ _3073_ _3145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7152_ _3067_ _3068_ _3077_ _3078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_228_3245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6618__A2 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6103_ core_0.execute.rf.reg_outputs\[14\]\[2\] _1802_ _1776_ core_0.execute.rf.reg_outputs\[4\]\[2\]
+ _2093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7083_ _2839_ _3009_ _3010_ _0206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_225_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_241_3401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5826__B1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6094__A3 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6034_ _2016_ _2021_ _2022_ _2023_ _2024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_174_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_2266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_241_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4991__C _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer11 net238 net239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xrebuffer22 _0709_ net316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xrebuffer33 net259 net261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer44 _2986_ net272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer55 net267 net283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7985_ _3472_ _3673_ _3692_ _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5054__A1 net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer66 net197 net294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xrebuffer77 net304 net305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8791__A2 net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8035__I _3714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6936_ _1894_ _2859_ _2866_ _2810_ _2867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_49_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer88 _1796_ net335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_77_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer99 net345 net346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_194_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_239_3385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6867_ _1880_ _2792_ _2798_ _1292_ _2799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6003__B1 _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7874__I _3627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8606_ _4165_ _4178_ _4180_ _4181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_81_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5818_ _1805_ _0950_ _1790_ _1806_ _1807_ _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_64_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5357__A2 _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6554__A1 _2074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9586_ _0596_ clknet_leaf_110_i_clk core_0.execute.sreg_scratch.o_d\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6798_ _1899_ _2360_ _2730_ _2731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer101 core_0.dec_r_reg_sel\[1\] net348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_134_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8537_ _0765_ _4048_ _3192_ _2133_ _3197_ _4120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_51_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4565__B1 _0707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_2395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5749_ _1226_ _1738_ _1739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_2551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8468_ _4058_ _4059_ _4060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7419_ _3336_ _3337_ _3338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output176_I net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8399_ _3828_ _4008_ _4009_ _4010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4868__A1 _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_217_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7806__A1 core_0.execute.rf.reg_outputs\[9\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__A4 _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_181_2680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9188__D _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5045__A1 _1031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_127_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clone6_A1 net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4556__B1 _0710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_212_3057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9322__CLK clknet_leaf_1_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput109 net109 o_instr_long_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6848__A2 _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4859__A1 _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5520__A2 _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9472__CLK clknet_leaf_37_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput80 net80 dbg_pc[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput91 net91 dbg_r0[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_207_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_208_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7273__A2 _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8470__A1 _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_222_Left_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6863__I core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_1814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_223_3186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6084__I0 _1687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8773__A2 _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7770_ _3421_ _3563_ _3569_ _0334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4982_ _1080_ _1162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__5587__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6784__A1 _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6721_ _2422_ _2656_ _2657_ _0196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_2849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9440_ _0450_ clknet_leaf_44_i_clk core_0.execute.rf.reg_outputs\[3\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_190_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6652_ _2588_ _2590_ _2593_ _2594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_73_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_231_Left_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5603_ core_0.decode.i_instr_l\[13\] _1616_ _1635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9371_ _0381_ clknet_leaf_4_i_clk core_0.execute.rf.reg_outputs\[7\]\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_27_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6583_ _2428_ _2054_ _2525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8322_ core_0.execute.alu_mul_div.mul_res\[9\] _3938_ _3863_ _3939_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_30_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8289__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ _1595_ net160 _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8739__B _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7643__B _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8253_ _3862_ _3863_ _3827_ net218 _3874_ _0512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__6839__A2 _2770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5465_ core_0.fetch.out_buffer_data_instr\[2\] net59 _1556_ _1557_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7204_ _2710_ _3120_ _3127_ _3128_ _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_246_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5511__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_124_i_clk clknet_4_5__leaf_i_clk clknet_leaf_124_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8184_ _1674_ _1749_ _1851_ _2372_ _2140_ _3810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5396_ core_0.decode.i_imm_pass\[3\] _1488_ _1494_ core_0.decode.i_instr_l\[14\]
+ _1495_ _1500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_7135_ _3060_ _2585_ _3061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_240_Left_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7066_ core_0.execute.alu_mul_div.div_cur\[6\] _1317_ _2991_ _2993_ _2994_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6017_ net313 _1404_ _2007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_139_i_clk clknet_4_1__leaf_i_clk clknet_leaf_139_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_2_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8213__A1 _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8764__A2 _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7968_ _3446_ _3672_ _3683_ _0418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5578__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_2424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4786__B1 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6919_ _2849_ _2510_ _2850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7818__B _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7899_ core_0.execute.rf.reg_outputs\[7\]\[11\] _3634_ _3636_ _3643_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6527__A1 net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9638_ _0648_ clknet_leaf_96_i_clk net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_174_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4538__B1 _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9569_ _0579_ clknet_leaf_63_i_clk core_0.execute.sreg_jtr_buff.o_d\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_53_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5502__A2 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_229_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8452__A1 _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8755__A2 _4300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6766__A1 _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5569__A2 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6632__B _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_103_1744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_172_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6518__A1 _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4529__B1 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7191__A1 _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer2 net229 net230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5741__A2 _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_41_i_clk clknet_4_10__leaf_i_clk clknet_leaf_41_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_239_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5250_ _1006_ _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__8691__A1 core_0.execute.sreg_irq_pc.o_d\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4701__B1 net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5181_ _1328_ _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_225_3215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_56_i_clk clknet_4_11__leaf_i_clk clknet_leaf_56_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_208_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8443__A1 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8940_ core_0.decode.i_imm_pass\[2\] _1293_ _4438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_2225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8871_ _0905_ _4387_ _4391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5009__A1 _1180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_207_2992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4480__A2 core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8746__A2 _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7822_ core_0.execute.rf.reg_outputs\[9\]\[10\] _3591_ _3595_ _3599_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7753_ core_0.execute.rf.reg_outputs\[11\]\[13\] _3548_ _3554_ _3559_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ _1133_ _1141_ _1144_ _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_164_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6704_ net133 _2642_ _2643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_236_3344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__A1 _1759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7684_ core_0.ew_reg_ie\[12\] _3395_ _3519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_191_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4896_ _1067_ _1070_ _1071_ _1076_ _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_116_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9423_ _0433_ clknet_leaf_23_i_clk core_0.execute.rf.reg_outputs\[4\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6635_ _2571_ _2573_ _2576_ _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_fanout1_I _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9354_ _0364_ clknet_leaf_0_i_clk core_0.execute.rf.reg_outputs\[8\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_2365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6566_ _1895_ _2505_ _2506_ _2507_ _2508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_144_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer25_I _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8469__B _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8305_ _3919_ _3921_ _3922_ _3923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5517_ _1035_ _1552_ _1585_ _0065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9285_ _0295_ clknet_leaf_153_i_clk core_0.execute.rf.reg_outputs\[13\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6497_ _1841_ _2054_ _2439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__8188__C _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7_0_i_clk clknet_0_i_clk clknet_3_7_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8236_ _3853_ _3857_ _3858_ _3859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8682__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5448_ _1542_ _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input52_I i_req_data[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__A1 net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8167_ _0891_ _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_245_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5379_ _1482_ _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_100_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7118_ core_0.execute.pc_high_buff_out\[7\] _2771_ _3044_ core_0.execute.sreg_scratch.o_d\[7\]
+ _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_242_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8098_ _3472_ _3738_ _3757_ _0474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5248__A1 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7049_ _2010_ _2806_ _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_29_Right_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6996__A1 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5799__A2 _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_2494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__A2 _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8737__A2 _1418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6748__A1 core_0.execute.sreg_priv_control.o_d\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6452__B _2404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5971__A2 _0951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Right_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5023__I1 _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6920__A1 _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5723__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8673__A1 _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7228__A2 _3150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8425__A1 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_47_Right_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8976__A2 _4456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4926__I core_0.fetch.prev_request_pc\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5023__S _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8189__B1 _1837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_220_3156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8728__A2 _4283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_199_Right_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_200_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5411__A1 _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6754__A4 _2687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_192_2819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4750_ _0668_ _0675_ _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XPHY_EDGE_ROW_56_Right_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_64_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5962__A2 _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4681_ core_0.execute.rf.reg_outputs\[9\]\[2\] _0705_ _0708_ core_0.execute.rf.reg_outputs\[13\]\[2\]
+ _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_119_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8900__A2 _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6420_ net78 _2389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_40_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_231_3285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _1547_ _2318_ _2224_ _2327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_141_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4610__B _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ net180 net183 net182 _1423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__8664__A1 _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9070_ _0095_ clknet_leaf_104_i_clk core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6282_ _2182_ _2266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8021_ core_0.execute.rf.reg_outputs\[4\]\[15\] _3693_ _3704_ _3713_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5233_ core_0.ew_data\[4\] core_0.ew_data\[12\] _1349_ _1362_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_65_Right_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7219__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8416__A1 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ _1314_ _1250_ _1315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ core_0.decode.oc_alu_mode\[1\] _1251_ _1252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8923_ _1450_ _1525_ _4426_ _4427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_196_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8719__A2 _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8854_ core_0.execute.pc_high_out\[7\] _4376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_182_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7805_ _3415_ _3585_ _3589_ _0349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8785_ core_0.execute.sreg_irq_flags.o_d\[1\] _4317_ core_0.execute.prev_sys _4318_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_166_Right_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _1979_ _1986_ _1987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_74_Right_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_148_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7736_ core_0.execute.rf.reg_outputs\[11\]\[5\] _3548_ _3539_ _3550_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4948_ _1087_ _1103_ _1120_ _1127_ _1128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_19_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5953__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7667_ _3451_ _3497_ _3509_ _0291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4879_ _1017_ net47 _1059_ _1060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_9406_ _0416_ clknet_leaf_36_i_clk core_0.execute.rf.reg_outputs\[5\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_34_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6618_ net212 _1829_ _2483_ _2558_ _2559_ _2560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__6902__A1 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7598_ core_0.execute.rf.reg_outputs\[15\]\[13\] _3429_ _3467_ _3468_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5705__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9337_ _0347_ clknet_leaf_5_i_clk core_0.execute.rf.reg_outputs\[9\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6549_ _2490_ _2438_ _2491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_104_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9268_ _0278_ clknet_leaf_7_i_clk core_0.execute.rf.reg_outputs\[14\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Right_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_167_2512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8219_ _2341_ _3833_ _3842_ _3843_ _3844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_246_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9199_ _0210_ clknet_leaf_56_i_clk core_0.ew_data\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8407__A1 _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4692__A2 _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6969__A1 _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7630__A2 _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_214_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_92_Right_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_2652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_133_Right_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_182_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__A2 net322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7146__A1 _1766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8894__A1 _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7697__A2 _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7449__A2 _3120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8646__A1 _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__S _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_209_3018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_2781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__A2 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8556__C _2136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4683__A2 net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_2039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_221_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7621__A2 _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5920_ _1904_ _1909_ _1910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_204_2962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7188__B _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5851_ net313 net206 _1840_ _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_152_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_201_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5235__I1 core_0.ew_data\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ core_0.ew_reg_ie\[0\] _0963_ _0966_ core_0.ew_reg_ie\[2\] _0948_ core_0.ew_reg_ie\[3\]
+ _0983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XPHY_EDGE_ROW_100_Right_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_172_Left_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_8570_ _1163_ _4133_ _4149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5396__B1 _1494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ _1771_ _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_233_3303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5935__A2 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_233_3314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7521_ core_0.execute.rf.reg_outputs\[15\]\[0\] _3403_ _2404_ _3404_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4733_ core_0.execute.pc_high_out\[6\] _0901_ _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__8798__I _4326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7916__B _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7452_ net116 _2419_ _3359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8885__A1 core_0.execute.pc_high_buff_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7688__A2 _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4664_ core_0.execute.rf.reg_outputs\[14\]\[3\] net262 net302 core_0.execute.rf.reg_outputs\[1\]\[3\]
+ _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_4_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_2324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6403_ _2206_ _2376_ _2217_ _2377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7383_ _1684_ _3301_ _3302_ _3303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4595_ _0783_ _0784_ _0785_ _0786_ _0787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_24_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9122_ _0134_ clknet_leaf_108_i_clk core_0.execute.sreg_priv_control.o_d\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6334_ _1546_ _2311_ _2312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_228_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9053_ _0079_ clknet_leaf_84_i_clk core_0.fetch.prev_request_pc\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7651__B _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_181_Left_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6265_ _1547_ _2240_ _2250_ _2251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6112__A2 _1772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8004_ _3647_ _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5216_ _1353_ net147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_244_3443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7860__A2 _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6196_ core_0.execute.alu_mul_div.div_cur\[7\] _2185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5871__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_235_Right_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_149_2297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5147_ _1267_ _1296_ _1299_ _1300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_rebuffer92_I _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7612__A2 _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_2453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5078_ core_0.decode.i_instr_l\[2\] _1235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input15_I i_core_int_sreg[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_223_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5623__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5474__I1 net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8906_ _4415_ _0624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_196_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_190_Left_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_8837_ _4316_ _4361_ _0609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5397__I _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8768_ core_0.execute.sreg_scratch.o_d\[10\] _4300_ _4308_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5926__A2 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7826__B _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7128__A1 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7719_ _3512_ _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_212_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8699_ _4219_ _4122_ _4260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8876__A1 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7679__A2 _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5154__A3 _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7117__I _2768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8628__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output83_I net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__A2 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5860__I net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7851__A2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_234_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4665__A2 net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A1 _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_202_Right_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8800__A1 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7603__A2 _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5614__A1 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__I1 net59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7367__A1 _2979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9429__CLK clknet_leaf_144_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5917__A2 _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7736__B _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8867__A1 _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9579__CLK clknet_leaf_21_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_215_3088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8619__A1 _2816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8095__A2 _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6050_ _2039_ _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7842__A2 _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I i_core_int_sreg[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _1145_ _1154_ _1177_ _1178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_72_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A2 _0673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5853__A1 net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5605__A1 _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6952_ _2711_ _2882_ _2883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ _1878_ _1879_ _1881_ _1892_ _1893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_88_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6883_ _2337_ _2755_ _2759_ net282 _2815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ core_0.execute.rf.reg_outputs\[2\]\[15\] _1797_ _1781_ core_0.execute.rf.reg_outputs\[10\]\[15\]
+ _1824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8622_ _4165_ _4194_ _4195_ _4196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5010__I net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6030__A1 core_0.execute.rf.reg_outputs\[11\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8553_ _1175_ _4126_ _1170_ _4134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5765_ net313 net177 _1755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__6581__A2 _2521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7504_ _3381_ _3387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_8
X_4716_ net19 net18 core_0.execute.irq_en _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8858__A1 core_0.execute.pc_high_buff_out\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8484_ net244 _4048_ _2923_ _2133_ _2895_ _4074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__7365__C _3073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5696_ _1700_ _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_20_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7435_ _2839_ _2821_ _3350_ _0218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4647_ _0831_ _0832_ _0833_ _0834_ _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__7530__A1 net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout2 _1746_ net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__5541__B1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7366_ _1885_ _3283_ _2423_ _1880_ _3285_ _3286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4578_ core_0.execute.rf.reg_outputs\[2\]\[10\] _0672_ _0707_ core_0.execute.rf.reg_outputs\[13\]\[10\]
+ _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4895__A2 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6776__I _2708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9105_ _0008_ clknet_leaf_113_i_clk core_0.execute.alu_mul_div.i_div vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6317_ core_0.execute.alu_mul_div.div_cur\[9\] _2220_ _2295_ _2296_ _2256_ _2297_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__8086__A2 _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5680__I _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7297_ _2564_ _2900_ _3218_ _1768_ _3219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_229_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6097__A1 core_0.execute.rf.reg_outputs\[3\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_9036_ _0063_ clknet_leaf_87_i_clk core_0.fetch.out_buffer_data_instr\[24\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7833__A2 _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ core_0.execute.alu_mul_div.div_cur\[1\] _2220_ _2235_ _2236_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_216_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5844__A1 _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6179_ core_0.execute.alu_mul_div.div_cur\[7\] net342 _2168_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8010__A2 _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_175_2611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8849__A1 _4335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_97_1679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_123_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8077__A2 _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_2740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6088__A1 core_0.execute.rf.reg_outputs\[9\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7824__A2 _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A2 net303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_235_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9251__CLK clknet_leaf_7_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_201_2921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_48_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8537__B1 _3192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_2__f_i_clk_I clknet_3_1_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8001__A2 _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_217_3117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_197_2880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8552__A3 net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5366__A3 _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5550_ _1597_ _1604_ _0079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4574__A1 core_0.execute.rf.reg_outputs\[5\]\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4501_ net326 net291 _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_14_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5481_ _1565_ _0049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_170_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7220_ net247 _1942_ _3144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7151_ _2004_ _3069_ _3075_ _3076_ _3077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_21_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8068__A2 _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6079__A1 net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_3246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6102_ core_0.execute.rf.reg_outputs\[12\]\[2\] _1819_ _1961_ _2092_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7082_ core_0.ew_data\[6\] _2642_ _3010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_241_3402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5826__B2 core_0.execute.rf.reg_outputs\[9\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6033_ core_0.execute.rf.reg_outputs\[6\]\[4\] net219 _1787_ core_0.execute.rf.reg_outputs\[3\]\[4\]
+ _2023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5005__I _1057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6094__A4 _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7028__B1 _2768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7579__B2 net36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer12 _1837_ net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_240_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer23 _0836_ net251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_206_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer34 _1848_ net319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7984_ core_0.execute.rf.reg_outputs\[5\]\[15\] _3671_ _3689_ _3692_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xrebuffer45 core_0.dec_r_reg_sel\[1\] net273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5054__A2 _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer56 _1759_ net325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6251__A1 core_0.execute.alu_mul_div.div_cur\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer67 net294 net295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6935_ _1894_ _2865_ _2866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_76_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer78 _1775_ net331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_25_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer89 _1796_ net336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_138_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_3375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_239_3386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6866_ _2449_ _2792_ _2798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_159_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6003__A1 core_0.execute.rf.reg_outputs\[1\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8605_ _1974_ _4179_ _4180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7376__B _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5817_ core_0.execute.rf.reg_outputs\[15\]\[0\] _1807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6797_ _1882_ _1925_ _2730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9585_ _0595_ clknet_leaf_108_i_clk core_0.execute.sreg_scratch.o_d\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_174_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6554__A2 _2349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8536_ _4053_ _4118_ _4119_ _4051_ _0550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5748_ _1400_ _1737_ _1738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xrebuffer102 _2528_ net349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4565__B2 core_0.execute.rf.reg_outputs\[13\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_2396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7503__A1 net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5679_ _1683_ _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8467_ _2389_ _2384_ _2391_ _4059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_170_2552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7418_ core_0.execute.sreg_priv_control.o_d\[15\] _1693_ _2996_ net7 _2689_ _3337_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_60_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9124__CLK clknet_leaf_108_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8398_ _4001_ _3996_ _4007_ _4009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7349_ _3263_ _3268_ _3201_ _3232_ _3270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__8059__A2 _3714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output169_I net169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8000__B _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7806__A2 _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9274__CLK clknet_leaf_155_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4955__S _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9019_ _0046_ clknet_leaf_80_i_clk core_0.fetch.out_buffer_data_instr\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_244_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_181_2681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5045__A2 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6242__A1 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7990__A1 _3401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire218_I _2025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clone6_A2 net246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_165_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6545__A2 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A1 core_0.execute.rf.reg_outputs\[6\]\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8298__A2 _3866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_212_3058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4859__A2 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__I core_0.fetch.prev_request_pc\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput81 net81 dbg_pc[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5808__A1 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput92 net92 dbg_r0[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_37_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__A1 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_1804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4492__B1 _0686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_223_3187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6084__I1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ net77 _1085_ _1161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_188_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7981__A1 _3465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6720_ net135 _2642_ _2657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5992__B1 _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6651_ _2588_ _2592_ _2593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Left_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_rebuffer5_I net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5602_ _1632_ _1634_ _0101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6582_ _2523_ _2522_ _2524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_9370_ _0380_ clknet_leaf_0_i_clk core_0.execute.rf.reg_outputs\[7\]\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_26_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5533_ _1082_ _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8321_ net213 _3827_ _3936_ _3937_ _3938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_119_1944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8252_ _3871_ _3873_ _3874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5464_ _1550_ _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7203_ _3093_ _3126_ _2710_ _3128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8183_ _1543_ net261 _3808_ _1545_ _3809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_100_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5395_ _0663_ _1486_ _1499_ _1497_ _0028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6259__C _2229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7134_ _2074_ _2562_ _3060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_0_226_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7065_ _2992_ _1314_ _2128_ _2993_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_clone75_I _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6016_ _1749_ _2005_ _2006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5275__A2 _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4483__B1 _0680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8213__A2 core_0.execute.alu_mul_div.mul_res\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7967_ core_0.execute.rf.reg_outputs\[5\]\[7\] _3679_ _3677_ _3683_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_3_3_0_i_clk clknet_0_i_clk clknet_3_3_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7972__A1 _3453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_2425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6918_ _2444_ _2449_ _2450_ _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4786__B2 core_0.ew_reg_ie\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7898_ _3457_ _3629_ _3642_ _0389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9637_ _0647_ clknet_leaf_96_i_clk net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6849_ _2776_ _2779_ _2781_ _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6527__A2 _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__A1 core_0.execute.rf.reg_outputs\[5\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__B2 core_0.execute.rf.reg_outputs\[4\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5735__B1 _1727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9568_ _0578_ clknet_leaf_21_i_clk core_0.execute.sreg_jtr_buff.o_d\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8519_ _0801_ _4048_ _3086_ _4104_ _4105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_9499_ _0509_ clknet_leaf_125_i_clk core_0.execute.alu_mul_div.mul_res\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_94_1638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_229_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_217_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_2710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6463__A1 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_6__f_i_clk clknet_3_3_0_i_clk clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_213_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_197_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6766__A2 _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7963__A1 core_0.execute.rf.reg_outputs\[5\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5974__B1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__B _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7715__A1 core_0.execute.rf.reg_outputs\[12\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6518__A2 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4529__B2 core_0.execute.rf.reg_outputs\[9\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5726__B1 _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7191__A2 core_0.execute.alu_mul_div.mul_res\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer3 net199 net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8140__A1 _3401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8691__A2 _4210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4701__A1 core_0.execute.rf.reg_outputs\[9\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5180_ core_0.decode.oc_alu_mode\[12\] _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_114_1885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_225_3216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5257__A2 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_2226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_147_Right_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_223_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8870_ _4386_ _4389_ _4390_ _0613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_207_2993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_69_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A2 _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6206__A1 core_0.execute.alu_mul_div.div_cur\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7821_ _3454_ _3585_ _3598_ _0356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7954__A1 _3408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4768__A1 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4964_ _1080_ _1143_ _1074_ _1140_ _1144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_2
X_7752_ _3463_ _3543_ _3558_ _0327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_80_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6703_ _2421_ _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_175_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_236_3345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4895_ _1072_ _1073_ _1075_ _1076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7683_ _3473_ _3498_ _3518_ _0298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6509__A2 _2349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7706__A1 _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9422_ _0432_ clknet_leaf_22_i_clk core_0.execute.rf.reg_outputs\[4\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_15_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6634_ _2571_ _2575_ _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5717__B1 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7182__A2 _2758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_2355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9353_ _0363_ clknet_leaf_5_i_clk core_0.execute.rf.reg_outputs\[8\]\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6565_ _2008_ _2337_ _2507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_154_2366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4997__C _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8304_ _3919_ _3921_ _3802_ _3922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5516_ net55 _1556_ _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9284_ _0294_ clknet_leaf_6_i_clk core_0.execute.rf.reg_outputs\[13\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6496_ net214 _1843_ _2438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__8131__A1 _3465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5447_ _1541_ _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8235_ _3853_ _3857_ _3828_ _3858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_219_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8682__A2 _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__A2 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Left_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5378_ _1464_ _1485_ _0025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8166_ _3462_ _3781_ _3796_ _0503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input45_I i_req_data[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7117_ _2768_ _3044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_238_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8097_ core_0.execute.rf.reg_outputs\[2\]\[15\] _3736_ _3756_ _3757_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8434__A2 _4031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7048_ _1292_ _2974_ _2975_ _2976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_165_2495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_114_Right_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8198__A1 _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9312__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4471__A3 _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7945__A1 _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8999_ _0026_ clknet_leaf_133_i_clk core_0.dec_r_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6748__A2 _1405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output201_I net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_Left_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5956__B1 _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5708__B1 _1709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8370__A1 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6920__A2 _2349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4479__I net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Left_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8189__A1 _1674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_220_3157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Left_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5947__B1 _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_123_i_clk clknet_4_5__leaf_i_clk clknet_leaf_123_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5411__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ core_0.execute.rf.reg_outputs\[11\]\[2\] _0680_ net341 core_0.execute.rf.reg_outputs\[3\]\[2\]
+ _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_83_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6911__A2 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_138_i_clk clknet_4_1__leaf_i_clk clknet_leaf_138_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_116_1903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6350_ _2221_ _2325_ _2326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_94_Left_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_231_3286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8113__A1 core_0.execute.rf.reg_outputs\[1\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ _1419_ net191 _1420_ _1421_ _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XPHY_EDGE_ROW_216_Right_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6281_ _2258_ _2265_ _0149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_121_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5232_ _1361_ net140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8020_ _3469_ _3695_ _3712_ _0441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6818__B _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5163_ core_0.execute.alu_mul_div.i_div _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_236_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_223_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5094_ _1250_ _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8922_ _4424_ _1322_ _4425_ _1507_ _4426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_223_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8853_ _4316_ _4375_ _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_182_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8324__I _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7804_ core_0.execute.rf.reg_outputs\[9\]\[2\] _3586_ _3580_ _3589_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8784_ _0899_ _4317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5996_ _1772_ _1980_ _1985_ _1986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_93_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_96_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7735_ _3428_ _3542_ _3549_ _0319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4947_ core_0.fetch.prev_request_pc\[7\] _1029_ _1126_ _1127_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_176_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7666_ core_0.execute.rf.reg_outputs\[13\]\[8\] _3504_ _3500_ _3509_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4878_ _0892_ _1058_ _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9405_ _0415_ clknet_leaf_49_i_clk core_0.execute.rf.reg_outputs\[5\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_6_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6617_ _2143_ _1973_ _2556_ _2559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_62_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__I net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7597_ _1430_ _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_171_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4913__A1 core_0.fetch.prev_request_pc\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9336_ _0346_ clknet_leaf_148_i_clk core_0.execute.rf.reg_outputs\[10\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6548_ _1851_ _2040_ _2490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8104__A1 core_0.execute.rf.reg_outputs\[1\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9267_ _0277_ clknet_leaf_10_i_clk core_0.execute.rf.reg_outputs\[14\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6479_ _2418_ _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6666__A1 _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8218_ _3834_ _3841_ _3802_ _3843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_167_2513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9198_ _0209_ clknet_leaf_51_i_clk core_0.ew_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4677__B1 net321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_246_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8407__A2 _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8149_ net97 _3787_ _3785_ _3788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_215_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__I _2008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8662__C _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_i_clk clknet_4_10__leaf_i_clk clknet_leaf_40_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8966__I0 net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4762__I core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8591__A1 _4154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_2653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4601__B1 net316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_55_i_clk clknet_4_11__leaf_i_clk clknet_leaf_55_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8343__A1 core_0.execute.alu_mul_div.mul_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6657__A1 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_209_3019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_2782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4668__B1 _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7082__A1 core_0.ew_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_204_2963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7909__A1 core_0.execute.rf.reg_outputs\[7\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_118_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5850_ core_0.dec_r_bus_imm _1839_ _1840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_201_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7385__A2 _3303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_201_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4801_ core_0.ew_reg_ie\[1\] _0964_ _0982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5396__A1 core_0.decode.i_imm_pass\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5396__B2 core_0.decode.i_instr_l\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5781_ _1770_ _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_233_3304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7520_ _3396_ _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_61_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4732_ core_0.execute.prev_pc_high\[4\] _0913_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_232_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8334__A1 core_0.execute.alu_mul_div.mul_res\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_138_2169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5148__A1 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7451_ _2616_ _3155_ _3358_ _0226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4663_ core_0.execute.rf.reg_outputs\[3\]\[3\] _0698_ net321 core_0.execute.rf.reg_outputs\[12\]\[3\]
+ _0849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_160_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8885__A2 _4385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6896__A1 _2694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _2221_ _2174_ _2376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_151_2325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7382_ _1684_ core_0.execute.sreg_irq_pc.o_d\[14\] _3302_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4594_ core_0.execute.rf.reg_outputs\[2\]\[9\] _0672_ _0715_ _0786_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_77_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_9121_ _0133_ clknet_leaf_64_i_clk core_0.execute.sreg_priv_control.o_d\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6333_ _2153_ _2310_ _2311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_51_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8637__A2 _4202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6648__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8747__C _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9052_ _0078_ clknet_leaf_84_i_clk core_0.fetch.prev_request_pc\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6264_ _1546_ _2249_ _2250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5215_ core_0.ew_data\[3\] net156 _1353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_177_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8003_ _3440_ _3694_ _3703_ _0433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6195_ _2181_ _2182_ _2183_ _2184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_244_3444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5871__A2 _1855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5146_ _1232_ _1297_ _1298_ _1269_ _1299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_149_2298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_208_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7073__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7073__B2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _1232_ _1233_ _1234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_162_2454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_rebuffer85_I net331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6820__A1 _1309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8905_ core_0.dec_mem_width _1251_ _1293_ _4414_ _4415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6820__B2 _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__I _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8948__I0 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8836_ core_0.execute.pc_high_out\[4\] _4327_ _4360_ _4361_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7376__A2 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8767_ _0789_ _4294_ _4306_ _4307_ _0593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_136_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5979_ core_0.execute.rf.reg_outputs\[2\]\[14\] _1797_ _1781_ core_0.execute.rf.reg_outputs\[10\]\[14\]
+ _1969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7718_ _3470_ _3521_ _3538_ _0313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_212_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8698_ _4258_ _4259_ _1435_ _0572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_192_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output199_I net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7649_ _3402_ _3497_ _3499_ _0283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8876__A2 _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9500__CLK clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9319_ _0329_ clknet_leaf_148_i_clk core_0.execute.rf.reg_outputs\[11\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7842__B _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8628__A2 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6639__A1 _1769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8657__C _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output76_I net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7300__A2 _3220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5862__A2 net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8673__B _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8800__A2 _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6811__A1 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5614__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8564__A1 _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7367__A2 _3069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__A1 _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8316__A1 _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8867__A2 _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_215_3089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6878__A1 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5550__A1 _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8619__A2 _2868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8567__C _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_44_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5302__A1 net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5000_ core_0.fetch.prev_request_pc\[12\] _1153_ _1177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_72_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A2 net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7055__A1 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6802__A1 _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__A2 net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6951_ _2833_ _2881_ _2882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_178_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ _1285_ _1883_ _1884_ _1885_ _1891_ _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_48_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6882_ _2813_ _2586_ _2814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8555__A1 _4080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5369__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8621_ net243 _4165_ _4167_ _4195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7927__B _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5833_ core_0.execute.rf.reg_outputs\[5\]\[15\] _1785_ _1802_ core_0.execute.rf.reg_outputs\[14\]\[15\]
+ _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_76_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6030__A2 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8552_ net75 net74 net73 _4121_ _4133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_29_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8307__A1 _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5764_ core_0.dec_r_bus_imm _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_118_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7503_ net20 _3381_ _3386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4715_ net37 core_0.execute.sreg_irq_flags.i_d\[2\] _0897_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8483_ _4039_ _4072_ _4073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4592__A2 _0685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5695_ _1699_ _1697_ _1700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_20_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6869__A1 _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7434_ net122 _3168_ _3350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4646_ core_0.execute.rf.reg_outputs\[1\]\[5\] net302 net321 core_0.execute.rf.reg_outputs\[12\]\[5\]
+ _0834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_25_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7662__B _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5541__A1 core_0.fetch.prev_request_pc\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7365_ _2370_ _3072_ _3284_ _2143_ _3073_ _3285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4577_ _0766_ _0767_ _0768_ _0769_ _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_114_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5541__B2 net169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9104_ _0007_ clknet_leaf_130_i_clk core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6316_ _1547_ _2288_ _2246_ _2296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_97_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7296_ _3216_ _3217_ _2564_ _3218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_228_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A2 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9035_ _0062_ clknet_leaf_87_i_clk core_0.fetch.out_buffer_data_instr\[23\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_31_Left_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6247_ _1547_ _2222_ _2234_ _2224_ _2235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_244_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__A2 net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6178_ core_0.execute.alu_mul_div.div_cur\[6\] _1843_ _2167_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7046__A1 _2438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5129_ _1259_ _1267_ _1277_ _1283_ _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_99_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8794__A1 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4804__B1 _0960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7061__A4 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output114_I net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7349__A2 _3268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8546__A1 _4080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8819_ _4324_ _4345_ _4346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7837__B _3595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_2612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5780__A1 _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8668__B _4201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7521__A2 _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7572__B _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7291__C _3073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_2741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7285__A1 _2468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6088__A2 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7798__I _3584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7037__A1 core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8785__A1 core_0.execute.sreg_irq_flags.o_d\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5599__A1 core_0.decode.i_instr_l\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_201_2922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8537__A1 _0765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8537__B2 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7747__B _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_217_3118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5771__A1 _1749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4574__A2 net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4500_ _0697_ _0698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5480_ core_0.fetch.out_buffer_data_instr\[9\] net68 _1559_ _1565_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_1 _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5781__I _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7150_ _1880_ _2456_ _3076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6101_ _1899_ _2090_ _2091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6079__A2 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_3247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7081_ _2709_ _3007_ _3008_ _3009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_225_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5826__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6032_ core_0.execute.rf.reg_outputs\[9\]\[4\] net224 _1818_ core_0.execute.rf.reg_outputs\[12\]\[4\]
+ _2022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_241_3403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__B2 core_0.execute.sreg_scratch.o_d\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_2268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7579__A2 core_0.ew_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8776__A1 _1726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer13 net240 net241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer24 net251 net252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7983_ _3469_ _3673_ _3691_ _0425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xrebuffer35 _0662_ net263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_178_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer46 net273 net274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6251__A2 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer57 _0707_ net285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6934_ _2011_ _2861_ _2864_ _2865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer68 _1835_ net327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XTAP_TAPCELL_ROW_25_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer79 _0777_ net307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_25_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8760__C _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6561__B _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6865_ _1338_ _2337_ _1285_ _2797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_239_3376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7200__A1 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6003__A2 _1779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8604_ _1292_ _3311_ _3329_ _4179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5816_ _0942_ _0943_ _0957_ _0955_ _1806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_9584_ _0594_ clknet_leaf_108_i_clk core_0.execute.sreg_scratch.o_d\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6796_ _1894_ _2728_ _2729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7751__A2 _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8535_ net72 _4053_ _4119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5762__A1 _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4565__A2 _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5747_ core_0.dec_jump_cond_code\[4\] _1394_ core_0.dec_pc_inc _1737_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_161_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_2397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8466_ net79 net78 _1226_ _4058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5678_ _1401_ _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_60_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7503__A2 _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8700__A1 net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_2553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7417_ core_0.execute.sreg_irq_pc.o_d\[15\] _3042_ _3044_ core_0.execute.sreg_scratch.o_d\[15\]
+ _3336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4629_ _0814_ _0815_ _0816_ _0817_ _0818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8397_ _4001_ _3996_ _4007_ _4008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_103_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7348_ _3263_ _3268_ _3269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7267__A1 _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9419__CLK clknet_leaf_136_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7279_ _3163_ _3199_ _3202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_244_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8935__C _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9018_ _0045_ clknet_leaf_80_i_clk core_0.fetch.out_buffer_data_instr\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_229_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_218_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_216_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_216_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8767__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_2682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8519__A1 _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7990__A2 _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7742__A2 _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4556__A2 _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_212_3059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4859__A3 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_128_Right_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_2069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7258__A1 _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput71 net71 dbg_pc[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_56_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput82 net82 dbg_pc[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput93 net93 dbg_r0[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_208_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__A2 _2370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4492__A1 core_0.execute.rf.reg_outputs\[7\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_108_1805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8758__A1 _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4492__B2 core_0.execute.rf.reg_outputs\[14\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_223_3188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7430__A1 _2130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4980_ _1146_ _1157_ _1159_ _1160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_203_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7981__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5992__A1 core_0.execute.rf.reg_outputs\[5\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5992__B2 core_0.execute.rf.reg_outputs\[14\]\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6650_ net283 _2591_ _2592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_73_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_171_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8930__A1 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5601_ _1591_ net41 _1369_ _1633_ _1634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_80_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6581_ net320 _2521_ _2457_ _2523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8320_ _3927_ _3935_ _3828_ _3937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5532_ core_0.fetch.prev_request_pc\[0\] _1078_ _1081_ _1594_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_30_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_1945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8251_ _3822_ _3872_ _3873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5463_ _1012_ _1551_ _1555_ _0041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7202_ _3093_ _3126_ _3127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_111_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8182_ _1542_ _2428_ _3808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5394_ core_0.decode.i_imm_pass\[2\] _1488_ _1494_ core_0.decode.i_instr_l\[13\]
+ _1495_ _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_10_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7940__B _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7133_ _3057_ _2456_ _3058_ _3059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_226_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7064_ core_0.execute.alu_mul_div.div_res\[6\] _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_105_Left_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6015_ core_0.decode.oc_alu_mode\[1\] _1328_ _2005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_214_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8749__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4483__B2 core_0.execute.rf.reg_outputs\[11\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clone68_I _0682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7421__A1 _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7966_ _3440_ _3672_ _3682_ _0417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8490__C _4047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7972__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6917_ _2845_ _2508_ _2847_ _2848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_159_2415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_2426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7897_ core_0.execute.rf.reg_outputs\[7\]\[10\] _3634_ _3636_ _3642_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9636_ _0646_ clknet_leaf_95_i_clk net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6848_ core_0.execute.sreg_data_page _1692_ _2780_ net8 core_0.dec_sreg_jal_over
+ _2781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_49_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8921__A1 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_114_Left_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4538__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5735__A1 core_0.execute.sreg_priv_control.o_d\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_9567_ _0577_ clknet_leaf_70_i_clk core_0.execute.sreg_irq_pc.o_d\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6779_ core_0.execute.alu_mul_div.div_res\[1\] _2712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5735__B2 _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8518_ _4080_ _3085_ _4104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9498_ _0508_ clknet_leaf_125_i_clk core_0.execute.alu_mul_div.mul_res\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_33_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output181_I net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9241__CLK clknet_leaf_2_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8449_ _2389_ _1226_ _4042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8011__B _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_183_2711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_123_Left_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_245_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__A2 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4474__A1 _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7412__A1 _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6215__A2 _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7963__A2 _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5974__A1 core_0.execute.rf.reg_outputs\[13\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5974__B2 core_0.execute.rf.reg_outputs\[9\]\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_194_2840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7715__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8912__A1 _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4529__A2 net347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5726__A1 core_0.execute.sreg_priv_control.o_d\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5726__B2 _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer4 net231 net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8140__A2 _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_239_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8279__I0 core_0.execute.alu_mul_div.mul_res\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4701__A2 _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_1886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8575__C _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8979__A1 _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_225_3217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7651__A1 core_0.execute.rf.reg_outputs\[13\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6454__A2 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_2227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_69_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7820_ core_0.execute.rf.reg_outputs\[9\]\[9\] _3591_ _3595_ _3598_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7954__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7751_ core_0.execute.rf.reg_outputs\[11\]\[12\] _3548_ _3554_ _3558_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_35_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4963_ _0895_ net48 _1142_ _1143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_59_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4768__A2 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6702_ _2637_ _2640_ _2641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_236_3346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7682_ core_0.execute.rf.reg_outputs\[13\]\[15\] _3496_ _3513_ _3518_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4894_ _1015_ _1074_ _1075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_74_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8903__A1 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7706__A2 _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9421_ _0431_ clknet_leaf_21_i_clk core_0.execute.rf.reg_outputs\[4\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6633_ _1863_ _2574_ _2575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_74_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5717__A1 core_0.execute.sreg_priv_control.o_d\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5717__B2 _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9352_ _0362_ clknet_leaf_152_i_clk core_0.execute.rf.reg_outputs\[9\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_171_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6390__A1 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6564_ _2341_ _2503_ _2504_ _2506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_116_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_2356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8303_ _3901_ _3909_ _3920_ _3921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_131_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5515_ _1047_ _1552_ _1584_ _0064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9283_ _0293_ clknet_leaf_7_i_clk core_0.execute.rf.reg_outputs\[13\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6495_ _2433_ _2436_ _2437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8131__A2 _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8234_ core_0.execute.alu_mul_div.mul_res\[3\] _3856_ _3857_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_42_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ core_0.execute.alu_mul_div.cbit\[0\] _1541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7670__B _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6693__A2 _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7890__A1 _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8165_ net90 _3787_ _3785_ _3796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_92_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5377_ core_0.dec_rf_ie\[15\] _1482_ _1468_ _1472_ _1485_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_227_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7116_ core_0.execute.sreg_irq_pc.o_d\[7\] _3042_ _2775_ core_0.execute.pc_high_out\[7\]
+ _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8096_ _3647_ _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_input38_I i_req_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6445__A2 _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7642__A1 _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7493__I1 core_0.ew_reg_ie\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ _2438_ _2973_ _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_198_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_165_2496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8198__A2 core_0.execute.alu_mul_div.cbit\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__A4 _0664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8998_ _0025_ clknet_leaf_127_i_clk core_0.dec_rf_ie\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7945__A2 _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6748__A3 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7949_ _3671_ _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_38_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5956__A1 core_0.execute.rf.reg_outputs\[13\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9619_ _0629_ clknet_leaf_109_i_clk core_0.dec_sreg_load vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_135_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5708__B2 _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__A2 _1031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8122__A2 _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7881__A1 core_0.execute.rf.reg_outputs\[7\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4695__A1 _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4495__I _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_232_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8189__A2 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_220_3147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_220_3158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7936__A2 _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7755__B _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5175__A2 _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6911__A3 _2756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4922__A2 _1016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_231_3287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_180_Right_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8113__A2 _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5300_ net188 net187 net190 net189 _1421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_24_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_114_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6280_ core_0.execute.alu_mul_div.div_cur\[5\] _2219_ _2264_ _2265_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_219_Left_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5231_ core_0.ew_data\[3\] core_0.ew_data\[11\] _1349_ _1361_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6675__A2 _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7872__A1 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ _1312_ _1313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_166_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6427__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7624__A1 core_0.execute.rf.reg_outputs\[14\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7475__I1 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5093_ _1249_ _1229_ _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_8921_ _1240_ _1302_ _4425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_235_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8852_ core_0.execute.pc_high_out\[6\] _4327_ _4374_ _4375_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_189_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_228_Left_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7927__A2 _3657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7803_ _3409_ _3585_ _3588_ _0348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8783_ _1249_ _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_176_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5938__A1 net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5995_ core_0.execute.rf.reg_outputs\[15\]\[13\] _0945_ _1821_ core_0.execute.rf.reg_outputs\[7\]\[13\]
+ _1984_ _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_148_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6060__B1 _1818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7734_ core_0.execute.rf.reg_outputs\[11\]\[4\] _3548_ _3539_ _3549_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4946_ _1091_ _1094_ _1122_ _1125_ _1126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_19_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A1 net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7665_ _3447_ _3497_ _3508_ _0290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4877_ core_0.fetch.out_buffer_data_instr\[19\] _1058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_191_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9404_ _0414_ clknet_leaf_36_i_clk core_0.execute.rf.reg_outputs\[5\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_46_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6616_ _2555_ _2557_ _2558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_rebuffer30_I _1843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7596_ _3465_ _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_132_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9335_ _0345_ clknet_leaf_148_i_clk core_0.execute.rf.reg_outputs\[10\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6547_ _2439_ _2488_ _2489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4913__A2 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8104__A2 _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_237_Left_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6115__A1 core_0.execute.rf.reg_outputs\[12\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_9266_ _0276_ clknet_leaf_9_i_clk core_0.execute.rf.reg_outputs\[14\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6478_ _2420_ _0190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6666__A2 _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8217_ _3834_ _3841_ _3842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7863__A1 _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5429_ _1277_ _1524_ _1525_ _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
X_9197_ _0208_ clknet_leaf_53_i_clk core_0.ew_data\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_167_2514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4677__A1 core_0.execute.rf.reg_outputs\[1\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4677__B2 core_0.execute.rf.reg_outputs\[12\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8148_ _3779_ _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_246_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8079_ _3440_ _3737_ _3747_ _0465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_226_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_246_Left_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_214_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5229__I0 core_0.ew_data\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7379__B1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7918__A2 _3652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8040__A1 core_0.execute.rf.reg_outputs\[3\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_242_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_2643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8591__A2 _4164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_178_2654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_194_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_191_2810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5874__I _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7854__A1 _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_2783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A1 core_0.execute.rf.reg_outputs\[5\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_1845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7082__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5093__A1 _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_204_2964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7909__A2 _3627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8031__A1 core_0.execute.rf.reg_outputs\[3\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_40_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _0978_ _0979_ _0980_ _0981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6593__A1 _2155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5780_ _0963_ _0962_ _1770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__5396__A2 _1488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_1974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5640__I0 _1016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_233_3305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _0912_ net111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_185_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8334__A2 _3830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7450_ net130 _2419_ _3358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4662_ _0848_ net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_142_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6401_ _1537_ _2353_ _2374_ _2375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7381_ net76 _2995_ _3300_ _2893_ _3301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_151_2326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4593_ core_0.execute.rf.reg_outputs\[6\]\[9\] net223 _0699_ core_0.execute.rf.reg_outputs\[12\]\[9\]
+ _0785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_77_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9120_ _0132_ clknet_leaf_67_i_clk core_0.execute.sreg_priv_control.o_d\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8098__A1 _3472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6332_ _2307_ _2309_ _2310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9051_ _0077_ clknet_leaf_92_i_clk core_0.fetch.prev_request_pc\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7845__A1 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6263_ _2247_ _2248_ _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5225__S net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7504__I _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8002_ core_0.execute.rf.reg_outputs\[4\]\[6\] _3700_ _3689_ _3703_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5214_ _1352_ net146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6194_ core_0.execute.alu_mul_div.div_cur\[4\] _1749_ _2183_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_177_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_244_3445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5145_ _1243_ _1273_ _1298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__9452__CLK clknet_leaf_16_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7440__S _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7073__A2 _2995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8270__A1 _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5076_ core_0.decode.i_instr_l\[0\] _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XTAP_TAPCELL_ROW_162_2455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8904_ _1257_ _1305_ _1520_ _4414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_223_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7379__C _2689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8022__A1 _3472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8835_ net244 _4328_ _4326_ _4359_ _4360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_35_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6033__B1 _1787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8766_ _1249_ _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5978_ core_0.execute.rf.reg_outputs\[5\]\[14\] _1785_ _1802_ core_0.execute.rf.reg_outputs\[14\]\[14\]
+ _1968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7717_ core_0.execute.rf.reg_outputs\[12\]\[14\] _3519_ _3528_ _3538_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4929_ core_0.fetch.prev_request_pc\[4\] _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_176_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8697_ core_0.execute.sreg_irq_pc.o_d\[10\] _4202_ _4259_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5694__I _1417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7648_ core_0.execute.rf.reg_outputs\[13\]\[0\] _3498_ _3486_ _3499_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7579_ _3387_ core_0.ew_data\[9\] _3449_ net36 _3453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_15_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9318_ _0328_ clknet_leaf_154_i_clk core_0.execute.rf.reg_outputs\[11\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8089__A1 _3459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8628__A3 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6639__A2 _2580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9249_ _0259_ clknet_leaf_38_i_clk core_0.execute.rf.reg_outputs\[15\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_122_i_clk clknet_4_5__leaf_i_clk clknet_leaf_122_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_137_i_clk clknet_4_1__leaf_i_clk clknet_leaf_137_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_215_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6024__B1 net331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6575__A1 _2438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4586__B1 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8316__A2 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6327__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4889__A1 _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6649__B _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7827__A1 _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9475__CLK clknet_leaf_16_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_238_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5302__A2 net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8864__B _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5779__I _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6950_ _2874_ _2880_ _2881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_178_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5901_ _1889_ _1890_ _1812_ _1891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6881_ _2571_ _2581_ _2717_ _1865_ _2813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_159_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8555__A2 _3261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8620_ _4185_ _4189_ _4193_ _4194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_88_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ core_0.execute.rf.reg_outputs\[1\]\[15\] _1779_ _1804_ core_0.execute.rf.reg_outputs\[11\]\[15\]
+ _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5369__A2 core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_0_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6566__A1 _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8551_ _4053_ _4131_ _4132_ _1702_ _0552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_174_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6030__A3 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5763_ _1519_ net215 _1752_ _1753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__8104__B _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7502_ _0946_ _0199_ _3385_ _0250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4714_ net69 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8482_ _4041_ _4070_ _4071_ _4072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6318__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5694_ _1417_ _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_20_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7433_ _2839_ _2766_ _3349_ _0217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4645_ core_0.execute.rf.reg_outputs\[14\]\[5\] net262 net341 core_0.execute.rf.reg_outputs\[3\]\[5\]
+ _0833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_114_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8758__C _4287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7364_ _1338_ _1973_ _1285_ _3284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5541__A2 _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4576_ core_0.execute.rf.reg_outputs\[7\]\[10\] net297 _0697_ core_0.execute.rf.reg_outputs\[3\]\[10\]
+ _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_114_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9103_ _0006_ clknet_leaf_112_i_clk core_0.decode.oc_alu_mode\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_97_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4858__I _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6315_ _2221_ _2294_ _2295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7295_ _2568_ _2594_ _3217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9034_ _0061_ clknet_leaf_86_i_clk core_0.fetch.out_buffer_data_instr\[22\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_229_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8491__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6246_ _1546_ _2233_ _2234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6097__A3 _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ core_0.execute.alu_mul_div.div_cur\[7\] net342 _2166_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_54_i_clk clknet_4_11__leaf_i_clk clknet_leaf_54_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5128_ _1278_ _1282_ _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input20_I i_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6294__B _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8794__A2 _1738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5059_ _1086_ _1223_ _1224_ _1162_ net167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_196_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4804__A1 core_0.ew_reg_ie\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4804__B2 core_0.ew_reg_ie\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69_i_clk clknet_4_12__leaf_i_clk clknet_leaf_69_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_149_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8546__A2 _3225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8818_ _4335_ _4342_ _4343_ _4344_ _4345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_0_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_2613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8749_ net215 _4294_ _4297_ _4287_ _0585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_164_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_109_Right_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6309__A1 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_180_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5780__A2 _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7853__B _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_8_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7809__A1 core_0.execute.rf.reg_outputs\[9\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8482__A1 _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_186_2742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8684__B _4201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7037__A2 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8234__A1 core_0.execute.alu_mul_div.mul_res\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6796__A1 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5599__A2 _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9011__D _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_201_2923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8537__A2 _4048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6548__A1 _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_217_3119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_197_2882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5771__A2 _1760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_2 _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6100_ net96 _1813_ _2080_ _2089_ _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_10_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_228_3248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7080_ _2708_ net289 _3008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8473__A1 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5287__A1 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6031_ _2017_ _2018_ _2019_ _2020_ _2021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_67_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_241_3404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__A2 _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5039__A1 _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8776__A2 _4295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_169_Left_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xrebuffer14 net240 net242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6787__A1 _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7982_ core_0.execute.rf.reg_outputs\[5\]\[14\] _3671_ _3689_ _3691_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer25 _0836_ net253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer36 _1835_ net264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xrebuffer47 _0688_ net275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6933_ _2011_ _2863_ _2864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4798__B1 _0960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7938__B _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer58 net285 net286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_194_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer69 _0682_ net297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_25_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6539__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6864_ _2508_ _2794_ _2795_ _2796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_193_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_3377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7200__A2 core_0.execute.sreg_irq_pc.o_d\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8603_ _1326_ _2556_ _4178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5815_ core_0.execute.rf.reg_outputs\[12\]\[0\] _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_92_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9583_ _0593_ clknet_leaf_109_i_clk core_0.execute.sreg_scratch.o_d\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6795_ _2011_ _2719_ _2727_ _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5211__A1 core_0.ew_data\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8534_ _4115_ _4117_ _4118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5746_ _1420_ _1735_ _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_32_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5762__A2 net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_2398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8465_ _2133_ _2821_ _4056_ _4057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_178_Left_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5677_ _1672_ _1681_ _1682_ _0128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8700__A2 _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_2554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7416_ _0997_ _3333_ _3334_ _3335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_142_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4628_ core_0.execute.rf.reg_outputs\[7\]\[6\] net297 _0697_ core_0.execute.rf.reg_outputs\[3\]\[6\]
+ _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5514__A2 _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8396_ _4000_ _4006_ _4007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input68_I i_req_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7347_ _3264_ _3267_ _1403_ _3268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _0753_ net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_13_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8464__A1 _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7267__A2 core_0.execute.alu_mul_div.mul_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7278_ _3200_ _3201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_4_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5278__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9017_ _0044_ clknet_leaf_80_i_clk core_0.fetch.out_buffer_data_instr\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6229_ _2217_ _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_244_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_187_Left_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_244_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__B _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8009__B _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8767__A2 _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_181_2683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9170__CLK clknet_leaf_42_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8519__A2 _4048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_87_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5202__A1 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5053__I1 _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_196_Left_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8679__B _4201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4859__A4 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8455__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__A1 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput72 net72 dbg_pc[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_56_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput83 net83 dbg_pc[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_207_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput94 net94 dbg_r0[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5808__A3 _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9513__CLK clknet_leaf_122_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4492__A2 net296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8758__A2 _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_2900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_223_3189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8861__C _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7430__A2 _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_203_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_203_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_2199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5992__A2 _1785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8391__C2 _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5600_ _1591_ _1569_ _1633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6580_ net320 _2521_ _2457_ _2522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_TAPCELL_ROW_80_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6941__A1 _2871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8589__B _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5531_ _1593_ _0071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_1935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_119_1946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8250_ _3865_ _3870_ _3872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_124_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7497__A2 _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8694__A1 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ net48 _1554_ _1555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_200_Left_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7201_ _1683_ _3124_ _3125_ _3126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_111_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4704__B1 _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8181_ _1674_ _1875_ _2372_ _2076_ _1540_ _3807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_10_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5393_ _0668_ _1486_ _1498_ _1497_ _0027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_100_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7132_ _3057_ _2456_ _2480_ _3058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_238_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7063_ _1290_ _2989_ _2990_ _1742_ _2991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__5233__S _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7512__I _3394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6014_ _1751_ _1960_ _2003_ _2004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_94_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8749__A2 _4294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8771__C _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7668__B _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7965_ core_0.execute.rf.reg_outputs\[5\]\[6\] _3679_ _3677_ _3682_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5432__A1 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_109_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6916_ _2508_ _2846_ _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_rebuffer60_I _0825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_2416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7896_ _3454_ _3628_ _3641_ _0388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5983__A2 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_194_Right_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9635_ _0645_ clknet_leaf_98_i_clk net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_193_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7185__A1 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6847_ _2692_ _2693_ _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__7185__B2 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6778_ _2710_ _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9566_ _0576_ clknet_leaf_103_i_clk core_0.execute.sreg_irq_pc.o_d\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6932__A1 _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5735__A2 _1700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8517_ _4039_ _4102_ _4103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5729_ core_0.execute.sreg_priv_control.o_d\[11\] _1701_ _1723_ _1698_ _1724_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9497_ _0507_ clknet_leaf_121_i_clk core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_162_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8685__A1 _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8448_ _4040_ _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_60_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output174_I net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8379_ core_0.execute.alu_mul_div.mul_res\[13\] _3830_ _3992_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6160__A2 _1837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8437__A1 _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_183_2712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6999__A1 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7660__A2 _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5671__A1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4474__A2 net301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7412__A2 core_0.execute.alu_mul_div.mul_res\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7297__C _1768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5974__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_161_Right_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_194_2841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8912__A2 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6923__A1 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5726__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4934__B1 _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9066__CLK clknet_leaf_110_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xrebuffer5 net234 net233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8676__A1 core_0.execute.sreg_irq_pc.o_d\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_210_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5117__I _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8428__A1 _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_225_3207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_225_3218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7100__A1 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5053__S _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7651__A2 _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5662__A1 _1668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4892__S _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_143_2228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_207_2995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8600__A1 core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__B _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_110_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5414__A1 core_0.decode.i_instr_l\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__B2 core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4962_ _0895_ _1012_ _1142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_35_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7750_ _3460_ _3543_ _3557_ _0326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6701_ _2638_ _2639_ _2640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_47_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7681_ _3470_ _3498_ _3517_ _0297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7167__A1 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4893_ _1072_ _1073_ _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_236_3347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8903__A2 _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6632_ _2055_ _1926_ _1329_ _2574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_74_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9420_ _0430_ clknet_leaf_17_i_clk core_0.execute.rf.reg_outputs\[4\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5717__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9351_ _0361_ clknet_leaf_152_i_clk core_0.execute.rf.reg_outputs\[9\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6563_ _2503_ _2504_ _2341_ _2505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_42_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_2357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5514_ net54 _1556_ _1584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6411__I net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8302_ core_0.execute.alu_mul_div.mul_res\[7\] _3908_ _3920_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8667__A1 _4203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9282_ _0292_ clknet_leaf_9_i_clk core_0.execute.rf.reg_outputs\[13\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6494_ _2434_ _2435_ _2436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6678__B1 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7951__B _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8233_ _1535_ _3855_ _3856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_14_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5445_ _1539_ _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_112_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6142__A2 _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8419__A1 _2921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_35_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5350__B1 _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8164_ _3459_ _3781_ _3795_ _0502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7890__A2 _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ _1464_ _1484_ _0024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_112_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7115_ _2774_ _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_227_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8095_ _3469_ _3738_ _3755_ _0473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ _2438_ _2973_ _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7642__A2 _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5653__A1 _1662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_214_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_2497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8997_ _0024_ clknet_leaf_141_i_clk core_0.dec_rf_ie\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5405__A1 _1313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6748__A4 _2680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7948_ core_0.ew_reg_ie\[5\] _3394_ _3671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_49_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5956__A2 _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7879_ core_0.execute.rf.reg_outputs\[7\]\[2\] _3629_ _3621_ _3632_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9618_ _0628_ clknet_leaf_20_i_clk core_0.dec_sreg_store vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__6905__A1 _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5708__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4916__B1 _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4550__B _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9549_ _0559_ clknet_leaf_131_i_clk core_0.execute.alu_flag_reg.o_d\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_92_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8658__A1 _4212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output99_I net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7330__A1 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7330__B2 _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7881__A2 _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4776__I core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8830__A1 _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7633__A2 _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_230_Right_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_189_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_220_3148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7397__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_213_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5947__A2 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7149__A1 _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7149__B2 _1885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8897__A1 core_0.execute.pc_high_buff_out\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6372__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5175__A3 _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5048__S _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6231__I _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_25_Right_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_231_3288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__S _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7172__I1 _3097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5230_ _1360_ net139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7872__A2 _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5161_ _1232_ _1256_ _1270_ _1312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_224_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__A2 _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5092_ net70 _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5635__A1 _1057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8920_ _1267_ _1296_ _4424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_34_Right_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_223_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_142_Left_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_8851_ net288 _4328_ _4326_ _4373_ _4374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_182_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7388__A1 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7802_ core_0.execute.rf.reg_outputs\[9\]\[1\] _3586_ _3580_ _3588_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8782_ _2413_ _4315_ _0600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5310__I _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5994_ _1981_ _1982_ _1983_ _1984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5938__A2 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7946__B _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4945_ _1090_ _1099_ _1124_ _1125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7733_ _3541_ _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4610__A2 net324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8888__A1 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4876_ _0893_ net56 _1056_ _1057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7664_ core_0.execute.rf.reg_outputs\[13\]\[7\] _3504_ _3500_ _3508_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9381__CLK clknet_leaf_155_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9403_ _0413_ clknet_leaf_35_i_clk core_0.execute.rf.reg_outputs\[5\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_6_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ _2143_ _1973_ _2556_ _2557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7595_ _3387_ core_0.ew_data\[13\] _3449_ net25 _3465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XPHY_EDGE_ROW_43_Right_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7560__A1 net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__A2 _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6141__I _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9334_ _0344_ clknet_leaf_155_i_clk core_0.execute.rf.reg_outputs\[10\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6546_ net258 _2487_ _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_151_Left_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_rebuffer23_I _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6477_ core_0.dec_mem_we net158 _2419_ _2420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6115__A2 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9265_ _0275_ clknet_leaf_30_i_clk core_0.execute.rf.reg_outputs\[14\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8216_ _3839_ _3840_ _3841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5428_ _1241_ _1243_ _1316_ _1502_ _1525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_9196_ _0207_ clknet_leaf_76_i_clk core_0.ew_data\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7863__A2 _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input50_I i_req_data[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_2515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4677__A2 net302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5359_ _1464_ _1473_ _0018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8147_ _3420_ _3780_ _3786_ _0494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8812__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7615__A2 _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8078_ core_0.execute.rf.reg_outputs\[2\]\[6\] _3743_ _3745_ _3747_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_52_Right_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_226_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7029_ _2955_ _2956_ _2957_ _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_output137_I net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7379__A1 core_0.execute.sreg_priv_control.o_d\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7379__B2 net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8017__B _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8040__A2 _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5929__A2 _1801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6051__A1 _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_2644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4601__A2 _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8879__A1 _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_2800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7551__A1 core_0.execute.rf.reg_outputs\[15\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5562__B1 _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5890__I core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7303__A1 _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6657__A3 _1862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7854__A2 _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_2784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A1 net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4668__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Right_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_111_1846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8803__A1 _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7606__A2 _3396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5617__A1 core_0.decode.i_imm_pass\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7610__I _3475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5093__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_204_2965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8031__A2 _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5130__I core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A1 _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7766__B _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6593__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5640__I1 core_0.decode.i_imm_pass\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ core_0.execute.pc_high_out\[4\] net104 _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_56_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_233_3306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4661_ net97 net324 _0847_ _0848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_126_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6345__A2 _2218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6400_ _1540_ _2364_ _2369_ _2373_ _1536_ _2374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5553__B1 _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7380_ _3298_ _3299_ _3300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4592_ core_0.execute.rf.reg_outputs\[14\]\[9\] _0685_ net285 core_0.execute.rf.reg_outputs\[13\]\[9\]
+ _0784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_141_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_151_2327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6331_ core_0.execute.alu_mul_div.div_cur\[11\] net327 _2300_ _2293_ _2308_ _2309_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__8098__A2 _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5506__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9050_ _0076_ clknet_leaf_92_i_clk core_0.fetch.prev_request_pc\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6262_ _2207_ _2239_ _2180_ _2248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7845__A2 _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5856__A1 net314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ core_0.ew_data\[2\] net156 _1352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8001_ _3434_ _3694_ _3702_ _0432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_177_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6193_ core_0.execute.alu_mul_div.div_cur\[5\] _1851_ _2182_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_244_3435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_244_3446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5144_ _1241_ _1260_ _1266_ _1297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_208_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A1 _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8270__A2 _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ core_0.decode.i_instr_l\[1\] _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7520__I _3396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6281__A1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_2456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8903_ _1229_ _1305_ _4413_ _4307_ _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_223_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8834_ _4324_ _4358_ _4359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8022__A2 _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7676__B _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6033__B2 core_0.execute.rf.reg_outputs\[3\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8765_ core_0.execute.sreg_scratch.o_d\[9\] _4300_ _4306_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7781__A1 _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5977_ core_0.execute.rf.reg_outputs\[15\]\[14\] _0945_ _1821_ core_0.execute.rf.reg_outputs\[7\]\[14\]
+ _1967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_164_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7716_ _3466_ _3521_ _3537_ _0312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_212_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4928_ core_0.fetch.prev_request_pc\[4\] _1032_ _1034_ core_0.fetch.prev_request_pc\[5\]
+ _1108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5792__B1 _1781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8696_ _4249_ core_0.execute.mem_stage_pc\[10\] _4255_ _4257_ _4209_ _4258_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_19_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7647_ _3496_ _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_7_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4859_ _1032_ _1034_ _1037_ _1039_ _1040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_7_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6336__A2 _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7578_ _3397_ _3451_ _3452_ _0259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_105_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9317_ _0327_ clknet_leaf_1_i_clk core_0.execute.rf.reg_outputs\[11\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6529_ net235 _1999_ _2471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8089__A2 _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9248_ _0258_ clknet_leaf_37_i_clk core_0.execute.rf.reg_outputs\[15\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_219_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5847__A1 net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9179_ _0190_ clknet_leaf_44_i_clk net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_208_3010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8261__A2 _2349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4822__A2 core_0.ew_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8013__A2 _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6024__A1 core_0.execute.rf.reg_outputs\[13\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_195_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7772__A1 core_0.execute.rf.reg_outputs\[10\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5885__I _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__B2 core_0.execute.rf.reg_outputs\[9\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6327__A2 _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9009__D _0036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4889__A2 _1069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__I _3472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7827__A2 _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5838__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5302__A3 net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5900_ _1338_ _1883_ _1890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5861__I1 _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6880_ _2796_ _2800_ _2811_ _2812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_88_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6015__A1 core_0.decode.oc_alu_mode\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5831_ _1773_ _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_158_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5369__A3 core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7763__A1 _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8550_ net74 _4053_ _4132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_173_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5762_ _1519_ net184 _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6030__A4 _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7501_ net154 _0199_ _3385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4713_ _0894_ _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_29_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7515__A1 net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_4_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8481_ net81 _4040_ _4071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6318__A2 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5693_ _1697_ _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_44_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7432_ net115 _3168_ _3349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4644_ core_0.execute.rf.reg_outputs\[5\]\[5\] _0677_ net318 core_0.execute.rf.reg_outputs\[4\]\[5\]
+ _0832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_13_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7363_ _2143_ _2370_ _3283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4575_ core_0.execute.rf.reg_outputs\[4\]\[10\] _0719_ _0709_ core_0.execute.rf.reg_outputs\[8\]\[10\]
+ _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_12_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9102_ _0005_ clknet_leaf_112_i_clk core_0.decode.oc_alu_mode\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6314_ _2156_ _2293_ _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7294_ _2587_ _2577_ _3216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7818__A2 _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9033_ _0060_ clknet_leaf_87_i_clk core_0.fetch.out_buffer_data_instr\[21\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6245_ _2176_ _2232_ _2233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8491__A2 _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8774__C _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6176_ _2154_ _2164_ _2165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5127_ _1247_ _1281_ _1282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_207_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_rebuffer90_I _1798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Right_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6254__A1 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5058_ net78 _1085_ _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8790__B _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input13_I i_core_int_sreg[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8817_ core_0.execute.pc_high_buff_out\[2\] _4334_ _4344_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7754__A1 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_175_2614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8748_ core_0.execute.sreg_scratch.o_d\[1\] _4295_ _4297_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_165_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8679_ _4212_ core_0.execute.mem_stage_pc\[7\] _4201_ _4243_ _4244_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7506__A1 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5654__B _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_214_3080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7809__A2 _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output81_I net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_83_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_186_2743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6493__A1 net254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_201_2924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__A2 _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_1789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_213_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8170__A1 net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4959__I _1071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_3 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6720__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8473__A2 _4041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_3249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6030_ core_0.execute.rf.reg_outputs\[11\]\[4\] _0942_ _0947_ _0948_ _2020_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5287__A2 net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input5_I i_core_int_sreg[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_146_2259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5039__A2 _1149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6236__A1 _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_175_Right_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xrebuffer15 _0848_ net243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7981_ _3465_ _3673_ _3690_ _0424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_178_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__A2 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer26 _1745_ net254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_221_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer37 net264 net265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xrebuffer48 net349 net276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6932_ _1930_ _2722_ _2862_ _2863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4798__A1 core_0.ew_reg_ie\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5995__B1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4798__B2 core_0.ew_reg_ie\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer59 _1841_ net287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_25_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ core_0.decode.oc_alu_mode\[11\] _2795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_159_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8115__B _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6539__A2 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_239_3378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8602_ _1974_ _3330_ _4177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6414__I _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5814_ _1803_ _1804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_201_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9582_ _0592_ clknet_leaf_20_i_clk core_0.execute.sreg_scratch.o_d\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6794_ _2010_ _2726_ _2727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6944__C1 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5211__A2 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_121_i_clk clknet_4_5__leaf_i_clk clknet_leaf_121_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8533_ _2133_ _3155_ _4116_ _4046_ _4117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_17_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5745_ _1734_ _1394_ _1412_ _1403_ _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__7446__S _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8769__C _4307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_2399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4970__A1 core_0.fetch.prev_request_pc\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8464_ _1403_ core_0.execute.sreg_irq_pc.o_d\[2\] _2132_ _4055_ _4056_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_17_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5676_ _1537_ _1534_ _1682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8161__A1 net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7415_ core_0.execute.alu_mul_div.div_cur\[15\] _0997_ _3334_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_170_2555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4627_ core_0.execute.rf.reg_outputs\[4\]\[6\] _0719_ net316 core_0.execute.rf.reg_outputs\[8\]\[6\]
+ _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8395_ _1537_ _4004_ _4005_ _4006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_136_i_clk clknet_4_1__leaf_i_clk clknet_leaf_136_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_4_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7346_ _3265_ _3266_ _2673_ _3267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4558_ _0742_ _0716_ _0747_ _0752_ _0753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_12_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7277_ _3163_ _3199_ _3200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4489_ core_0.execute.rf.reg_outputs\[4\]\[15\] _0687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_217_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6475__A1 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9016_ _0043_ clknet_leaf_79_i_clk core_0.fetch.out_buffer_data_instr\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_218_17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _2141_ _2215_ _2216_ _2217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6159_ core_0.execute.alu_mul_div.div_cur\[13\] _1837_ _2148_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_232_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9112__D _0002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6227__A1 core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9315__CLK clknet_leaf_10_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_142_Right_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7975__A1 core_0.execute.rf.reg_outputs\[5\]\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_2684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5202__A2 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7864__B _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8152__A1 _3434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6702__A2 _2640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8695__B _4249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8455__A2 _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6466__A1 _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__A2 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput73 net73 dbg_pc[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_56_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput84 net84 dbg_pc[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__5808__A4 _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput95 net95 dbg_r0[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6218__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_1807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_199_2901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7966__A1 _3440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5977__B1 _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7718__A1 _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_224_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__B1 _1723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8391__A1 _1674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7194__A2 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8391__B2 _1973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7774__B _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6941__A2 _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5530_ core_0.decode.i_flush _1253_ _1008_ _1592_ _1593_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xclkbuf_leaf_53_i_clk clknet_4_11__leaf_i_clk clknet_leaf_53_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8143__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_1936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_11__f_i_clk clknet_3_5_0_i_clk clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5461_ _1550_ _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8694__A2 _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7200_ _1683_ core_0.execute.sreg_irq_pc.o_d\[9\] _3125_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8180_ _1543_ _2011_ _3805_ _1545_ _3806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4704__B2 core_0.execute.rf.reg_outputs\[10\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ core_0.decode.i_imm_pass\[1\] _1488_ _1494_ core_0.decode.i_instr_l\[12\]
+ _1495_ _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XPHY_EDGE_ROW_244_Right_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_99_Right_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7131_ _2432_ _2441_ _2455_ _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
Xclkbuf_leaf_68_i_clk clknet_4_12__leaf_i_clk clknet_leaf_68_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_239_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9338__CLK clknet_leaf_155_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7062_ _1743_ core_0.execute.alu_mul_div.mul_res\[6\] _2990_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6013_ _1751_ _2002_ _2003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5313__I _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_206_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Left_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7964_ _3434_ _3672_ _3681_ _0416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_38_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _2510_ _2509_ _2846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7895_ core_0.execute.rf.reg_outputs\[7\]\[9\] _3634_ _3636_ _3641_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4640__B1 net284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_2417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_31_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9634_ _0644_ clknet_leaf_95_i_clk net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_76_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6846_ core_0.execute.sreg_irq_flags.o_d\[1\] _2777_ _2778_ core_0.execute.trap_flag
+ _2779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_159_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8382__A1 core_0.execute.alu_mul_div.mul_res\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5196__A1 _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9565_ _0575_ clknet_leaf_81_i_clk core_0.execute.sreg_irq_pc.o_d\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6777_ core_0.dec_sreg_load _2673_ _2710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_18_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8516_ _4041_ _4100_ _4101_ _4102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4943__A1 core_0.fetch.prev_request_pc\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5728_ _0765_ _1699_ _1723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8134__A1 core_0.execute.rf.reg_outputs\[1\]\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_9496_ _0506_ clknet_leaf_18_i_clk net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_45_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8447_ _1371_ _1737_ _4040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XPHY_EDGE_ROW_28_Left_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5659_ _1543_ _1545_ _1667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_211_3050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5499__A2 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8378_ _1988_ _3833_ _3988_ _3990_ _3991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_102_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_211_Right_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output167_I net167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_1__f_i_clk_I clknet_3_0_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7329_ _2371_ _3072_ _3249_ net240 _3073_ _3250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_229_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_217_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_2713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_245_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5671__A2 _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Left_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7859__B _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7948__A1 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6620__A1 _2008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4631__B1 net286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8373__A1 _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_194_2842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5187__A1 _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5187__B2 _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4934__A1 core_0.fetch.prev_request_pc\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Left_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4934__B2 core_0.fetch.prev_request_pc\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8125__A1 _3456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer6 _1853_ net315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__8676__A2 _4209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6687__A1 _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4698__B1 net347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8428__A2 _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_225_3208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5111__A1 core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6229__I _2217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7769__B _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7939__A1 _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_207_2996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4961_ _1075_ _1138_ _1140_ _1141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_35_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6700_ core_0.execute.rf.reg_outputs\[7\]\[3\] _2611_ _2612_ core_0.execute.rf.reg_outputs\[5\]\[3\]
+ _2639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_129_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7680_ core_0.execute.rf.reg_outputs\[13\]\[14\] _3496_ _3513_ _3517_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4892_ net62 core_0.fetch.out_buffer_data_instr\[3\] _0894_ _1073_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7167__A2 _3091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8364__A1 _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_236_3348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6631_ _1769_ _2572_ _1863_ _2573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5178__A1 _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9350_ _0360_ clknet_leaf_152_i_clk core_0.execute.rf.reg_outputs\[9\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6562_ _1869_ _1873_ _1877_ _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__8116__A1 _3440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_2358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8301_ core_0.execute.alu_mul_div.mul_res\[8\] _3918_ _3919_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5513_ _1044_ _1552_ _1583_ _0063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9281_ _0291_ clknet_leaf_32_i_clk core_0.execute.rf.reg_outputs\[13\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6493_ net254 _2040_ _2435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6678__A1 core_0.execute.rf.reg_outputs\[7\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6678__B2 core_0.execute.rf.reg_outputs\[5\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8232_ core_0.execute.alu_mul_div.cbit\[2\] _3854_ _3855_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5444_ _1538_ _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_2_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4689__B1 net284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8163_ net89 _3787_ _3785_ _3795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5375_ core_0.dec_rf_ie\[14\] _1482_ _1466_ _1472_ _1484_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_227_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7114_ core_0.execute.sreg_priv_control.o_d\[7\] _1693_ _2996_ net14 _3041_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_227_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8094_ core_0.execute.rf.reg_outputs\[2\]\[14\] _3736_ _3745_ _3755_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5102__A1 _1257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7045_ _2902_ _2454_ _2437_ _2973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_242_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_2487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_2498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8996_ _0023_ clknet_leaf_140_i_clk core_0.dec_rf_ie\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_210_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7947_ _3473_ _3652_ _3670_ _0410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4613__B1 _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8355__A1 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7878_ _3409_ _3628_ _3631_ _0380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7158__A2 _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5169__A1 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9617_ _0627_ clknet_leaf_132_i_clk core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_42_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6829_ _2713_ _2761_ _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6905__A2 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4916__A1 core_0.fetch.prev_request_pc\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9548_ _0558_ clknet_leaf_134_i_clk core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__8107__A1 _3414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4916__B2 core_0.fetch.prev_request_pc\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6118__B1 _1797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9479_ _0489_ clknet_leaf_144_i_clk core_0.execute.rf.reg_outputs\[1\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6669__A1 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__A1 _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5644__A2 _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6841__A1 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7589__B _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_220_3149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7397__A2 _1974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8594__A1 net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4604__B1 _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8346__A1 core_0.execute.alu_mul_div.mul_res\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_54_Left_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8897__A2 _4386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4907__A1 core_0.fetch.prev_request_pc\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_181_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6109__B1 _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5580__A1 core_0.decode.i_instr_l\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_231_3289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4967__I core_0.fetch.prev_request_pc\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5332__A1 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5160_ _1253_ _1309_ _1229_ _1256_ _1311_ _0012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5091_ _1237_ _1240_ _1244_ _1247_ _1248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8821__A2 _4327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__A1 _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5635__A2 _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5798__I _1787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8850_ _4324_ _4372_ _4373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_189_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7801_ _3402_ _3585_ _3587_ _0347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5399__A1 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8781_ core_0.execute.irq_en net18 _4217_ core_0.execute.sreg_irq_flags.o_d\[0\]
+ _4315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_204_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5993_ core_0.execute.rf.reg_outputs\[2\]\[13\] _1797_ _1781_ core_0.execute.rf.reg_outputs\[10\]\[13\]
+ _1983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6060__A2 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7732_ _3421_ _3542_ _3547_ _0318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4944_ _1087_ _1102_ _1123_ _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_176_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8337__A1 _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7663_ _3441_ _3497_ _3507_ _0289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ _0893_ _1055_ _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8888__A2 _4387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5239__S _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6899__A1 _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9402_ _0412_ clknet_leaf_36_i_clk core_0.execute.rf.reg_outputs\[5\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_28_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6614_ net212 _1974_ _2556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_7594_ _3403_ _3463_ _3464_ _0263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9333_ _0343_ clknet_leaf_155_i_clk core_0.execute.rf.reg_outputs\[10\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6545_ _2484_ _1962_ _2485_ _2486_ _2487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_171_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7454__S _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9264_ _0274_ clknet_leaf_33_i_clk core_0.execute.rf.reg_outputs\[14\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6476_ _2418_ _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_rebuffer16_I _0848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8215_ _1679_ _3837_ core_0.execute.alu_mul_div.mul_res\[1\] _3840_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_112_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5323__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _1294_ _1269_ _1303_ _1305_ _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_112_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9195_ _0206_ clknet_leaf_55_i_clk core_0.ew_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_2_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_2516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8146_ net96 _3781_ _3785_ _3786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5358_ core_0.dec_rf_ie\[8\] _1438_ _1470_ _1472_ _1473_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_100_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input43_I i_req_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8812__A2 _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8077_ _3434_ _3737_ _3746_ _0464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5289_ net184 net177 _1409_ _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_215_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5626__A2 _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6823__A1 _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7028_ core_0.execute.pc_high_buff_out\[5\] _2771_ _2768_ core_0.execute.sreg_scratch.o_d\[5\]
+ _2957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7379__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8576__A1 _3079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8979_ _1497_ _4457_ _0655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_222_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6051__A2 _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_2645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8328__A1 core_0.execute.alu_mul_div.mul_res\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8879__A2 _4383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8033__B _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_191_2801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7000__A1 _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7551__A2 _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5562__A1 core_0.fetch.prev_request_pc\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5562__B2 net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8500__A1 _4039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7303__A2 _3223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_153_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_189_2785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5865__A2 net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8803__A2 _4328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__A1 _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5617__A2 _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7112__B _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8567__A1 _4053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_2955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_2966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_78_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_233_3307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _0841_ _0846_ _0847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7782__B _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5553__A1 core_0.fetch.prev_request_pc\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5553__B2 net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4591_ core_0.execute.rf.reg_outputs\[1\]\[9\] _0692_ _0702_ core_0.execute.rf.reg_outputs\[15\]\[9\]
+ _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_151_2328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6330_ core_0.execute.alu_mul_div.div_cur\[10\] _1833_ _2308_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_40_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4697__I net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ _2179_ _2183_ _2247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5305__B2 _1425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8000_ core_0.execute.rf.reg_outputs\[4\]\[5\] _3700_ _3689_ _3702_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5212_ _1351_ net145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6192_ _2178_ _2179_ _2180_ _2181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_110_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_244_3436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5143_ _1294_ _1295_ _1296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6805__A1 _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5074_ _1230_ _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_224_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8902_ core_0.dec_mem_long _1229_ _4413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6417__I _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_2457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5321__I core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8833_ _4335_ _4356_ _4357_ _4358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_204_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6033__A2 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8764_ _0801_ _4294_ _4305_ _4287_ _0592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5976_ core_0.execute.rf.reg_outputs\[6\]\[14\] net322 _1819_ core_0.execute.rf.reg_outputs\[12\]\[14\]
+ _1788_ core_0.execute.rf.reg_outputs\[3\]\[14\] _1966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_94_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7781__A2 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7715_ core_0.execute.rf.reg_outputs\[12\]\[13\] _3526_ _3528_ _3537_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4927_ _1105_ _1033_ _1038_ _1106_ _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5792__A1 core_0.execute.rf.reg_outputs\[1\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8695_ _4224_ _4256_ _4249_ _4257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5792__B2 core_0.execute.rf.reg_outputs\[10\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7646_ _3496_ _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4858_ _1038_ _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7533__A2 core_0.ew_data\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5544__A1 _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7577_ core_0.execute.rf.reg_outputs\[15\]\[8\] _3429_ _3422_ _3452_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4789_ _0952_ _0961_ _0969_ _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9316_ _0326_ clknet_leaf_3_i_clk core_0.execute.rf.reg_outputs\[11\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ net235 _1999_ _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__7297__A1 _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9247_ _0257_ clknet_leaf_38_i_clk core_0.execute.rf.reg_outputs\[15\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6459_ _1249_ _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_189_Right_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5847__A2 net197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_9178_ _0189_ clknet_leaf_41_i_clk core_0.execute.prev_sys vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_208_3011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8129_ _3462_ _3760_ _3775_ _0487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_237_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_237_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8797__A1 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_126_2021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_187_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_214_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6771__B core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7221__A1 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6024__A2 _1791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7772__A2 _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_219_3140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5783__A1 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__A2 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8698__B _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__A2 _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8721__A1 net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6732__B1 _2609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8210__C core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_156_Right_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_238_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A2 _1813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8788__A1 _4316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_148_2290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_221_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6015__A2 _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ core_0.execute.rf.reg_outputs\[6\]\[15\] net322 _1819_ core_0.execute.rf.reg_outputs\[12\]\[15\]
+ _1788_ core_0.execute.rf.reg_outputs\[3\]\[15\] _1820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_57_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7763__A2 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5774__A1 _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5761_ _1519_ net216 _1750_ _1751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__7068__I _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7500_ _3384_ _0249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4712_ _0893_ _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8480_ _1211_ _4069_ _4070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5692_ _1685_ _1696_ _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__8712__A1 _4224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7431_ _1366_ _2422_ _3348_ _0216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_182_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5526__A1 net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4643_ core_0.execute.rf.reg_outputs\[7\]\[5\] _0683_ _0695_ core_0.execute.rf.reg_outputs\[10\]\[5\]
+ _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6723__B1 _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7362_ _3279_ _3281_ _3282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_188_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4574_ core_0.execute.rf.reg_outputs\[5\]\[10\] net222 _0679_ core_0.execute.rf.reg_outputs\[11\]\[10\]
+ _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9101_ _0004_ clknet_leaf_130_i_clk core_0.decode.oc_alu_mode\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_24_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6313_ _2196_ _2287_ _2197_ _2293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_142_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8476__B1 _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7293_ _1254_ _2472_ _2909_ _3069_ _3214_ _3215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_40_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9032_ _0059_ clknet_leaf_87_i_clk core_0.fetch.out_buffer_data_instr\[20\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_229_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_228_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6244_ _2170_ _2171_ _2231_ _2232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_123_Right_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_229_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4888__I0 net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6175_ _2156_ _2159_ _2160_ _2163_ _2164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_209_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8779__A1 core_0.execute.sreg_scratch.o_d\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5126_ _1279_ _1280_ _1281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_34_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7451__A1 _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5057_ _1222_ _1043_ _1145_ _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer83_I _2528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7687__B _3513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_101_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8816_ core_0.execute.pc_high_out\[1\] core_0.execute.pc_high_out\[0\] core_0.execute.pc_high_out\[2\]
+ _4343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_177_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7754__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8951__A1 _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_2615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4568__A2 _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5765__A1 net313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8747_ _0890_ _4294_ _4296_ _4287_ _0584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_192_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5959_ _1772_ _1948_ _1949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_192_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8678_ _4203_ _4092_ _4242_ _1661_ _4243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_75_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7506__A2 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7629_ core_0.execute.rf.reg_outputs\[14\]\[8\] _3482_ _3486_ _3488_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output197_I net294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9244__CLK clknet_leaf_10_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_3081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9394__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_26_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output74_I net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_186_2744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7690__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6493__A2 _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7993__A2 _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_9__f_i_clk clknet_3_4_0_i_clk clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_201_2925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8942__A1 core_0.decode.i_imm_pass\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7745__A2 _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_197_2873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_225_Right_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_4 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5136__I core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6484__A2 _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7681__A1 _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7433__A1 _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7980_ core_0.execute.rf.reg_outputs\[5\]\[13\] _3679_ _3689_ _3690_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9117__CLK clknet_leaf_64_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer16 _0848_ net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_179_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer27 net254 net255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7984__A2 _3671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer38 net264 net266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6931_ _1857_ _1896_ _2731_ _2862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_77_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer49 _0813_ net277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_85_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _2792_ _2793_ _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7197__B1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8933__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7736__A2 _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8601_ _4167_ _4175_ _4176_ _0558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_159_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5813_ _0971_ _0943_ _0960_ _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_239_3379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9581_ _0591_ clknet_leaf_21_i_clk core_0.execute.sreg_scratch.o_d\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6793_ _2722_ _2725_ _1895_ _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__9267__CLK clknet_leaf_10_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6944__B1 _2768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6944__C2 _1411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8532_ net194 _2134_ _3156_ _4116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5744_ core_0.dec_jump_cond_code\[4\] _1734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_32_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8463_ _1403_ net216 _4055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4970__A2 core_0.fetch.prev_request_pc\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ _1679_ _1680_ _1676_ _1681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_127_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8161__A2 _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7414_ core_0.execute.alu_mul_div.div_res\[15\] _1742_ _3332_ _3333_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4626_ core_0.execute.rf.reg_outputs\[5\]\[6\] net222 _0679_ core_0.execute.rf.reg_outputs\[11\]\[6\]
+ _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_170_2556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8394_ _1537_ _3907_ _4005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7345_ core_0.execute.sreg_priv_control.o_d\[13\] _1693_ _2996_ net5 _2689_ _3266_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4722__A2 _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4557_ _0748_ _0749_ _0750_ _0751_ _0752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7462__S _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_229_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7276_ _3198_ _3199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6586__B _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4488_ _0685_ _0686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_9015_ _0042_ clknet_leaf_84_i_clk core_0.fetch.out_buffer_data_instr\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6227_ core_0.execute.alu_mul_div.comp _0998_ _2216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__6475__A2 _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__A1 _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6158_ core_0.execute.alu_mul_div.div_cur\[15\] _2146_ _2147_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_5_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7424__A1 _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6227__A2 _0998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5109_ _1259_ _1262_ _1264_ _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_225_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6089_ core_0.execute.rf.reg_outputs\[12\]\[3\] _1818_ _1793_ core_0.execute.rf.reg_outputs\[8\]\[3\]
+ _2079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7975__A2 _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_2685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7727__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8924__A1 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_216_3110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8152__A2 _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5910__A1 core_0.execute.rf.reg_outputs\[7\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6466__A2 _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7663__A1 _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput74 net74 dbg_pc[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_235_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput85 net85 dbg_pc[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_235_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput96 net96 dbg_r0[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_101_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6218__A2 _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7415__A1 core_0.execute.alu_mul_div.div_cur\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_1808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_2902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7966__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7718__A2 _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8915__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__A1 core_0.execute.sreg_priv_control.o_d\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5729__B2 _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8391__A2 _1829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8143__A2 _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_1937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5460_ _1009_ _1551_ _1553_ _0040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4704__A2 net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _0675_ _1486_ _1496_ _1497_ _0026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_112_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7282__S _2708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7130_ _2839_ _3055_ _3056_ _0207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7654__A1 _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6457__A2 _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7061_ _2972_ _2976_ _2985_ _2988_ _2989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_120_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4468__A1 _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6012_ _1976_ _2001_ _1930_ _2002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
.ends

