magic
tech sky130B
magscale 1 2
timestamp 1662647170
<< viali >>
rect 1869 30277 1903 30311
rect 2789 30277 2823 30311
rect 7481 30277 7515 30311
rect 13553 30277 13587 30311
rect 15117 30277 15151 30311
rect 15669 30277 15703 30311
rect 5549 30209 5583 30243
rect 6745 30209 6779 30243
rect 7205 30209 7239 30243
rect 9137 30209 9171 30243
rect 11713 30209 11747 30243
rect 14105 30209 14139 30243
rect 18153 30209 18187 30243
rect 19257 30209 19291 30243
rect 20085 30209 20119 30243
rect 21281 30209 21315 30243
rect 22017 30209 22051 30243
rect 24593 30209 24627 30243
rect 26985 30209 27019 30243
rect 27721 30209 27755 30243
rect 28457 30209 28491 30243
rect 2053 30073 2087 30107
rect 5365 30073 5399 30107
rect 9321 30073 9355 30107
rect 11897 30073 11931 30107
rect 14289 30073 14323 30107
rect 17509 30073 17543 30107
rect 18337 30073 18371 30107
rect 27169 30073 27203 30107
rect 28641 30073 28675 30107
rect 3065 30005 3099 30039
rect 15945 30005 15979 30039
rect 20269 30005 20303 30039
rect 22201 30005 22235 30039
rect 24777 30005 24811 30039
rect 26341 30005 26375 30039
rect 27905 30005 27939 30039
rect 2605 29801 2639 29835
rect 19993 29801 20027 29835
rect 22385 29801 22419 29835
rect 24501 29801 24535 29835
rect 3065 29733 3099 29767
rect 16313 29733 16347 29767
rect 12541 29665 12575 29699
rect 12817 29665 12851 29699
rect 17141 29665 17175 29699
rect 21373 29665 21407 29699
rect 22109 29665 22143 29699
rect 22845 29665 22879 29699
rect 1685 29597 1719 29631
rect 12449 29597 12483 29631
rect 16497 29597 16531 29631
rect 16589 29597 16623 29631
rect 17877 29597 17911 29631
rect 17969 29597 18003 29631
rect 18521 29597 18555 29631
rect 22017 29597 22051 29631
rect 27077 29597 27111 29631
rect 28733 29597 28767 29631
rect 16313 29529 16347 29563
rect 1501 29461 1535 29495
rect 9229 29461 9263 29495
rect 11529 29461 11563 29495
rect 17693 29461 17727 29495
rect 27629 29461 27663 29495
rect 28549 29461 28583 29495
rect 13001 29257 13035 29291
rect 1869 29189 1903 29223
rect 12909 29189 12943 29223
rect 18981 29189 19015 29223
rect 6745 29121 6779 29155
rect 7757 29121 7791 29155
rect 8769 29121 8803 29155
rect 15577 29121 15611 29155
rect 16865 29121 16899 29155
rect 16957 29121 16991 29155
rect 17141 29121 17175 29155
rect 17233 29121 17267 29155
rect 18245 29121 18279 29155
rect 19717 29121 19751 29155
rect 19901 29121 19935 29155
rect 20361 29121 20395 29155
rect 22109 29121 22143 29155
rect 22845 29121 22879 29155
rect 2513 29053 2547 29087
rect 6837 29053 6871 29087
rect 7849 29053 7883 29087
rect 8677 29053 8711 29087
rect 9689 29053 9723 29087
rect 13185 29053 13219 29087
rect 15669 29053 15703 29087
rect 2053 28985 2087 29019
rect 6377 28985 6411 29019
rect 8125 28985 8159 29019
rect 12541 28985 12575 29019
rect 21925 28985 21959 29019
rect 28273 28985 28307 29019
rect 9137 28917 9171 28951
rect 10241 28917 10275 28951
rect 15301 28917 15335 28951
rect 16681 28917 16715 28951
rect 19809 28917 19843 28951
rect 21281 28917 21315 28951
rect 22937 28917 22971 28951
rect 23305 28917 23339 28951
rect 23765 28917 23799 28951
rect 1685 28713 1719 28747
rect 6377 28713 6411 28747
rect 7205 28713 7239 28747
rect 19625 28713 19659 28747
rect 8953 28645 8987 28679
rect 16221 28645 16255 28679
rect 22109 28645 22143 28679
rect 6101 28577 6135 28611
rect 9229 28577 9263 28611
rect 11897 28577 11931 28611
rect 14841 28577 14875 28611
rect 18245 28577 18279 28611
rect 19717 28577 19751 28611
rect 20729 28577 20763 28611
rect 21925 28577 21959 28611
rect 6009 28509 6043 28543
rect 7113 28509 7147 28543
rect 7205 28509 7239 28543
rect 9321 28509 9355 28543
rect 11805 28509 11839 28543
rect 12817 28509 12851 28543
rect 13093 28509 13127 28543
rect 14565 28509 14599 28543
rect 16037 28509 16071 28543
rect 16313 28509 16347 28543
rect 19441 28509 19475 28543
rect 22109 28509 22143 28543
rect 22477 28509 22511 28543
rect 23121 28509 23155 28543
rect 23397 28509 23431 28543
rect 24409 28509 24443 28543
rect 24593 28509 24627 28543
rect 8309 28441 8343 28475
rect 10057 28441 10091 28475
rect 17417 28441 17451 28475
rect 17969 28441 18003 28475
rect 25053 28441 25087 28475
rect 6837 28373 6871 28407
rect 10517 28373 10551 28407
rect 11161 28373 11195 28407
rect 12173 28373 12207 28407
rect 12633 28373 12667 28407
rect 13001 28373 13035 28407
rect 19257 28373 19291 28407
rect 20177 28373 20211 28407
rect 21281 28373 21315 28407
rect 22937 28373 22971 28407
rect 23305 28373 23339 28407
rect 24501 28373 24535 28407
rect 7849 28169 7883 28203
rect 8953 28169 8987 28203
rect 10149 28169 10183 28203
rect 15853 28169 15887 28203
rect 19073 28169 19107 28203
rect 21925 28169 21959 28203
rect 22109 28169 22143 28203
rect 24225 28169 24259 28203
rect 24393 28169 24427 28203
rect 9413 28101 9447 28135
rect 19993 28101 20027 28135
rect 24593 28101 24627 28135
rect 7665 28033 7699 28067
rect 9137 28033 9171 28067
rect 11897 28033 11931 28067
rect 12909 28033 12943 28067
rect 13001 28033 13035 28067
rect 13185 28033 13219 28067
rect 13277 28033 13311 28067
rect 14473 28033 14507 28067
rect 15209 28033 15243 28067
rect 15372 28039 15406 28073
rect 15472 28036 15506 28070
rect 15577 28033 15611 28067
rect 18889 28033 18923 28067
rect 19165 28033 19199 28067
rect 20177 28033 20211 28067
rect 21189 28033 21223 28067
rect 22106 28033 22140 28067
rect 22569 28033 22603 28067
rect 23397 28033 23431 28067
rect 23581 28033 23615 28067
rect 25053 28033 25087 28067
rect 27997 28033 28031 28067
rect 28641 28033 28675 28067
rect 9229 27965 9263 27999
rect 11621 27965 11655 27999
rect 16681 27965 16715 27999
rect 22477 27965 22511 27999
rect 14013 27897 14047 27931
rect 28457 27897 28491 27931
rect 9413 27829 9447 27863
rect 10977 27829 11011 27863
rect 13461 27829 13495 27863
rect 18889 27829 18923 27863
rect 19809 27829 19843 27863
rect 20729 27829 20763 27863
rect 23213 27829 23247 27863
rect 24409 27829 24443 27863
rect 12633 27625 12667 27659
rect 14473 27625 14507 27659
rect 14657 27625 14691 27659
rect 19625 27625 19659 27659
rect 21005 27625 21039 27659
rect 25513 27625 25547 27659
rect 10701 27557 10735 27591
rect 16865 27557 16899 27591
rect 21741 27557 21775 27591
rect 20637 27489 20671 27523
rect 23765 27489 23799 27523
rect 10425 27421 10459 27455
rect 10517 27421 10551 27455
rect 11161 27421 11195 27455
rect 12449 27421 12483 27455
rect 12633 27421 12667 27455
rect 14657 27421 14691 27455
rect 15025 27421 15059 27455
rect 19809 27421 19843 27455
rect 19901 27421 19935 27455
rect 20085 27421 20119 27455
rect 20177 27421 20211 27455
rect 22017 27421 22051 27455
rect 23213 27421 23247 27455
rect 23673 27421 23707 27455
rect 23857 27421 23891 27455
rect 24593 27421 24627 27455
rect 25145 27421 25179 27455
rect 25605 27421 25639 27455
rect 11345 27353 11379 27387
rect 11529 27353 11563 27387
rect 13093 27353 13127 27387
rect 22937 27353 22971 27387
rect 8033 27285 8067 27319
rect 9321 27285 9355 27319
rect 9873 27285 9907 27319
rect 15761 27285 15795 27319
rect 16221 27285 16255 27319
rect 21005 27285 21039 27319
rect 21189 27285 21223 27319
rect 7389 27081 7423 27115
rect 12081 27081 12115 27115
rect 20453 27081 20487 27115
rect 23480 27081 23514 27115
rect 26249 27081 26283 27115
rect 11713 27013 11747 27047
rect 11805 27013 11839 27047
rect 12633 27013 12667 27047
rect 14749 27013 14783 27047
rect 15761 27013 15795 27047
rect 17693 27013 17727 27047
rect 19165 27013 19199 27047
rect 20085 27013 20119 27047
rect 20913 27013 20947 27047
rect 24501 27013 24535 27047
rect 25053 27013 25087 27047
rect 26341 27013 26375 27047
rect 1869 26945 1903 26979
rect 7573 26945 7607 26979
rect 7849 26945 7883 26979
rect 9781 26945 9815 26979
rect 10793 26945 10827 26979
rect 10977 26945 11011 26979
rect 11529 26945 11563 26979
rect 11897 26945 11931 26979
rect 12541 26945 12575 26979
rect 12725 26945 12759 26979
rect 14657 26945 14691 26979
rect 14933 26945 14967 26979
rect 15393 26945 15427 26979
rect 15577 26945 15611 26979
rect 16865 26945 16899 26979
rect 19349 26945 19383 26979
rect 19967 26945 20001 26979
rect 20177 26945 20211 26979
rect 20268 26945 20302 26979
rect 21097 26945 21131 26979
rect 21833 26945 21867 26979
rect 22753 26945 22787 26979
rect 23857 26945 23891 26979
rect 24869 26945 24903 26979
rect 24961 26945 24995 26979
rect 26157 26945 26191 26979
rect 7665 26877 7699 26911
rect 16957 26877 16991 26911
rect 18981 26877 19015 26911
rect 19809 26877 19843 26911
rect 21281 26877 21315 26911
rect 24317 26877 24351 26911
rect 25605 26877 25639 26911
rect 25789 26877 25823 26911
rect 10333 26809 10367 26843
rect 14933 26809 14967 26843
rect 1961 26741 1995 26775
rect 5273 26741 5307 26775
rect 7849 26741 7883 26775
rect 8309 26741 8343 26775
rect 10885 26741 10919 26775
rect 13185 26741 13219 26775
rect 14105 26741 14139 26775
rect 17141 26741 17175 26775
rect 18337 26741 18371 26775
rect 22569 26741 22603 26775
rect 23305 26741 23339 26775
rect 23489 26741 23523 26775
rect 28641 26741 28675 26775
rect 1593 26537 1627 26571
rect 5549 26537 5583 26571
rect 7113 26537 7147 26571
rect 10977 26537 11011 26571
rect 11989 26537 12023 26571
rect 14473 26537 14507 26571
rect 15209 26537 15243 26571
rect 16497 26537 16531 26571
rect 18061 26537 18095 26571
rect 19993 26537 20027 26571
rect 21005 26537 21039 26571
rect 22569 26537 22603 26571
rect 24501 26537 24535 26571
rect 6285 26469 6319 26503
rect 10517 26469 10551 26503
rect 16773 26469 16807 26503
rect 23121 26469 23155 26503
rect 4997 26401 5031 26435
rect 11253 26401 11287 26435
rect 11345 26401 11379 26435
rect 22109 26401 22143 26435
rect 4905 26333 4939 26367
rect 5089 26333 5123 26367
rect 5549 26333 5583 26367
rect 5733 26333 5767 26367
rect 7021 26333 7055 26367
rect 7205 26333 7239 26367
rect 7573 26333 7607 26367
rect 7849 26333 7883 26367
rect 9965 26333 9999 26367
rect 10103 26333 10137 26367
rect 10333 26333 10367 26367
rect 11161 26333 11195 26367
rect 11437 26333 11471 26367
rect 12173 26333 12207 26367
rect 12265 26333 12299 26367
rect 12449 26333 12483 26367
rect 12541 26333 12575 26367
rect 15393 26333 15427 26367
rect 15761 26333 15795 26367
rect 16681 26333 16715 26367
rect 16865 26333 16899 26367
rect 16957 26333 16991 26367
rect 17141 26333 17175 26367
rect 18245 26333 18279 26367
rect 18337 26333 18371 26367
rect 18586 26333 18620 26367
rect 18705 26333 18739 26367
rect 19349 26333 19383 26367
rect 19442 26333 19476 26367
rect 19625 26333 19659 26367
rect 19814 26333 19848 26367
rect 20453 26333 20487 26367
rect 20821 26333 20855 26367
rect 24409 26333 24443 26367
rect 24593 26333 24627 26367
rect 25789 26333 25823 26367
rect 25973 26333 26007 26367
rect 9505 26265 9539 26299
rect 10237 26265 10271 26299
rect 14105 26265 14139 26299
rect 14289 26265 14323 26299
rect 15485 26265 15519 26299
rect 15577 26265 15611 26299
rect 18429 26265 18463 26299
rect 19717 26265 19751 26299
rect 20637 26265 20671 26299
rect 20729 26265 20763 26299
rect 28273 26265 28307 26299
rect 28641 26265 28675 26299
rect 8309 26197 8343 26231
rect 13553 26197 13587 26231
rect 21465 26197 21499 26231
rect 25789 26197 25823 26231
rect 5181 25993 5215 26027
rect 7205 25993 7239 26027
rect 8769 25993 8803 26027
rect 11529 25993 11563 26027
rect 13369 25993 13403 26027
rect 15025 25993 15059 26027
rect 19441 25993 19475 26027
rect 19533 25993 19567 26027
rect 20729 25993 20763 26027
rect 23673 25993 23707 26027
rect 25872 25993 25906 26027
rect 5549 25925 5583 25959
rect 7665 25925 7699 25959
rect 13553 25925 13587 25959
rect 19809 25925 19843 25959
rect 22385 25925 22419 25959
rect 26249 25925 26283 25959
rect 4353 25857 4387 25891
rect 5365 25857 5399 25891
rect 5641 25857 5675 25891
rect 7021 25857 7055 25891
rect 7849 25857 7883 25891
rect 8033 25857 8067 25891
rect 8125 25857 8159 25891
rect 8677 25857 8711 25891
rect 8861 25857 8895 25891
rect 9321 25857 9355 25891
rect 10425 25857 10459 25891
rect 11713 25857 11747 25891
rect 13737 25857 13771 25891
rect 14381 25857 14415 25891
rect 15165 25857 15199 25891
rect 15301 25857 15335 25891
rect 15393 25857 15427 25891
rect 15576 25857 15610 25891
rect 15669 25857 15703 25891
rect 19257 25857 19291 25891
rect 19625 25857 19659 25891
rect 20729 25857 20763 25891
rect 20913 25857 20947 25891
rect 25605 25857 25639 25891
rect 4261 25789 4295 25823
rect 6745 25789 6779 25823
rect 11897 25789 11931 25823
rect 17233 25789 17267 25823
rect 18337 25789 18371 25823
rect 4721 25721 4755 25755
rect 7941 25721 7975 25755
rect 10977 25721 11011 25755
rect 14473 25721 14507 25755
rect 16773 25721 16807 25755
rect 21833 25721 21867 25755
rect 28641 25721 28675 25755
rect 6837 25653 6871 25687
rect 12817 25653 12851 25687
rect 17877 25653 17911 25687
rect 25881 25653 25915 25687
rect 27629 25653 27663 25687
rect 28181 25653 28215 25687
rect 4353 25449 4387 25483
rect 5273 25449 5307 25483
rect 7113 25449 7147 25483
rect 8217 25449 8251 25483
rect 13553 25449 13587 25483
rect 15761 25449 15795 25483
rect 17049 25449 17083 25483
rect 17417 25449 17451 25483
rect 19257 25449 19291 25483
rect 20821 25449 20855 25483
rect 21465 25449 21499 25483
rect 22385 25449 22419 25483
rect 23489 25449 23523 25483
rect 26893 25449 26927 25483
rect 28549 25449 28583 25483
rect 9689 25313 9723 25347
rect 17325 25313 17359 25347
rect 24685 25313 24719 25347
rect 4629 25245 4663 25279
rect 5089 25245 5123 25279
rect 5273 25245 5307 25279
rect 7389 25245 7423 25279
rect 7849 25245 7883 25279
rect 8033 25245 8067 25279
rect 8953 25245 8987 25279
rect 9137 25245 9171 25279
rect 12173 25245 12207 25279
rect 15393 25245 15427 25279
rect 15577 25245 15611 25279
rect 17417 25245 17451 25279
rect 19441 25245 19475 25279
rect 19625 25245 19659 25279
rect 19717 25245 19751 25279
rect 22569 25245 22603 25279
rect 24593 25245 24627 25279
rect 24777 25245 24811 25279
rect 25697 25245 25731 25279
rect 25881 25245 25915 25279
rect 26065 25245 26099 25279
rect 4353 25177 4387 25211
rect 7113 25177 7147 25211
rect 9045 25177 9079 25211
rect 10425 25177 10459 25211
rect 11253 25177 11287 25211
rect 17877 25177 17911 25211
rect 20177 25177 20211 25211
rect 21373 25177 21407 25211
rect 25237 25177 25271 25211
rect 26861 25177 26895 25211
rect 27077 25177 27111 25211
rect 4537 25109 4571 25143
rect 7297 25109 7331 25143
rect 10701 25109 10735 25143
rect 12725 25109 12759 25143
rect 14105 25109 14139 25143
rect 14841 25109 14875 25143
rect 16313 25109 16347 25143
rect 18429 25109 18463 25143
rect 26709 25109 26743 25143
rect 28089 25109 28123 25143
rect 8125 24905 8159 24939
rect 14841 24905 14875 24939
rect 22477 24905 22511 24939
rect 25881 24905 25915 24939
rect 22661 24837 22695 24871
rect 1409 24769 1443 24803
rect 4537 24769 4571 24803
rect 4721 24769 4755 24803
rect 8033 24769 8067 24803
rect 8217 24769 8251 24803
rect 13093 24769 13127 24803
rect 13461 24769 13495 24803
rect 13921 24769 13955 24803
rect 21833 24769 21867 24803
rect 22845 24769 22879 24803
rect 23397 24769 23431 24803
rect 25237 24769 25271 24803
rect 25421 24769 25455 24803
rect 25516 24775 25550 24809
rect 25651 24769 25685 24803
rect 12541 24701 12575 24735
rect 14013 24701 14047 24735
rect 10333 24633 10367 24667
rect 26341 24633 26375 24667
rect 27537 24633 27571 24667
rect 1593 24565 1627 24599
rect 4905 24565 4939 24599
rect 7481 24565 7515 24599
rect 9229 24565 9263 24599
rect 18797 24565 18831 24599
rect 19533 24565 19567 24599
rect 19993 24565 20027 24599
rect 24317 24565 24351 24599
rect 26985 24565 27019 24599
rect 28457 24565 28491 24599
rect 1409 24361 1443 24395
rect 10425 24361 10459 24395
rect 11621 24361 11655 24395
rect 12541 24361 12575 24395
rect 23765 24361 23799 24395
rect 5641 24293 5675 24327
rect 18613 24293 18647 24327
rect 22569 24293 22603 24327
rect 24869 24293 24903 24327
rect 18429 24225 18463 24259
rect 21741 24225 21775 24259
rect 25237 24225 25271 24259
rect 4261 24157 4295 24191
rect 4445 24157 4479 24191
rect 4905 24157 4939 24191
rect 5089 24157 5123 24191
rect 5549 24157 5583 24191
rect 5733 24157 5767 24191
rect 7665 24157 7699 24191
rect 9229 24157 9263 24191
rect 9321 24157 9355 24191
rect 10149 24157 10183 24191
rect 11805 24157 11839 24191
rect 14565 24157 14599 24191
rect 18705 24157 18739 24191
rect 19717 24157 19751 24191
rect 20085 24157 20119 24191
rect 21925 24157 21959 24191
rect 22748 24157 22782 24191
rect 22845 24157 22879 24191
rect 23120 24157 23154 24191
rect 23213 24157 23247 24191
rect 25513 24157 25547 24191
rect 25973 24157 26007 24191
rect 26709 24157 26743 24191
rect 4997 24089 5031 24123
rect 7021 24089 7055 24123
rect 8125 24089 8159 24123
rect 11069 24089 11103 24123
rect 11989 24089 12023 24123
rect 21097 24089 21131 24123
rect 22937 24089 22971 24123
rect 25028 24089 25062 24123
rect 25145 24089 25179 24123
rect 4353 24021 4387 24055
rect 9413 24021 9447 24055
rect 10609 24021 10643 24055
rect 14657 24021 14691 24055
rect 18429 24021 18463 24055
rect 20545 24021 20579 24055
rect 22109 24021 22143 24055
rect 26157 24021 26191 24055
rect 27353 24021 27387 24055
rect 28089 24021 28123 24055
rect 28733 24021 28767 24055
rect 4629 23817 4663 23851
rect 6745 23817 6779 23851
rect 9045 23817 9079 23851
rect 10241 23817 10275 23851
rect 12173 23817 12207 23851
rect 14657 23817 14691 23851
rect 18981 23817 19015 23851
rect 19901 23817 19935 23851
rect 21833 23817 21867 23851
rect 22937 23817 22971 23851
rect 6377 23749 6411 23783
rect 7849 23749 7883 23783
rect 14841 23749 14875 23783
rect 22477 23749 22511 23783
rect 4721 23681 4755 23715
rect 5181 23681 5215 23715
rect 5365 23681 5399 23715
rect 6561 23681 6595 23715
rect 6837 23681 6871 23715
rect 7665 23681 7699 23715
rect 8953 23681 8987 23715
rect 9137 23681 9171 23715
rect 9597 23681 9631 23715
rect 9690 23681 9724 23715
rect 9873 23681 9907 23715
rect 9965 23681 9999 23715
rect 10103 23681 10137 23715
rect 13001 23681 13035 23715
rect 13461 23681 13495 23715
rect 13645 23681 13679 23715
rect 13829 23681 13863 23715
rect 16957 23681 16991 23715
rect 17049 23681 17083 23715
rect 17141 23681 17175 23715
rect 17325 23681 17359 23715
rect 19165 23681 19199 23715
rect 19349 23681 19383 23715
rect 21005 23681 21039 23715
rect 24777 23681 24811 23715
rect 24961 23681 24995 23715
rect 25237 23681 25271 23715
rect 25973 23681 26007 23715
rect 28457 23681 28491 23715
rect 4261 23613 4295 23647
rect 7481 23613 7515 23647
rect 11621 23613 11655 23647
rect 20361 23613 20395 23647
rect 23949 23613 23983 23647
rect 5273 23545 5307 23579
rect 8401 23545 8435 23579
rect 12817 23545 12851 23579
rect 15209 23545 15243 23579
rect 15761 23545 15795 23579
rect 22753 23545 22787 23579
rect 24593 23545 24627 23579
rect 25789 23545 25823 23579
rect 27813 23545 27847 23579
rect 4445 23477 4479 23511
rect 10793 23477 10827 23511
rect 14841 23477 14875 23511
rect 16681 23477 16715 23511
rect 23397 23477 23431 23511
rect 25145 23477 25179 23511
rect 27077 23477 27111 23511
rect 28641 23477 28675 23511
rect 4353 23273 4387 23307
rect 6193 23273 6227 23307
rect 11345 23273 11379 23307
rect 14197 23273 14231 23307
rect 15853 23273 15887 23307
rect 17049 23273 17083 23307
rect 20729 23273 20763 23307
rect 22753 23273 22787 23307
rect 13185 23205 13219 23239
rect 10057 23137 10091 23171
rect 11069 23137 11103 23171
rect 12173 23137 12207 23171
rect 12633 23137 12667 23171
rect 16405 23137 16439 23171
rect 19257 23137 19291 23171
rect 24685 23137 24719 23171
rect 25513 23137 25547 23171
rect 26893 23137 26927 23171
rect 27537 23137 27571 23171
rect 27813 23137 27847 23171
rect 28089 23137 28123 23171
rect 28733 23137 28767 23171
rect 4261 23069 4295 23103
rect 4353 23069 4387 23103
rect 4721 23069 4755 23103
rect 6193 23069 6227 23103
rect 7619 23069 7653 23103
rect 7977 23069 8011 23103
rect 8125 23069 8159 23103
rect 9965 23069 9999 23103
rect 10185 23069 10219 23103
rect 10701 23069 10735 23103
rect 10885 23069 10919 23103
rect 10977 23069 11011 23103
rect 11161 23069 11195 23103
rect 12357 23069 12391 23103
rect 12541 23069 12575 23103
rect 13369 23069 13403 23103
rect 14381 23069 14415 23103
rect 15209 23069 15243 23103
rect 15357 23069 15391 23103
rect 15715 23069 15749 23103
rect 16497 23069 16531 23103
rect 16868 23069 16902 23103
rect 18429 23069 18463 23103
rect 18705 23069 18739 23103
rect 19487 23069 19521 23103
rect 19622 23069 19656 23103
rect 19722 23069 19756 23103
rect 19901 23069 19935 23103
rect 20913 23069 20947 23103
rect 21189 23069 21223 23103
rect 21925 23069 21959 23103
rect 24501 23069 24535 23103
rect 24777 23069 24811 23103
rect 25145 23069 25179 23103
rect 27696 23069 27730 23103
rect 28549 23069 28583 23103
rect 5733 23001 5767 23035
rect 6285 23001 6319 23035
rect 6469 23001 6503 23035
rect 7757 23001 7791 23035
rect 7849 23001 7883 23035
rect 9781 23001 9815 23035
rect 10057 23001 10091 23035
rect 15485 23001 15519 23035
rect 15577 23001 15611 23035
rect 23305 23001 23339 23035
rect 1501 22933 1535 22967
rect 4077 22933 4111 22967
rect 7021 22933 7055 22967
rect 7481 22933 7515 22967
rect 9321 22933 9355 22967
rect 16865 22933 16899 22967
rect 18245 22933 18279 22967
rect 18613 22933 18647 22967
rect 21097 22933 21131 22967
rect 22201 22933 22235 22967
rect 25973 22933 26007 22967
rect 4169 22729 4203 22763
rect 6837 22729 6871 22763
rect 9689 22729 9723 22763
rect 10241 22729 10275 22763
rect 12081 22729 12115 22763
rect 13001 22729 13035 22763
rect 15025 22729 15059 22763
rect 16681 22729 16715 22763
rect 18705 22729 18739 22763
rect 19349 22729 19383 22763
rect 21189 22729 21223 22763
rect 25329 22729 25363 22763
rect 26065 22729 26099 22763
rect 3341 22661 3375 22695
rect 7481 22661 7515 22695
rect 8861 22661 8895 22695
rect 11989 22661 12023 22695
rect 13645 22661 13679 22695
rect 14197 22661 14231 22695
rect 25446 22661 25480 22695
rect 26985 22661 27019 22695
rect 1593 22593 1627 22627
rect 2513 22593 2547 22627
rect 2973 22593 3007 22627
rect 3985 22593 4019 22627
rect 4261 22593 4295 22627
rect 6929 22593 6963 22627
rect 7389 22593 7423 22627
rect 7573 22593 7607 22627
rect 13001 22593 13035 22627
rect 15025 22593 15059 22627
rect 15209 22593 15243 22627
rect 16865 22593 16899 22627
rect 16957 22593 16991 22627
rect 17877 22593 17911 22627
rect 21833 22593 21867 22627
rect 22569 22593 22603 22627
rect 22661 22593 22695 22627
rect 22845 22593 22879 22627
rect 22937 22593 22971 22627
rect 23581 22593 23615 22627
rect 24961 22593 24995 22627
rect 27997 22593 28031 22627
rect 22109 22525 22143 22559
rect 25237 22525 25271 22559
rect 1777 22457 1811 22491
rect 20729 22457 20763 22491
rect 24133 22457 24167 22491
rect 3801 22389 3835 22423
rect 8217 22389 8251 22423
rect 10701 22389 10735 22423
rect 20085 22389 20119 22423
rect 23121 22389 23155 22423
rect 25605 22389 25639 22423
rect 28089 22389 28123 22423
rect 2237 22185 2271 22219
rect 11253 22185 11287 22219
rect 12449 22185 12483 22219
rect 19257 22185 19291 22219
rect 7389 22117 7423 22151
rect 2053 22049 2087 22083
rect 6837 22049 6871 22083
rect 9505 22049 9539 22083
rect 9689 22049 9723 22083
rect 14933 22049 14967 22083
rect 19901 22049 19935 22083
rect 21348 22049 21382 22083
rect 21465 22049 21499 22083
rect 21741 22049 21775 22083
rect 23029 22049 23063 22083
rect 24501 22049 24535 22083
rect 26157 22049 26191 22083
rect 28089 22049 28123 22083
rect 1961 21981 1995 22015
rect 2789 21981 2823 22015
rect 3985 21981 4019 22015
rect 7297 21981 7331 22015
rect 7481 21981 7515 22015
rect 14381 21981 14415 22015
rect 14473 21981 14507 22015
rect 14657 21981 14691 22015
rect 14749 21981 14783 22015
rect 18137 21981 18171 22015
rect 18337 21981 18371 22015
rect 18521 21981 18555 22015
rect 18613 21981 18647 22015
rect 19625 21981 19659 22015
rect 21189 21981 21223 22015
rect 22201 21981 22235 22015
rect 22385 21981 22419 22015
rect 23213 21981 23247 22015
rect 25513 21981 25547 22015
rect 7941 21913 7975 21947
rect 10609 21913 10643 21947
rect 18245 21913 18279 21947
rect 19717 21913 19751 21947
rect 25329 21913 25363 21947
rect 27905 21913 27939 21947
rect 3893 21845 3927 21879
rect 9781 21845 9815 21879
rect 10149 21845 10183 21879
rect 13185 21845 13219 21879
rect 17509 21845 17543 21879
rect 17969 21845 18003 21879
rect 20545 21845 20579 21879
rect 23121 21845 23155 21879
rect 23581 21845 23615 21879
rect 26617 21845 26651 21879
rect 27537 21845 27571 21879
rect 27997 21845 28031 21879
rect 4629 21641 4663 21675
rect 8677 21641 8711 21675
rect 9229 21641 9263 21675
rect 10885 21641 10919 21675
rect 14105 21641 14139 21675
rect 15761 21641 15795 21675
rect 18245 21641 18279 21675
rect 21833 21641 21867 21675
rect 27353 21641 27387 21675
rect 28549 21641 28583 21675
rect 12725 21573 12759 21607
rect 14473 21573 14507 21607
rect 15117 21573 15151 21607
rect 15209 21573 15243 21607
rect 18337 21573 18371 21607
rect 26157 21573 26191 21607
rect 3433 21505 3467 21539
rect 4261 21505 4295 21539
rect 4445 21505 4479 21539
rect 9408 21505 9442 21539
rect 9496 21505 9530 21539
rect 9597 21505 9631 21539
rect 9725 21505 9759 21539
rect 9873 21505 9907 21539
rect 12633 21505 12667 21539
rect 12817 21505 12851 21539
rect 13277 21505 13311 21539
rect 13461 21505 13495 21539
rect 14289 21505 14323 21539
rect 14381 21505 14415 21539
rect 14657 21505 14691 21539
rect 15485 21505 15519 21539
rect 17049 21505 17083 21539
rect 20821 21505 20855 21539
rect 21005 21505 21039 21539
rect 22477 21505 22511 21539
rect 23029 21505 23063 21539
rect 23397 21505 23431 21539
rect 24041 21505 24075 21539
rect 24133 21505 24167 21539
rect 25237 21505 25271 21539
rect 28733 21505 28767 21539
rect 3525 21437 3559 21471
rect 15577 21437 15611 21471
rect 17141 21437 17175 21471
rect 17325 21437 17359 21471
rect 18521 21437 18555 21471
rect 20269 21437 20303 21471
rect 24317 21437 24351 21471
rect 27445 21437 27479 21471
rect 27537 21437 27571 21471
rect 10333 21369 10367 21403
rect 16681 21369 16715 21403
rect 19073 21369 19107 21403
rect 19717 21369 19751 21403
rect 23305 21369 23339 21403
rect 25513 21369 25547 21403
rect 2513 21301 2547 21335
rect 3709 21301 3743 21335
rect 11529 21301 11563 21335
rect 13461 21301 13495 21335
rect 17877 21301 17911 21335
rect 20913 21301 20947 21335
rect 24225 21301 24259 21335
rect 26985 21301 27019 21335
rect 9321 21097 9355 21131
rect 11621 21097 11655 21131
rect 12449 21097 12483 21131
rect 13553 21097 13587 21131
rect 16589 21097 16623 21131
rect 17233 21097 17267 21131
rect 17877 21097 17911 21131
rect 26249 21097 26283 21131
rect 8401 21029 8435 21063
rect 26801 21029 26835 21063
rect 22569 20961 22603 20995
rect 26065 20961 26099 20995
rect 27445 20961 27479 20995
rect 27721 20961 27755 20995
rect 27997 20961 28031 20995
rect 9505 20893 9539 20927
rect 9670 20893 9704 20927
rect 9781 20893 9815 20927
rect 9873 20871 9907 20905
rect 11529 20893 11563 20927
rect 12449 20893 12483 20927
rect 12633 20893 12667 20927
rect 14284 20893 14318 20927
rect 14656 20893 14690 20927
rect 14749 20893 14783 20927
rect 16405 20893 16439 20927
rect 16589 20893 16623 20927
rect 17141 20893 17175 20927
rect 17325 20893 17359 20927
rect 20729 20893 20763 20927
rect 20913 20893 20947 20927
rect 21649 20893 21683 20927
rect 23397 20893 23431 20927
rect 23581 20893 23615 20927
rect 26341 20893 26375 20927
rect 27604 20893 27638 20927
rect 28457 20893 28491 20927
rect 28641 20893 28675 20927
rect 10885 20825 10919 20859
rect 14381 20825 14415 20859
rect 14473 20825 14507 20859
rect 20821 20825 20855 20859
rect 21925 20825 21959 20859
rect 6561 20757 6595 20791
rect 7849 20757 7883 20791
rect 10609 20757 10643 20791
rect 14105 20757 14139 20791
rect 18705 20757 18739 20791
rect 19257 20757 19291 20791
rect 23489 20757 23523 20791
rect 24685 20757 24719 20791
rect 25513 20757 25547 20791
rect 26065 20757 26099 20791
rect 1961 20553 1995 20587
rect 11989 20553 12023 20587
rect 12633 20553 12667 20587
rect 16773 20553 16807 20587
rect 17969 20553 18003 20587
rect 25053 20553 25087 20587
rect 4629 20485 4663 20519
rect 9689 20485 9723 20519
rect 14105 20485 14139 20519
rect 25421 20485 25455 20519
rect 26985 20485 27019 20519
rect 3157 20417 3191 20451
rect 3341 20417 3375 20451
rect 3617 20417 3651 20451
rect 4537 20417 4571 20451
rect 4721 20417 4755 20451
rect 7113 20417 7147 20451
rect 8769 20417 8803 20451
rect 8953 20417 8987 20451
rect 9505 20417 9539 20451
rect 9781 20417 9815 20451
rect 9873 20417 9907 20451
rect 12817 20417 12851 20451
rect 13093 20417 13127 20451
rect 13921 20417 13955 20451
rect 14197 20417 14231 20451
rect 14289 20417 14323 20451
rect 19257 20417 19291 20451
rect 19533 20417 19567 20451
rect 21833 20417 21867 20451
rect 24225 20417 24259 20451
rect 24501 20417 24535 20451
rect 25513 20417 25547 20451
rect 3525 20349 3559 20383
rect 7205 20349 7239 20383
rect 7573 20349 7607 20383
rect 8585 20349 8619 20383
rect 19441 20349 19475 20383
rect 23765 20349 23799 20383
rect 24593 20349 24627 20383
rect 25697 20349 25731 20383
rect 2513 20281 2547 20315
rect 3433 20281 3467 20315
rect 19073 20281 19107 20315
rect 23121 20281 23155 20315
rect 3801 20213 3835 20247
rect 5825 20213 5859 20247
rect 6469 20213 6503 20247
rect 6929 20213 6963 20247
rect 8033 20213 8067 20247
rect 10057 20213 10091 20247
rect 10609 20213 10643 20247
rect 13001 20213 13035 20247
rect 14473 20213 14507 20247
rect 17509 20213 17543 20247
rect 19349 20213 19383 20247
rect 19993 20213 20027 20247
rect 20729 20213 20763 20247
rect 26249 20213 26283 20247
rect 27813 20213 27847 20247
rect 28273 20213 28307 20247
rect 3065 20009 3099 20043
rect 3249 20009 3283 20043
rect 5917 20009 5951 20043
rect 6101 20009 6135 20043
rect 8309 20009 8343 20043
rect 9137 20009 9171 20043
rect 9965 20009 9999 20043
rect 21925 20009 21959 20043
rect 26157 20009 26191 20043
rect 3893 19941 3927 19975
rect 5273 19941 5307 19975
rect 10609 19941 10643 19975
rect 18429 19941 18463 19975
rect 27261 19941 27295 19975
rect 6193 19873 6227 19907
rect 13277 19873 13311 19907
rect 13461 19873 13495 19907
rect 17233 19873 17267 19907
rect 18521 19873 18555 19907
rect 19257 19873 19291 19907
rect 21097 19873 21131 19907
rect 1685 19805 1719 19839
rect 2145 19805 2179 19839
rect 2329 19805 2363 19839
rect 2789 19805 2823 19839
rect 4077 19805 4111 19839
rect 4261 19805 4295 19839
rect 4445 19805 4479 19839
rect 4537 19805 4571 19839
rect 4997 19805 5031 19839
rect 5273 19805 5307 19839
rect 5457 19805 5491 19839
rect 6469 19805 6503 19839
rect 7113 19805 7147 19839
rect 7205 19805 7239 19839
rect 7297 19805 7331 19839
rect 9781 19805 9815 19839
rect 10057 19805 10091 19839
rect 14289 19805 14323 19839
rect 14381 19805 14415 19839
rect 14565 19805 14599 19839
rect 14657 19805 14691 19839
rect 16129 19805 16163 19839
rect 16957 19805 16991 19839
rect 18305 19805 18339 19839
rect 18613 19805 18647 19839
rect 20269 19805 20303 19839
rect 21005 19805 21039 19839
rect 21281 19805 21315 19839
rect 21373 19805 21407 19839
rect 22661 19805 22695 19839
rect 22753 19805 22787 19839
rect 23857 19805 23891 19839
rect 24869 19805 24903 19839
rect 25513 19805 25547 19839
rect 27997 19805 28031 19839
rect 4169 19737 4203 19771
rect 9689 19737 9723 19771
rect 10149 19737 10183 19771
rect 10793 19737 10827 19771
rect 10977 19737 11011 19771
rect 11529 19737 11563 19771
rect 17049 19737 17083 19771
rect 1501 19669 1535 19703
rect 2329 19669 2363 19703
rect 6929 19669 6963 19703
rect 11989 19669 12023 19703
rect 12817 19669 12851 19703
rect 13185 19669 13219 19703
rect 14105 19669 14139 19703
rect 15577 19669 15611 19703
rect 16589 19669 16623 19703
rect 18153 19669 18187 19703
rect 20913 19669 20947 19703
rect 22477 19669 22511 19703
rect 28181 19669 28215 19703
rect 2789 19465 2823 19499
rect 4070 19465 4104 19499
rect 4721 19465 4755 19499
rect 5273 19465 5307 19499
rect 6821 19465 6855 19499
rect 10057 19465 10091 19499
rect 10241 19465 10275 19499
rect 16865 19465 16899 19499
rect 17325 19465 17359 19499
rect 19901 19465 19935 19499
rect 20361 19465 20395 19499
rect 27813 19465 27847 19499
rect 2421 19397 2455 19431
rect 3985 19397 4019 19431
rect 7021 19397 7055 19431
rect 9137 19397 9171 19431
rect 10701 19397 10735 19431
rect 20269 19397 20303 19431
rect 23489 19397 23523 19431
rect 1869 19329 1903 19363
rect 2329 19329 2363 19363
rect 2605 19329 2639 19363
rect 3893 19329 3927 19363
rect 4169 19329 4203 19363
rect 8953 19329 8987 19363
rect 9597 19329 9631 19363
rect 9689 19329 9723 19363
rect 10060 19329 10094 19363
rect 13829 19329 13863 19363
rect 14013 19329 14047 19363
rect 16681 19329 16715 19363
rect 16865 19329 16899 19363
rect 23305 19329 23339 19363
rect 24593 19329 24627 19363
rect 5825 19261 5859 19295
rect 8769 19261 8803 19295
rect 17969 19261 18003 19295
rect 20453 19261 20487 19295
rect 23949 19261 23983 19295
rect 24777 19261 24811 19295
rect 26341 19261 26375 19295
rect 27905 19261 27939 19295
rect 28089 19261 28123 19295
rect 1777 19125 1811 19159
rect 3249 19125 3283 19159
rect 6653 19125 6687 19159
rect 6837 19125 6871 19159
rect 7573 19125 7607 19159
rect 8217 19125 8251 19159
rect 13921 19125 13955 19159
rect 16129 19125 16163 19159
rect 19349 19125 19383 19159
rect 21281 19125 21315 19159
rect 23121 19125 23155 19159
rect 27445 19125 27479 19159
rect 28641 19125 28675 19159
rect 2237 18921 2271 18955
rect 4721 18921 4755 18955
rect 7205 18921 7239 18955
rect 7849 18921 7883 18955
rect 9505 18921 9539 18955
rect 10241 18921 10275 18955
rect 15485 18921 15519 18955
rect 17877 18921 17911 18955
rect 21649 18921 21683 18955
rect 23857 18921 23891 18955
rect 28549 18921 28583 18955
rect 5181 18853 5215 18887
rect 16129 18785 16163 18819
rect 17141 18785 17175 18819
rect 17325 18785 17359 18819
rect 18429 18785 18463 18819
rect 21005 18785 21039 18819
rect 26709 18785 26743 18819
rect 27905 18785 27939 18819
rect 2237 18717 2271 18751
rect 2329 18717 2363 18751
rect 5917 18717 5951 18751
rect 6009 18717 6043 18751
rect 6193 18717 6227 18751
rect 6285 18717 6319 18751
rect 7113 18717 7147 18751
rect 7297 18717 7331 18751
rect 8309 18717 8343 18751
rect 9321 18717 9355 18751
rect 9505 18717 9539 18751
rect 14105 18717 14139 18751
rect 14289 18717 14323 18751
rect 15945 18717 15979 18751
rect 19717 18717 19751 18751
rect 20637 18717 20671 18751
rect 21097 18717 21131 18751
rect 21833 18717 21867 18751
rect 24409 18717 24443 18751
rect 24593 18717 24627 18751
rect 26525 18717 26559 18751
rect 27721 18717 27755 18751
rect 28733 18717 28767 18751
rect 2513 18649 2547 18683
rect 19901 18649 19935 18683
rect 20729 18649 20763 18683
rect 1685 18581 1719 18615
rect 5733 18581 5767 18615
rect 14105 18581 14139 18615
rect 15853 18581 15887 18615
rect 16681 18581 16715 18615
rect 17049 18581 17083 18615
rect 18245 18581 18279 18615
rect 18337 18581 18371 18615
rect 19533 18581 19567 18615
rect 20361 18581 20395 18615
rect 20821 18581 20855 18615
rect 24501 18581 24535 18615
rect 26157 18581 26191 18615
rect 26617 18581 26651 18615
rect 27353 18581 27387 18615
rect 27813 18581 27847 18615
rect 9137 18377 9171 18411
rect 9965 18377 9999 18411
rect 14473 18377 14507 18411
rect 16681 18377 16715 18411
rect 17785 18377 17819 18411
rect 20545 18377 20579 18411
rect 28181 18377 28215 18411
rect 2237 18309 2271 18343
rect 4997 18309 5031 18343
rect 14749 18309 14783 18343
rect 14841 18309 14875 18343
rect 18245 18309 18279 18343
rect 23489 18309 23523 18343
rect 23673 18309 23707 18343
rect 1869 18241 1903 18275
rect 4077 18241 4111 18275
rect 6745 18241 6779 18275
rect 6929 18241 6963 18275
rect 7665 18241 7699 18275
rect 7849 18241 7883 18275
rect 8309 18241 8343 18275
rect 11805 18241 11839 18275
rect 12081 18241 12115 18275
rect 14657 18241 14691 18275
rect 15025 18241 15059 18275
rect 16865 18241 16899 18275
rect 17049 18241 17083 18275
rect 17141 18241 17175 18275
rect 20729 18241 20763 18275
rect 21189 18241 21223 18275
rect 27169 18241 27203 18275
rect 27261 18241 27295 18275
rect 3985 18173 4019 18207
rect 6837 18173 6871 18207
rect 11897 18173 11931 18207
rect 16957 18173 16991 18207
rect 20821 18173 20855 18207
rect 23765 18173 23799 18207
rect 26985 18173 27019 18207
rect 11989 18105 12023 18139
rect 23213 18105 23247 18139
rect 4445 18037 4479 18071
rect 5273 18037 5307 18071
rect 7757 18037 7791 18071
rect 10425 18037 10459 18071
rect 11621 18037 11655 18071
rect 14013 18037 14047 18071
rect 16129 18037 16163 18071
rect 19993 18037 20027 18071
rect 21097 18037 21131 18071
rect 27077 18037 27111 18071
rect 10977 17833 11011 17867
rect 17877 17833 17911 17867
rect 18613 17833 18647 17867
rect 26985 17833 27019 17867
rect 28733 17833 28767 17867
rect 1593 17765 1627 17799
rect 4169 17765 4203 17799
rect 13185 17765 13219 17799
rect 16681 17765 16715 17799
rect 20545 17765 20579 17799
rect 22385 17765 22419 17799
rect 6469 17697 6503 17731
rect 7113 17697 7147 17731
rect 7297 17697 7331 17731
rect 7389 17697 7423 17731
rect 11069 17697 11103 17731
rect 17141 17697 17175 17731
rect 17325 17697 17359 17731
rect 25421 17697 25455 17731
rect 27629 17697 27663 17731
rect 4353 17629 4387 17663
rect 4629 17629 4663 17663
rect 5733 17629 5767 17663
rect 6377 17629 6411 17663
rect 6561 17629 6595 17663
rect 7205 17629 7239 17663
rect 8217 17629 8251 17663
rect 9500 17629 9534 17663
rect 9817 17629 9851 17663
rect 9965 17629 9999 17663
rect 10793 17629 10827 17663
rect 10885 17629 10919 17663
rect 13093 17629 13127 17663
rect 13277 17629 13311 17663
rect 13369 17629 13403 17663
rect 14289 17629 14323 17663
rect 16037 17629 16071 17663
rect 16221 17629 16255 17663
rect 19349 17629 19383 17663
rect 19717 17629 19751 17663
rect 21649 17629 21683 17663
rect 21833 17629 21867 17663
rect 24777 17629 24811 17663
rect 24961 17629 24995 17663
rect 27721 17629 27755 17663
rect 4261 17561 4295 17595
rect 4997 17561 5031 17595
rect 8401 17561 8435 17595
rect 9597 17561 9631 17595
rect 9689 17561 9723 17595
rect 14473 17561 14507 17595
rect 15577 17561 15611 17595
rect 17049 17561 17083 17595
rect 5825 17493 5859 17527
rect 7573 17493 7607 17527
rect 8033 17493 8067 17527
rect 9321 17493 9355 17527
rect 11621 17493 11655 17527
rect 12909 17493 12943 17527
rect 14105 17493 14139 17527
rect 16129 17493 16163 17527
rect 21741 17493 21775 17527
rect 24777 17493 24811 17527
rect 26341 17493 26375 17527
rect 27813 17493 27847 17527
rect 28181 17493 28215 17527
rect 4813 17289 4847 17323
rect 7573 17289 7607 17323
rect 13185 17289 13219 17323
rect 16773 17289 16807 17323
rect 21281 17289 21315 17323
rect 23397 17289 23431 17323
rect 28273 17289 28307 17323
rect 9873 17221 9907 17255
rect 20361 17221 20395 17255
rect 24133 17221 24167 17255
rect 2145 17153 2179 17187
rect 7573 17153 7607 17187
rect 7757 17153 7791 17187
rect 9505 17153 9539 17187
rect 9597 17153 9631 17187
rect 9781 17153 9815 17187
rect 9965 17153 9999 17187
rect 11897 17153 11931 17187
rect 11989 17153 12023 17187
rect 12081 17153 12115 17187
rect 12265 17153 12299 17187
rect 13369 17153 13403 17187
rect 13645 17153 13679 17187
rect 19349 17153 19383 17187
rect 19533 17153 19567 17187
rect 21833 17153 21867 17187
rect 22109 17153 22143 17187
rect 22845 17153 22879 17187
rect 23121 17153 23155 17187
rect 23213 17153 23247 17187
rect 27261 17153 27295 17187
rect 27353 17153 27387 17187
rect 2237 17085 2271 17119
rect 10057 17085 10091 17119
rect 13461 17085 13495 17119
rect 21925 17085 21959 17119
rect 27077 17085 27111 17119
rect 6469 17017 6503 17051
rect 8493 17017 8527 17051
rect 24317 17017 24351 17051
rect 1869 16949 1903 16983
rect 5825 16949 5859 16983
rect 7113 16949 7147 16983
rect 9045 16949 9079 16983
rect 10609 16949 10643 16983
rect 11621 16949 11655 16983
rect 13645 16949 13679 16983
rect 21833 16949 21867 16983
rect 22293 16949 22327 16983
rect 22937 16949 22971 16983
rect 27169 16949 27203 16983
rect 1777 16745 1811 16779
rect 2881 16745 2915 16779
rect 5181 16745 5215 16779
rect 7205 16745 7239 16779
rect 7941 16745 7975 16779
rect 9505 16745 9539 16779
rect 9689 16745 9723 16779
rect 10333 16745 10367 16779
rect 12633 16745 12667 16779
rect 19809 16745 19843 16779
rect 21281 16745 21315 16779
rect 27813 16745 27847 16779
rect 11529 16677 11563 16711
rect 18153 16677 18187 16711
rect 2237 16609 2271 16643
rect 9045 16609 9079 16643
rect 13093 16609 13127 16643
rect 14841 16609 14875 16643
rect 23121 16609 23155 16643
rect 23305 16609 23339 16643
rect 25237 16609 25271 16643
rect 25421 16609 25455 16643
rect 27077 16609 27111 16643
rect 27629 16609 27663 16643
rect 2145 16541 2179 16575
rect 11713 16541 11747 16575
rect 11897 16541 11931 16575
rect 11989 16541 12023 16575
rect 12817 16541 12851 16575
rect 13001 16541 13035 16575
rect 19717 16541 19751 16575
rect 19993 16541 20027 16575
rect 20821 16541 20855 16575
rect 21005 16541 21039 16575
rect 21097 16541 21131 16575
rect 21373 16541 21407 16575
rect 21833 16541 21867 16575
rect 23029 16541 23063 16575
rect 25145 16541 25179 16575
rect 27905 16541 27939 16575
rect 28733 16541 28767 16575
rect 9873 16473 9907 16507
rect 14657 16473 14691 16507
rect 26801 16473 26835 16507
rect 26893 16473 26927 16507
rect 27629 16473 27663 16507
rect 9673 16405 9707 16439
rect 14289 16405 14323 16439
rect 14749 16405 14783 16439
rect 17509 16405 17543 16439
rect 22661 16405 22695 16439
rect 24777 16405 24811 16439
rect 26433 16405 26467 16439
rect 28549 16405 28583 16439
rect 9229 16201 9263 16235
rect 10057 16201 10091 16235
rect 15117 16201 15151 16235
rect 17141 16201 17175 16235
rect 20177 16201 20211 16235
rect 22845 16201 22879 16235
rect 23489 16201 23523 16235
rect 24133 16201 24167 16235
rect 24501 16201 24535 16235
rect 27353 16201 27387 16235
rect 3801 16133 3835 16167
rect 3985 16133 4019 16167
rect 15025 16133 15059 16167
rect 17049 16133 17083 16167
rect 28181 16133 28215 16167
rect 1409 16065 1443 16099
rect 2053 16065 2087 16099
rect 4077 16065 4111 16099
rect 6745 16065 6779 16099
rect 6837 16065 6871 16099
rect 7021 16065 7055 16099
rect 7113 16065 7147 16099
rect 7573 16065 7607 16099
rect 11897 16065 11931 16099
rect 12081 16065 12115 16099
rect 12817 16065 12851 16099
rect 13737 16065 13771 16099
rect 13921 16065 13955 16099
rect 18429 16065 18463 16099
rect 18613 16065 18647 16099
rect 18705 16065 18739 16099
rect 18889 16065 18923 16099
rect 19349 16065 19383 16099
rect 20545 16065 20579 16099
rect 22753 16065 22787 16099
rect 22937 16065 22971 16099
rect 27445 16065 27479 16099
rect 28365 16065 28399 16099
rect 28457 16065 28491 16099
rect 13093 15997 13127 16031
rect 15209 15997 15243 16031
rect 17325 15997 17359 16031
rect 18245 15997 18279 16031
rect 18521 15997 18555 16031
rect 20637 15997 20671 16031
rect 20729 15997 20763 16031
rect 24593 15997 24627 16031
rect 24685 15997 24719 16031
rect 27537 15997 27571 16031
rect 28181 15997 28215 16031
rect 1593 15929 1627 15963
rect 7665 15929 7699 15963
rect 8309 15929 8343 15963
rect 13553 15929 13587 15963
rect 16681 15929 16715 15963
rect 4077 15861 4111 15895
rect 6561 15861 6595 15895
rect 11897 15861 11931 15895
rect 12909 15861 12943 15895
rect 13001 15861 13035 15895
rect 13921 15861 13955 15895
rect 14657 15861 14691 15895
rect 21833 15861 21867 15895
rect 26985 15861 27019 15895
rect 4813 15657 4847 15691
rect 5641 15657 5675 15691
rect 10149 15657 10183 15691
rect 16405 15657 16439 15691
rect 17877 15657 17911 15691
rect 20361 15657 20395 15691
rect 22477 15657 22511 15691
rect 23489 15657 23523 15691
rect 28733 15657 28767 15691
rect 15301 15589 15335 15623
rect 6193 15521 6227 15555
rect 15393 15521 15427 15555
rect 17049 15521 17083 15555
rect 25881 15521 25915 15555
rect 3801 15453 3835 15487
rect 4077 15453 4111 15487
rect 6469 15453 6503 15487
rect 11253 15453 11287 15487
rect 15209 15453 15243 15487
rect 15485 15453 15519 15487
rect 16773 15453 16807 15487
rect 18061 15453 18095 15487
rect 19257 15453 19291 15487
rect 24593 15453 24627 15487
rect 25237 15453 25271 15487
rect 25421 15453 25455 15487
rect 27261 15453 27295 15487
rect 3893 15385 3927 15419
rect 4261 15385 4295 15419
rect 15669 15385 15703 15419
rect 18245 15385 18279 15419
rect 10701 15317 10735 15351
rect 12173 15317 12207 15351
rect 16865 15317 16899 15351
rect 24685 15317 24719 15351
rect 25237 15317 25271 15351
rect 27537 15317 27571 15351
rect 3801 15113 3835 15147
rect 5457 15113 5491 15147
rect 6469 15113 6503 15147
rect 11897 15113 11931 15147
rect 16773 15113 16807 15147
rect 17141 15113 17175 15147
rect 24501 15113 24535 15147
rect 27353 15113 27387 15147
rect 5089 15045 5123 15079
rect 5289 15045 5323 15079
rect 7573 15045 7607 15079
rect 9873 15045 9907 15079
rect 13645 15045 13679 15079
rect 15117 15045 15151 15079
rect 20085 15045 20119 15079
rect 3617 14977 3651 15011
rect 3801 14977 3835 15011
rect 4629 14977 4663 15011
rect 6837 14977 6871 15011
rect 7941 14977 7975 15011
rect 9689 14977 9723 15011
rect 9965 14977 9999 15011
rect 10057 14977 10091 15011
rect 10701 14977 10735 15011
rect 10793 14977 10827 15011
rect 10977 14977 11011 15011
rect 11713 14977 11747 15011
rect 11989 14977 12023 15011
rect 13553 14977 13587 15011
rect 14013 14977 14047 15011
rect 14381 14977 14415 15011
rect 14565 14977 14599 15011
rect 17233 14977 17267 15011
rect 17969 14977 18003 15011
rect 18245 14977 18279 15011
rect 20637 14977 20671 15011
rect 20729 14977 20763 15011
rect 20913 14977 20947 15011
rect 28181 14977 28215 15011
rect 4537 14909 4571 14943
rect 6929 14909 6963 14943
rect 14105 14909 14139 14943
rect 17325 14909 17359 14943
rect 18797 14909 18831 14943
rect 20821 14909 20855 14943
rect 21097 14909 21131 14943
rect 24593 14909 24627 14943
rect 24685 14909 24719 14943
rect 27445 14909 27479 14943
rect 27537 14909 27571 14943
rect 4261 14841 4295 14875
rect 18061 14841 18095 14875
rect 26985 14841 27019 14875
rect 4629 14773 4663 14807
rect 5273 14773 5307 14807
rect 9229 14773 9263 14807
rect 10241 14773 10275 14807
rect 10977 14773 11011 14807
rect 11529 14773 11563 14807
rect 24133 14773 24167 14807
rect 28365 14773 28399 14807
rect 5273 14569 5307 14603
rect 6561 14569 6595 14603
rect 7389 14569 7423 14603
rect 9505 14569 9539 14603
rect 10701 14569 10735 14603
rect 14105 14569 14139 14603
rect 18245 14569 18279 14603
rect 18429 14569 18463 14603
rect 19717 14569 19751 14603
rect 19809 14569 19843 14603
rect 21557 14569 21591 14603
rect 23213 14569 23247 14603
rect 26893 14569 26927 14603
rect 14381 14501 14415 14535
rect 2237 14433 2271 14467
rect 5365 14433 5399 14467
rect 19901 14433 19935 14467
rect 20637 14433 20671 14467
rect 20821 14433 20855 14467
rect 23765 14433 23799 14467
rect 24409 14433 24443 14467
rect 25053 14433 25087 14467
rect 27997 14433 28031 14467
rect 28641 14433 28675 14467
rect 2145 14365 2179 14399
rect 4353 14365 4387 14399
rect 4537 14365 4571 14399
rect 4629 14365 4663 14399
rect 5089 14365 5123 14399
rect 5181 14365 5215 14399
rect 6469 14365 6503 14399
rect 6561 14365 6595 14399
rect 7113 14365 7147 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 10425 14365 10459 14399
rect 10517 14365 10551 14399
rect 11345 14365 11379 14399
rect 11621 14365 11655 14399
rect 14289 14365 14323 14399
rect 14473 14365 14507 14399
rect 14565 14365 14599 14399
rect 15577 14365 15611 14399
rect 15945 14365 15979 14399
rect 17877 14365 17911 14399
rect 18245 14365 18279 14399
rect 19625 14365 19659 14399
rect 20913 14365 20947 14399
rect 23673 14365 23707 14399
rect 23857 14365 23891 14399
rect 24567 14365 24601 14399
rect 24869 14365 24903 14399
rect 27813 14365 27847 14399
rect 2881 14297 2915 14331
rect 8033 14297 8067 14331
rect 9137 14297 9171 14331
rect 9321 14297 9355 14331
rect 12081 14297 12115 14331
rect 17417 14297 17451 14331
rect 20453 14297 20487 14331
rect 21525 14297 21559 14331
rect 21741 14297 21775 14331
rect 24685 14297 24719 14331
rect 24777 14297 24811 14331
rect 26433 14297 26467 14331
rect 27905 14297 27939 14331
rect 1777 14229 1811 14263
rect 4169 14229 4203 14263
rect 6193 14229 6227 14263
rect 7573 14229 7607 14263
rect 11161 14229 11195 14263
rect 11529 14229 11563 14263
rect 21373 14229 21407 14263
rect 27445 14229 27479 14263
rect 4261 14025 4295 14059
rect 4905 14025 4939 14059
rect 5457 14025 5491 14059
rect 8861 14025 8895 14059
rect 10609 14025 10643 14059
rect 15577 14025 15611 14059
rect 19809 14025 19843 14059
rect 28641 14025 28675 14059
rect 6929 13957 6963 13991
rect 7573 13957 7607 13991
rect 12633 13957 12667 13991
rect 24501 13957 24535 13991
rect 24593 13957 24627 13991
rect 27445 13957 27479 13991
rect 1961 13889 1995 13923
rect 3709 13889 3743 13923
rect 4169 13889 4203 13923
rect 6837 13889 6871 13923
rect 9045 13889 9079 13923
rect 9229 13889 9263 13923
rect 10241 13889 10275 13923
rect 12081 13889 12115 13923
rect 15485 13889 15519 13923
rect 15669 13889 15703 13923
rect 19717 13889 19751 13923
rect 19901 13889 19935 13923
rect 20729 13889 20763 13923
rect 22937 13889 22971 13923
rect 23121 13889 23155 13923
rect 24409 13889 24443 13923
rect 24711 13889 24745 13923
rect 24869 13889 24903 13923
rect 27721 13889 27755 13923
rect 28457 13889 28491 13923
rect 1869 13821 1903 13855
rect 10149 13821 10183 13855
rect 10333 13821 10367 13855
rect 10425 13821 10459 13855
rect 19165 13821 19199 13855
rect 20821 13821 20855 13855
rect 27445 13821 27479 13855
rect 11529 13753 11563 13787
rect 27629 13753 27663 13787
rect 2237 13685 2271 13719
rect 20453 13685 20487 13719
rect 23029 13685 23063 13719
rect 24225 13685 24259 13719
rect 10333 13481 10367 13515
rect 10793 13481 10827 13515
rect 25697 13481 25731 13515
rect 26525 13481 26559 13515
rect 28365 13481 28399 13515
rect 19349 13413 19383 13447
rect 20269 13413 20303 13447
rect 22753 13413 22787 13447
rect 25053 13413 25087 13447
rect 8953 13345 8987 13379
rect 21465 13345 21499 13379
rect 1685 13277 1719 13311
rect 7757 13277 7791 13311
rect 7941 13277 7975 13311
rect 8309 13277 8343 13311
rect 12633 13277 12667 13311
rect 12817 13277 12851 13311
rect 21189 13277 21223 13311
rect 21373 13277 21407 13311
rect 22937 13277 22971 13311
rect 23121 13277 23155 13311
rect 24409 13277 24443 13311
rect 25605 13277 25639 13311
rect 25789 13277 25823 13311
rect 26433 13277 26467 13311
rect 26617 13277 26651 13311
rect 9689 13209 9723 13243
rect 11345 13209 11379 13243
rect 1501 13141 1535 13175
rect 2237 13141 2271 13175
rect 7941 13141 7975 13175
rect 12725 13141 12759 13175
rect 15853 13141 15887 13175
rect 21005 13141 21039 13175
rect 23029 13141 23063 13175
rect 23305 13141 23339 13175
rect 24501 13141 24535 13175
rect 27813 13141 27847 13175
rect 7481 12937 7515 12971
rect 10333 12937 10367 12971
rect 14657 12937 14691 12971
rect 17509 12937 17543 12971
rect 20177 12937 20211 12971
rect 20729 12937 20763 12971
rect 23949 12937 23983 12971
rect 25329 12937 25363 12971
rect 27261 12937 27295 12971
rect 27629 12937 27663 12971
rect 8401 12869 8435 12903
rect 11989 12869 12023 12903
rect 18061 12869 18095 12903
rect 20913 12869 20947 12903
rect 5825 12801 5859 12835
rect 6377 12801 6411 12835
rect 7113 12801 7147 12835
rect 8033 12801 8067 12835
rect 8309 12801 8343 12835
rect 8861 12801 8895 12835
rect 9045 12801 9079 12835
rect 10509 12823 10543 12857
rect 10609 12801 10643 12835
rect 10793 12801 10827 12835
rect 10885 12801 10919 12835
rect 13001 12801 13035 12835
rect 13461 12801 13495 12835
rect 13645 12801 13679 12835
rect 14565 12801 14599 12835
rect 14749 12801 14783 12835
rect 15301 12801 15335 12835
rect 16957 12801 16991 12835
rect 19073 12801 19107 12835
rect 19165 12801 19199 12835
rect 19349 12801 19383 12835
rect 19441 12801 19475 12835
rect 21097 12801 21131 12835
rect 23213 12801 23247 12835
rect 23305 12801 23339 12835
rect 23949 12801 23983 12835
rect 24133 12801 24167 12835
rect 24961 12801 24995 12835
rect 25145 12801 25179 12835
rect 25421 12801 25455 12835
rect 28457 12801 28491 12835
rect 7205 12733 7239 12767
rect 15393 12733 15427 12767
rect 16681 12733 16715 12767
rect 23489 12733 23523 12767
rect 27721 12733 27755 12767
rect 27813 12733 27847 12767
rect 16773 12665 16807 12699
rect 16865 12665 16899 12699
rect 19625 12665 19659 12699
rect 23397 12665 23431 12699
rect 5733 12597 5767 12631
rect 8953 12597 8987 12631
rect 9781 12597 9815 12631
rect 13553 12597 13587 12631
rect 15301 12597 15335 12631
rect 15669 12597 15703 12631
rect 18521 12597 18555 12631
rect 28641 12597 28675 12631
rect 7481 12393 7515 12427
rect 12081 12393 12115 12427
rect 19625 12393 19659 12427
rect 26157 12393 26191 12427
rect 5089 12325 5123 12359
rect 5825 12325 5859 12359
rect 10517 12325 10551 12359
rect 11069 12325 11103 12359
rect 14197 12325 14231 12359
rect 15117 12325 15151 12359
rect 26893 12325 26927 12359
rect 2053 12257 2087 12291
rect 9413 12257 9447 12291
rect 14381 12257 14415 12291
rect 14841 12257 14875 12291
rect 20085 12257 20119 12291
rect 25513 12257 25547 12291
rect 27997 12257 28031 12291
rect 2145 12189 2179 12223
rect 4353 12189 4387 12223
rect 4629 12189 4663 12223
rect 5273 12189 5307 12223
rect 5365 12189 5399 12223
rect 5825 12189 5859 12223
rect 5917 12189 5951 12223
rect 7113 12189 7147 12223
rect 7941 12189 7975 12223
rect 8125 12189 8159 12223
rect 9873 12189 9907 12223
rect 9966 12189 10000 12223
rect 10241 12189 10275 12223
rect 10338 12189 10372 12223
rect 11253 12189 11287 12223
rect 11345 12189 11379 12223
rect 11529 12189 11563 12223
rect 11621 12167 11655 12201
rect 12265 12189 12299 12223
rect 12357 12189 12391 12223
rect 12541 12189 12575 12223
rect 12633 12189 12667 12223
rect 13369 12189 13403 12223
rect 13553 12189 13587 12223
rect 14105 12189 14139 12223
rect 15025 12189 15059 12223
rect 15209 12189 15243 12223
rect 15301 12189 15335 12223
rect 16037 12189 16071 12223
rect 16221 12189 16255 12223
rect 16313 12189 16347 12223
rect 16405 12189 16439 12223
rect 19441 12189 19475 12223
rect 19625 12189 19659 12223
rect 25237 12189 25271 12223
rect 27813 12189 27847 12223
rect 4537 12121 4571 12155
rect 5089 12121 5123 12155
rect 6101 12121 6135 12155
rect 7297 12121 7331 12155
rect 8309 12121 8343 12155
rect 10149 12121 10183 12155
rect 21189 12121 21223 12155
rect 26709 12121 26743 12155
rect 27721 12121 27755 12155
rect 28549 12121 28583 12155
rect 2513 12053 2547 12087
rect 4169 12053 4203 12087
rect 6653 12053 6687 12087
rect 13461 12053 13495 12087
rect 14381 12053 14415 12087
rect 16681 12053 16715 12087
rect 17785 12053 17819 12087
rect 18613 12053 18647 12087
rect 19257 12053 19291 12087
rect 24869 12053 24903 12087
rect 25329 12053 25363 12087
rect 27353 12053 27387 12087
rect 3157 11849 3191 11883
rect 5457 11849 5491 11883
rect 6377 11849 6411 11883
rect 7297 11849 7331 11883
rect 9229 11849 9263 11883
rect 10885 11849 10919 11883
rect 11529 11849 11563 11883
rect 14565 11849 14599 11883
rect 24501 11849 24535 11883
rect 27261 11849 27295 11883
rect 27629 11849 27663 11883
rect 28457 11849 28491 11883
rect 8677 11781 8711 11815
rect 10425 11781 10459 11815
rect 11681 11781 11715 11815
rect 11897 11781 11931 11815
rect 22109 11781 22143 11815
rect 22293 11781 22327 11815
rect 2329 11713 2363 11747
rect 2605 11713 2639 11747
rect 4997 11713 5031 11747
rect 7297 11713 7331 11747
rect 7481 11713 7515 11747
rect 12817 11713 12851 11747
rect 13001 11713 13035 11747
rect 13093 11713 13127 11747
rect 13277 11713 13311 11747
rect 17049 11713 17083 11747
rect 17325 11713 17359 11747
rect 18429 11713 18463 11747
rect 19257 11713 19291 11747
rect 20545 11713 20579 11747
rect 20637 11713 20671 11747
rect 20821 11713 20855 11747
rect 20913 11713 20947 11747
rect 23029 11713 23063 11747
rect 23213 11713 23247 11747
rect 23857 11713 23891 11747
rect 24041 11713 24075 11747
rect 24685 11713 24719 11747
rect 24777 11713 24811 11747
rect 24961 11713 24995 11747
rect 25053 11713 25087 11747
rect 19165 11645 19199 11679
rect 21097 11645 21131 11679
rect 22477 11645 22511 11679
rect 23397 11645 23431 11679
rect 27721 11645 27755 11679
rect 27905 11645 27939 11679
rect 12909 11577 12943 11611
rect 17509 11577 17543 11611
rect 19257 11577 19291 11611
rect 4537 11509 4571 11543
rect 4721 11509 4755 11543
rect 7941 11509 7975 11543
rect 9873 11509 9907 11543
rect 11713 11509 11747 11543
rect 12633 11509 12667 11543
rect 13737 11509 13771 11543
rect 20085 11509 20119 11543
rect 23949 11509 23983 11543
rect 1777 11305 1811 11339
rect 17233 11305 17267 11339
rect 18337 11305 18371 11339
rect 19257 11305 19291 11339
rect 19717 11305 19751 11339
rect 21281 11305 21315 11339
rect 22661 11305 22695 11339
rect 24501 11305 24535 11339
rect 27629 11305 27663 11339
rect 27721 11305 27755 11339
rect 4537 11237 4571 11271
rect 18153 11237 18187 11271
rect 20729 11237 20763 11271
rect 23213 11237 23247 11271
rect 2237 11169 2271 11203
rect 4629 11169 4663 11203
rect 8033 11169 8067 11203
rect 8217 11169 8251 11203
rect 9045 11169 9079 11203
rect 10425 11169 10459 11203
rect 10977 11169 11011 11203
rect 12909 11169 12943 11203
rect 13001 11169 13035 11203
rect 14473 11169 14507 11203
rect 19349 11169 19383 11203
rect 21833 11169 21867 11203
rect 27813 11169 27847 11203
rect 2145 11101 2179 11135
rect 4261 11101 4295 11135
rect 4353 11101 4387 11135
rect 7941 11101 7975 11135
rect 8125 11101 8159 11135
rect 8953 11101 8987 11135
rect 9137 11101 9171 11135
rect 13093 11101 13127 11135
rect 13185 11101 13219 11135
rect 14197 11101 14231 11135
rect 14289 11101 14323 11135
rect 14381 11101 14415 11135
rect 17141 11101 17175 11135
rect 17325 11101 17359 11135
rect 18337 11101 18371 11135
rect 18429 11101 18463 11135
rect 19257 11101 19291 11135
rect 19533 11101 19567 11135
rect 27537 11101 27571 11135
rect 2881 11033 2915 11067
rect 7205 11033 7239 11067
rect 9597 11033 9631 11067
rect 11713 11033 11747 11067
rect 16589 11033 16623 11067
rect 18613 11033 18647 11067
rect 20177 11033 20211 11067
rect 4445 10965 4479 10999
rect 7757 10965 7791 10999
rect 12725 10965 12759 10999
rect 14657 10965 14691 10999
rect 1501 10761 1535 10795
rect 5657 10761 5691 10795
rect 5825 10761 5859 10795
rect 11529 10761 11563 10795
rect 14013 10761 14047 10795
rect 17325 10761 17359 10795
rect 18245 10761 18279 10795
rect 20637 10761 20671 10795
rect 25605 10761 25639 10795
rect 27629 10761 27663 10795
rect 5457 10693 5491 10727
rect 23673 10693 23707 10727
rect 1685 10625 1719 10659
rect 4629 10625 4663 10659
rect 6377 10625 6411 10659
rect 7941 10625 7975 10659
rect 8309 10625 8343 10659
rect 8677 10625 8711 10659
rect 9045 10625 9079 10659
rect 9505 10625 9539 10659
rect 13277 10625 13311 10659
rect 13461 10625 13495 10659
rect 13645 10625 13679 10659
rect 14565 10625 14599 10659
rect 17233 10625 17267 10659
rect 17417 10625 17451 10659
rect 18245 10625 18279 10659
rect 18429 10625 18463 10659
rect 19717 10625 19751 10659
rect 21097 10625 21131 10659
rect 21833 10625 21867 10659
rect 21925 10625 21959 10659
rect 22109 10625 22143 10659
rect 22569 10625 22603 10659
rect 22753 10625 22787 10659
rect 23305 10625 23339 10659
rect 23489 10625 23523 10659
rect 24133 10625 24167 10659
rect 24317 10625 24351 10659
rect 24869 10625 24903 10659
rect 25053 10625 25087 10659
rect 25421 10625 25455 10659
rect 26985 10625 27019 10659
rect 27169 10625 27203 10659
rect 27905 10625 27939 10659
rect 4537 10557 4571 10591
rect 4721 10557 4755 10591
rect 4813 10557 4847 10591
rect 19809 10557 19843 10591
rect 19993 10557 20027 10591
rect 20729 10557 20763 10591
rect 20821 10557 20855 10591
rect 23213 10557 23247 10591
rect 25145 10557 25179 10591
rect 25237 10557 25271 10591
rect 27629 10557 27663 10591
rect 9413 10489 9447 10523
rect 19349 10489 19383 10523
rect 21833 10489 21867 10523
rect 24225 10489 24259 10523
rect 27077 10489 27111 10523
rect 2513 10421 2547 10455
rect 4997 10421 5031 10455
rect 5641 10421 5675 10455
rect 12817 10421 12851 10455
rect 13553 10421 13587 10455
rect 13737 10421 13771 10455
rect 21005 10421 21039 10455
rect 22569 10421 22603 10455
rect 27813 10421 27847 10455
rect 9045 10217 9079 10251
rect 13001 10217 13035 10251
rect 17417 10217 17451 10251
rect 19993 10217 20027 10251
rect 20913 10217 20947 10251
rect 22293 10217 22327 10251
rect 24409 10217 24443 10251
rect 25329 10217 25363 10251
rect 10977 10149 11011 10183
rect 23213 10149 23247 10183
rect 25421 10149 25455 10183
rect 4813 10081 4847 10115
rect 7665 10081 7699 10115
rect 11437 10081 11471 10115
rect 18061 10081 18095 10115
rect 21833 10081 21867 10115
rect 25237 10081 25271 10115
rect 27077 10081 27111 10115
rect 28181 10081 28215 10115
rect 28273 10081 28307 10115
rect 4537 10013 4571 10047
rect 7573 10013 7607 10047
rect 8953 10013 8987 10047
rect 10333 10013 10367 10047
rect 10517 10013 10551 10047
rect 10793 10013 10827 10047
rect 12357 10013 12391 10047
rect 12450 10013 12484 10047
rect 12822 10013 12856 10047
rect 14657 10013 14691 10047
rect 17877 10013 17911 10047
rect 19349 10013 19383 10047
rect 20545 10013 20579 10047
rect 21373 10013 21407 10047
rect 21649 10013 21683 10047
rect 23581 10013 23615 10047
rect 24409 10013 24443 10047
rect 24501 10013 24535 10047
rect 25513 10013 25547 10047
rect 26893 10013 26927 10047
rect 28089 10013 28123 10047
rect 12633 9945 12667 9979
rect 12725 9945 12759 9979
rect 14105 9945 14139 9979
rect 16405 9945 16439 9979
rect 20729 9945 20763 9979
rect 21465 9945 21499 9979
rect 22477 9945 22511 9979
rect 22661 9945 22695 9979
rect 23397 9945 23431 9979
rect 25973 9945 26007 9979
rect 2605 9877 2639 9911
rect 7941 9877 7975 9911
rect 13461 9877 13495 9911
rect 16865 9877 16899 9911
rect 17785 9877 17819 9911
rect 18705 9877 18739 9911
rect 24777 9877 24811 9911
rect 26525 9877 26559 9911
rect 26985 9877 27019 9911
rect 27721 9877 27755 9911
rect 10977 9673 11011 9707
rect 12357 9673 12391 9707
rect 17417 9673 17451 9707
rect 21833 9673 21867 9707
rect 22937 9673 22971 9707
rect 27813 9673 27847 9707
rect 2145 9605 2179 9639
rect 3157 9605 3191 9639
rect 7297 9605 7331 9639
rect 8033 9605 8067 9639
rect 14381 9605 14415 9639
rect 15853 9605 15887 9639
rect 17877 9605 17911 9639
rect 18705 9605 18739 9639
rect 23673 9605 23707 9639
rect 24317 9605 24351 9639
rect 24961 9605 24995 9639
rect 2329 9537 2363 9571
rect 3341 9537 3375 9571
rect 4353 9537 4387 9571
rect 7113 9537 7147 9571
rect 7941 9537 7975 9571
rect 8217 9537 8251 9571
rect 9045 9537 9079 9571
rect 9137 9537 9171 9571
rect 9321 9537 9355 9571
rect 10609 9537 10643 9571
rect 12909 9537 12943 9571
rect 15117 9537 15151 9571
rect 15301 9537 15335 9571
rect 17785 9537 17819 9571
rect 20453 9537 20487 9571
rect 20913 9537 20947 9571
rect 23857 9537 23891 9571
rect 25237 9537 25271 9571
rect 25329 9537 25363 9571
rect 25421 9537 25455 9571
rect 25605 9537 25639 9571
rect 27629 9537 27663 9571
rect 28733 9537 28767 9571
rect 10333 9469 10367 9503
rect 10517 9469 10551 9503
rect 12633 9469 12667 9503
rect 18061 9469 18095 9503
rect 23489 9469 23523 9503
rect 27353 9469 27387 9503
rect 3893 9401 3927 9435
rect 27445 9401 27479 9435
rect 2513 9333 2547 9367
rect 2973 9333 3007 9367
rect 4445 9333 4479 9367
rect 8401 9333 8435 9367
rect 11529 9333 11563 9367
rect 12541 9333 12575 9367
rect 13461 9333 13495 9367
rect 15301 9333 15335 9367
rect 16957 9333 16991 9367
rect 19257 9333 19291 9367
rect 22477 9333 22511 9367
rect 28549 9333 28583 9367
rect 1961 9129 1995 9163
rect 3893 9129 3927 9163
rect 4813 9129 4847 9163
rect 5549 9129 5583 9163
rect 7021 9129 7055 9163
rect 8309 9129 8343 9163
rect 9689 9129 9723 9163
rect 11069 9129 11103 9163
rect 15669 9129 15703 9163
rect 23121 9129 23155 9163
rect 24961 9129 24995 9163
rect 27261 9129 27295 9163
rect 27997 9129 28031 9163
rect 28733 9129 28767 9163
rect 13001 9061 13035 9095
rect 21281 9061 21315 9095
rect 2421 8993 2455 9027
rect 4905 8993 4939 9027
rect 6561 8993 6595 9027
rect 10241 8993 10275 9027
rect 25605 8993 25639 9027
rect 2329 8925 2363 8959
rect 4537 8925 4571 8959
rect 7205 8925 7239 8959
rect 7297 8925 7331 8959
rect 7481 8925 7515 8959
rect 7573 8925 7607 8959
rect 9505 8925 9539 8959
rect 9689 8925 9723 8959
rect 14565 8925 14599 8959
rect 14713 8925 14747 8959
rect 15030 8925 15064 8959
rect 17049 8925 17083 8959
rect 17693 8925 17727 8959
rect 25329 8925 25363 8959
rect 5365 8857 5399 8891
rect 14841 8857 14875 8891
rect 14933 8857 14967 8891
rect 17877 8857 17911 8891
rect 4629 8789 4663 8823
rect 4721 8789 4755 8823
rect 5565 8789 5599 8823
rect 5733 8789 5767 8823
rect 9045 8789 9079 8823
rect 13553 8789 13587 8823
rect 15209 8789 15243 8823
rect 17509 8789 17543 8823
rect 23673 8789 23707 8823
rect 25421 8789 25455 8823
rect 4629 8585 4663 8619
rect 6377 8585 6411 8619
rect 7481 8585 7515 8619
rect 11529 8585 11563 8619
rect 14013 8585 14047 8619
rect 18061 8585 18095 8619
rect 21189 8585 21223 8619
rect 23029 8585 23063 8619
rect 23673 8585 23707 8619
rect 25237 8585 25271 8619
rect 25605 8585 25639 8619
rect 26985 8585 27019 8619
rect 27353 8585 27387 8619
rect 1593 8517 1627 8551
rect 5733 8517 5767 8551
rect 8033 8517 8067 8551
rect 10149 8517 10183 8551
rect 14933 8517 14967 8551
rect 20085 8517 20119 8551
rect 21925 8517 21959 8551
rect 2605 8449 2639 8483
rect 2881 8449 2915 8483
rect 4997 8449 5031 8483
rect 8217 8449 8251 8483
rect 13829 8449 13863 8483
rect 14013 8449 14047 8483
rect 14657 8449 14691 8483
rect 14749 8449 14783 8483
rect 15393 8449 15427 8483
rect 15485 8449 15519 8483
rect 15669 8449 15703 8483
rect 17233 8449 17267 8483
rect 17325 8449 17359 8483
rect 17417 8449 17451 8483
rect 17601 8449 17635 8483
rect 20269 8449 20303 8483
rect 20361 8449 20395 8483
rect 20545 8449 20579 8483
rect 20637 8449 20671 8483
rect 22385 8449 22419 8483
rect 2789 8381 2823 8415
rect 4813 8381 4847 8415
rect 4905 8381 4939 8415
rect 5089 8381 5123 8415
rect 9321 8381 9355 8415
rect 9597 8381 9631 8415
rect 13093 8381 13127 8415
rect 22293 8381 22327 8415
rect 25697 8381 25731 8415
rect 25789 8381 25823 8415
rect 27445 8381 27479 8415
rect 27537 8381 27571 8415
rect 14473 8313 14507 8347
rect 15669 8313 15703 8347
rect 1869 8245 1903 8279
rect 2421 8245 2455 8279
rect 2789 8245 2823 8279
rect 3433 8245 3467 8279
rect 14933 8245 14967 8279
rect 16957 8245 16991 8279
rect 22385 8245 22419 8279
rect 22569 8245 22603 8279
rect 1501 8041 1535 8075
rect 2237 8041 2271 8075
rect 8953 8041 8987 8075
rect 11253 8041 11287 8075
rect 15485 8041 15519 8075
rect 17141 8041 17175 8075
rect 21005 8041 21039 8075
rect 22477 8041 22511 8075
rect 25973 8041 26007 8075
rect 27169 8041 27203 8075
rect 2145 7973 2179 8007
rect 6009 7973 6043 8007
rect 14105 7973 14139 8007
rect 2329 7905 2363 7939
rect 4721 7905 4755 7939
rect 5089 7905 5123 7939
rect 6193 7905 6227 7939
rect 10793 7905 10827 7939
rect 15025 7905 15059 7939
rect 20545 7905 20579 7939
rect 22017 7905 22051 7939
rect 22109 7905 22143 7939
rect 26617 7905 26651 7939
rect 27721 7905 27755 7939
rect 1961 7837 1995 7871
rect 4629 7837 4663 7871
rect 4997 7837 5031 7871
rect 9137 7837 9171 7871
rect 9229 7837 9263 7871
rect 9413 7837 9447 7871
rect 9505 7837 9539 7871
rect 10885 7837 10919 7871
rect 14841 7837 14875 7871
rect 15664 7837 15698 7871
rect 15761 7837 15795 7871
rect 15981 7837 16015 7871
rect 16129 7837 16163 7871
rect 19257 7837 19291 7871
rect 19441 7837 19475 7871
rect 21281 7837 21315 7871
rect 22201 7837 22235 7871
rect 22292 7837 22326 7871
rect 22937 7837 22971 7871
rect 24409 7837 24443 7871
rect 27537 7837 27571 7871
rect 5273 7769 5307 7803
rect 5733 7769 5767 7803
rect 13553 7769 13587 7803
rect 15853 7769 15887 7803
rect 16681 7769 16715 7803
rect 21005 7769 21039 7803
rect 26341 7769 26375 7803
rect 27629 7769 27663 7803
rect 28457 7769 28491 7803
rect 28641 7769 28675 7803
rect 2053 7701 2087 7735
rect 2973 7701 3007 7735
rect 4905 7701 4939 7735
rect 10149 7701 10183 7735
rect 11713 7701 11747 7735
rect 13001 7701 13035 7735
rect 14657 7701 14691 7735
rect 17877 7701 17911 7735
rect 18613 7701 18647 7735
rect 19349 7701 19383 7735
rect 19993 7701 20027 7735
rect 21189 7701 21223 7735
rect 23581 7701 23615 7735
rect 26433 7701 26467 7735
rect 5365 7497 5399 7531
rect 7941 7497 7975 7531
rect 9229 7497 9263 7531
rect 9781 7497 9815 7531
rect 12265 7497 12299 7531
rect 14565 7497 14599 7531
rect 18337 7497 18371 7531
rect 19441 7497 19475 7531
rect 21925 7497 21959 7531
rect 25973 7497 26007 7531
rect 27261 7497 27295 7531
rect 27721 7497 27755 7531
rect 10701 7429 10735 7463
rect 12633 7429 12667 7463
rect 14197 7429 14231 7463
rect 14397 7429 14431 7463
rect 19717 7429 19751 7463
rect 19809 7429 19843 7463
rect 21189 7429 21223 7463
rect 28733 7429 28767 7463
rect 4997 7361 5031 7395
rect 6469 7361 6503 7395
rect 6561 7361 6595 7395
rect 8217 7361 8251 7395
rect 8769 7361 8803 7395
rect 9045 7361 9079 7395
rect 10333 7361 10367 7395
rect 10426 7361 10460 7395
rect 10609 7361 10643 7395
rect 10798 7361 10832 7395
rect 12403 7361 12437 7395
rect 12541 7361 12575 7395
rect 12761 7361 12795 7395
rect 12909 7361 12943 7395
rect 16957 7361 16991 7395
rect 17233 7361 17267 7395
rect 17785 7361 17819 7395
rect 18521 7361 18555 7395
rect 18797 7361 18831 7395
rect 18981 7361 19015 7395
rect 19620 7361 19654 7395
rect 19992 7361 20026 7395
rect 20085 7361 20119 7395
rect 22845 7361 22879 7395
rect 23489 7361 23523 7395
rect 23581 7361 23615 7395
rect 25697 7361 25731 7395
rect 26985 7361 27019 7395
rect 27997 7361 28031 7395
rect 4905 7293 4939 7327
rect 5089 7293 5123 7327
rect 5181 7293 5215 7327
rect 7389 7293 7423 7327
rect 7941 7293 7975 7327
rect 8125 7293 8159 7327
rect 8953 7293 8987 7327
rect 13369 7293 13403 7327
rect 16681 7293 16715 7327
rect 20637 7293 20671 7327
rect 22753 7293 22787 7327
rect 25973 7293 26007 7327
rect 27261 7293 27295 7327
rect 27721 7293 27755 7327
rect 8861 7225 8895 7259
rect 11713 7225 11747 7259
rect 15301 7225 15335 7259
rect 10977 7157 11011 7191
rect 14381 7157 14415 7191
rect 15853 7157 15887 7191
rect 22477 7157 22511 7191
rect 22845 7157 22879 7191
rect 23305 7157 23339 7191
rect 25789 7157 25823 7191
rect 27077 7157 27111 7191
rect 27905 7157 27939 7191
rect 4353 6953 4387 6987
rect 4905 6953 4939 6987
rect 11805 6953 11839 6987
rect 13185 6953 13219 6987
rect 14105 6953 14139 6987
rect 14473 6953 14507 6987
rect 16865 6953 16899 6987
rect 18705 6953 18739 6987
rect 22109 6953 22143 6987
rect 23489 6953 23523 6987
rect 25697 6953 25731 6987
rect 27353 6953 27387 6987
rect 27813 6953 27847 6987
rect 9413 6885 9447 6919
rect 10517 6885 10551 6919
rect 12725 6885 12759 6919
rect 15945 6885 15979 6919
rect 4261 6817 4295 6851
rect 9505 6817 9539 6851
rect 16957 6817 16991 6851
rect 20729 6817 20763 6851
rect 22661 6817 22695 6851
rect 25145 6817 25179 6851
rect 26801 6817 26835 6851
rect 28273 6817 28307 6851
rect 28365 6817 28399 6851
rect 4353 6749 4387 6783
rect 4813 6749 4847 6783
rect 4997 6749 5031 6783
rect 5825 6749 5859 6783
rect 6009 6749 6043 6783
rect 6285 6749 6319 6783
rect 7021 6749 7055 6783
rect 7205 6749 7239 6783
rect 7665 6749 7699 6783
rect 9321 6749 9355 6783
rect 9586 6749 9620 6783
rect 10333 6749 10367 6783
rect 10425 6749 10459 6783
rect 10609 6749 10643 6783
rect 10793 6749 10827 6783
rect 11253 6749 11287 6783
rect 11345 6749 11379 6783
rect 11529 6749 11563 6783
rect 11621 6749 11655 6783
rect 12449 6749 12483 6783
rect 13185 6749 13219 6783
rect 13369 6749 13403 6783
rect 14105 6749 14139 6783
rect 14197 6749 14231 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 16037 6749 16071 6783
rect 16221 6749 16255 6783
rect 16681 6749 16715 6783
rect 16773 6749 16807 6783
rect 18245 6749 18279 6783
rect 18337 6749 18371 6783
rect 18613 6749 18647 6783
rect 18705 6749 18739 6783
rect 19257 6749 19291 6783
rect 19350 6749 19384 6783
rect 19625 6749 19659 6783
rect 19763 6749 19797 6783
rect 20453 6749 20487 6783
rect 20545 6749 20579 6783
rect 22017 6749 22051 6783
rect 22201 6749 22235 6783
rect 22845 6749 22879 6783
rect 25329 6749 25363 6783
rect 7113 6681 7147 6715
rect 8401 6681 8435 6715
rect 9137 6681 9171 6715
rect 12725 6681 12759 6715
rect 15577 6681 15611 6715
rect 18429 6681 18463 6715
rect 19533 6681 19567 6715
rect 20729 6681 20763 6715
rect 23673 6681 23707 6715
rect 23857 6681 23891 6715
rect 26893 6681 26927 6715
rect 28181 6681 28215 6715
rect 3985 6613 4019 6647
rect 5181 6613 5215 6647
rect 6193 6613 6227 6647
rect 10149 6613 10183 6647
rect 12541 6613 12575 6647
rect 15025 6613 15059 6647
rect 17509 6613 17543 6647
rect 19901 6613 19935 6647
rect 21189 6613 21223 6647
rect 23029 6613 23063 6647
rect 24409 6613 24443 6647
rect 25237 6613 25271 6647
rect 26985 6613 27019 6647
rect 1593 6409 1627 6443
rect 6837 6409 6871 6443
rect 8677 6409 8711 6443
rect 10609 6409 10643 6443
rect 11897 6409 11931 6443
rect 12633 6409 12667 6443
rect 13277 6409 13311 6443
rect 14105 6409 14139 6443
rect 14565 6409 14599 6443
rect 15853 6409 15887 6443
rect 18429 6409 18463 6443
rect 19073 6409 19107 6443
rect 19625 6409 19659 6443
rect 23213 6409 23247 6443
rect 24133 6409 24167 6443
rect 26433 6409 26467 6443
rect 27077 6409 27111 6443
rect 28089 6409 28123 6443
rect 9597 6341 9631 6375
rect 10241 6341 10275 6375
rect 16681 6341 16715 6375
rect 17969 6341 18003 6375
rect 22661 6341 22695 6375
rect 25881 6341 25915 6375
rect 27629 6341 27663 6375
rect 28641 6341 28675 6375
rect 1409 6273 1443 6307
rect 5181 6273 5215 6307
rect 5365 6273 5399 6307
rect 5457 6273 5491 6307
rect 5549 6273 5583 6307
rect 7021 6273 7055 6307
rect 7205 6273 7239 6307
rect 7941 6273 7975 6307
rect 8861 6273 8895 6307
rect 9045 6273 9079 6307
rect 10057 6273 10091 6307
rect 10333 6273 10367 6307
rect 10425 6273 10459 6307
rect 12541 6273 12575 6307
rect 12725 6273 12759 6307
rect 13185 6273 13219 6307
rect 13369 6273 13403 6307
rect 13829 6273 13863 6307
rect 15393 6273 15427 6307
rect 15669 6273 15703 6307
rect 16865 6273 16899 6307
rect 17049 6273 17083 6307
rect 18245 6273 18279 6307
rect 19165 6273 19199 6307
rect 20361 6273 20395 6307
rect 20545 6273 20579 6307
rect 22017 6273 22051 6307
rect 22201 6273 22235 6307
rect 7297 6205 7331 6239
rect 7849 6205 7883 6239
rect 14105 6205 14139 6239
rect 15485 6205 15519 6239
rect 18153 6205 18187 6239
rect 20177 6205 20211 6239
rect 5825 6137 5859 6171
rect 15577 6137 15611 6171
rect 24869 6137 24903 6171
rect 4629 6069 4663 6103
rect 13921 6069 13955 6103
rect 18245 6069 18279 6103
rect 21097 6069 21131 6103
rect 21833 6069 21867 6103
rect 22017 6069 22051 6103
rect 1409 5865 1443 5899
rect 5733 5865 5767 5899
rect 7205 5865 7239 5899
rect 9137 5865 9171 5899
rect 10609 5865 10643 5899
rect 13093 5865 13127 5899
rect 15209 5865 15243 5899
rect 15761 5865 15795 5899
rect 18337 5865 18371 5899
rect 19901 5865 19935 5899
rect 21189 5865 21223 5899
rect 22569 5865 22603 5899
rect 28549 5865 28583 5899
rect 6561 5797 6595 5831
rect 17693 5797 17727 5831
rect 19257 5797 19291 5831
rect 21373 5797 21407 5831
rect 27997 5797 28031 5831
rect 16129 5729 16163 5763
rect 16589 5729 16623 5763
rect 20545 5729 20579 5763
rect 5549 5661 5583 5695
rect 5917 5661 5951 5695
rect 6009 5661 6043 5695
rect 6469 5661 6503 5695
rect 6653 5661 6687 5695
rect 7941 5661 7975 5695
rect 13277 5661 13311 5695
rect 13461 5661 13495 5695
rect 15945 5661 15979 5695
rect 19257 5661 19291 5695
rect 19441 5661 19475 5695
rect 21833 5661 21867 5695
rect 28733 5661 28767 5695
rect 11161 5593 11195 5627
rect 12081 5593 12115 5627
rect 14197 5593 14231 5627
rect 14749 5593 14783 5627
rect 21005 5593 21039 5627
rect 21205 5593 21239 5627
rect 7849 5525 7883 5559
rect 17233 5525 17267 5559
rect 6837 5321 6871 5355
rect 8033 5321 8067 5355
rect 10057 5321 10091 5355
rect 10885 5321 10919 5355
rect 13829 5321 13863 5355
rect 14657 5321 14691 5355
rect 15485 5321 15519 5355
rect 17877 5321 17911 5355
rect 18613 5321 18647 5355
rect 28733 5321 28767 5355
rect 22109 5253 22143 5287
rect 22201 5253 22235 5287
rect 7205 5185 7239 5219
rect 21833 5185 21867 5219
rect 21925 5185 21959 5219
rect 22293 5185 22327 5219
rect 23673 5185 23707 5219
rect 24133 5185 24167 5219
rect 24685 5185 24719 5219
rect 7113 5117 7147 5151
rect 22937 5117 22971 5151
rect 22477 5049 22511 5083
rect 23397 5049 23431 5083
rect 5825 4981 5859 5015
rect 7205 4981 7239 5015
rect 19165 4981 19199 5015
rect 19809 4981 19843 5015
rect 2145 4777 2179 4811
rect 6653 4777 6687 4811
rect 6745 4777 6779 4811
rect 7297 4777 7331 4811
rect 10517 4777 10551 4811
rect 14381 4777 14415 4811
rect 15761 4777 15795 4811
rect 19901 4777 19935 4811
rect 23397 4777 23431 4811
rect 16221 4709 16255 4743
rect 17785 4709 17819 4743
rect 22017 4709 22051 4743
rect 24409 4709 24443 4743
rect 6561 4641 6595 4675
rect 9321 4641 9355 4675
rect 20545 4641 20579 4675
rect 21005 4641 21039 4675
rect 6837 4573 6871 4607
rect 9505 4573 9539 4607
rect 9689 4573 9723 4607
rect 14197 4573 14231 4607
rect 14381 4573 14415 4607
rect 15117 4573 15151 4607
rect 15209 4573 15243 4607
rect 20085 4573 20119 4607
rect 20407 4573 20441 4607
rect 22569 4573 22603 4607
rect 22753 4573 22787 4607
rect 23213 4573 23247 4607
rect 1869 4505 1903 4539
rect 10149 4505 10183 4539
rect 10333 4505 10367 4539
rect 10977 4505 11011 4539
rect 20177 4505 20211 4539
rect 20269 4505 20303 4539
rect 14565 4437 14599 4471
rect 22753 4437 22787 4471
rect 10885 4233 10919 4267
rect 12725 4233 12759 4267
rect 15945 4233 15979 4267
rect 20637 4233 20671 4267
rect 22293 4233 22327 4267
rect 1593 4165 1627 4199
rect 13185 4165 13219 4199
rect 15193 4165 15227 4199
rect 15393 4165 15427 4199
rect 16865 4165 16899 4199
rect 23397 4165 23431 4199
rect 2421 4097 2455 4131
rect 10057 4097 10091 4131
rect 10241 4097 10275 4131
rect 10425 4097 10459 4131
rect 11529 4097 11563 4131
rect 11713 4097 11747 4131
rect 12909 4097 12943 4131
rect 14289 4097 14323 4131
rect 14565 4097 14599 4131
rect 17325 4097 17359 4131
rect 17509 4097 17543 4131
rect 18153 4097 18187 4131
rect 19073 4097 19107 4131
rect 19533 4097 19567 4131
rect 20913 4097 20947 4131
rect 21833 4097 21867 4131
rect 21925 4097 21959 4131
rect 22109 4097 22143 4131
rect 23213 4097 23247 4131
rect 23305 4097 23339 4131
rect 24133 4097 24167 4131
rect 24317 4097 24351 4131
rect 24777 4097 24811 4131
rect 2973 4029 3007 4063
rect 12173 4029 12207 4063
rect 13093 4029 13127 4063
rect 14473 4029 14507 4063
rect 18337 4029 18371 4063
rect 18429 4029 18463 4063
rect 18981 4029 19015 4063
rect 20637 4029 20671 4063
rect 20821 4029 20855 4063
rect 23673 4029 23707 4063
rect 24225 4029 24259 4063
rect 9597 3961 9631 3995
rect 15025 3961 15059 3995
rect 2237 3893 2271 3927
rect 11529 3893 11563 3927
rect 12909 3893 12943 3927
rect 14105 3893 14139 3927
rect 15209 3893 15243 3927
rect 17509 3893 17543 3927
rect 17969 3893 18003 3927
rect 22937 3893 22971 3927
rect 23581 3893 23615 3927
rect 28641 3893 28675 3927
rect 10977 3689 11011 3723
rect 13553 3689 13587 3723
rect 14197 3689 14231 3723
rect 14657 3689 14691 3723
rect 15669 3689 15703 3723
rect 16865 3689 16899 3723
rect 20085 3689 20119 3723
rect 20821 3689 20855 3723
rect 21741 3689 21775 3723
rect 23305 3689 23339 3723
rect 24409 3689 24443 3723
rect 11989 3621 12023 3655
rect 15853 3621 15887 3655
rect 17325 3621 17359 3655
rect 18613 3621 18647 3655
rect 28457 3621 28491 3655
rect 11529 3553 11563 3587
rect 16589 3553 16623 3587
rect 17601 3553 17635 3587
rect 19533 3553 19567 3587
rect 22293 3553 22327 3587
rect 23765 3553 23799 3587
rect 1685 3485 1719 3519
rect 10517 3485 10551 3519
rect 10793 3485 10827 3519
rect 11621 3485 11655 3519
rect 12633 3485 12667 3519
rect 13093 3485 13127 3519
rect 13277 3485 13311 3519
rect 14105 3485 14139 3519
rect 14473 3485 14507 3519
rect 16405 3485 16439 3519
rect 16497 3485 16531 3519
rect 16684 3485 16718 3519
rect 17693 3485 17727 3519
rect 18337 3485 18371 3519
rect 19441 3485 19475 3519
rect 19960 3485 19994 3519
rect 20913 3485 20947 3519
rect 21005 3485 21039 3519
rect 21465 3485 21499 3519
rect 21649 3485 21683 3519
rect 21741 3485 21775 3519
rect 22201 3485 22235 3519
rect 22937 3485 22971 3519
rect 10609 3417 10643 3451
rect 15485 3417 15519 3451
rect 18613 3417 18647 3451
rect 23121 3417 23155 3451
rect 28641 3417 28675 3451
rect 1501 3349 1535 3383
rect 12541 3349 12575 3383
rect 13369 3349 13403 3383
rect 15695 3349 15729 3383
rect 18429 3349 18463 3383
rect 19901 3349 19935 3383
rect 20637 3349 20671 3383
rect 27905 3349 27939 3383
rect 10333 3145 10367 3179
rect 10885 3145 10919 3179
rect 11529 3145 11563 3179
rect 12725 3145 12759 3179
rect 13921 3145 13955 3179
rect 14933 3145 14967 3179
rect 18061 3145 18095 3179
rect 20729 3145 20763 3179
rect 23397 3145 23431 3179
rect 15117 3077 15151 3111
rect 18981 3077 19015 3111
rect 19165 3077 19199 3111
rect 19349 3077 19383 3111
rect 21281 3077 21315 3111
rect 28457 3077 28491 3111
rect 1685 3009 1719 3043
rect 11713 3009 11747 3043
rect 11897 3009 11931 3043
rect 11989 3009 12023 3043
rect 14381 3009 14415 3043
rect 14841 3009 14875 3043
rect 18153 3009 18187 3043
rect 20545 3009 20579 3043
rect 20729 3009 20763 3043
rect 27169 3009 27203 3043
rect 27721 3009 27755 3043
rect 28641 3009 28675 3043
rect 21833 2941 21867 2975
rect 15117 2873 15151 2907
rect 27905 2873 27939 2907
rect 1501 2805 1535 2839
rect 14105 2805 14139 2839
rect 16865 2805 16899 2839
rect 19809 2805 19843 2839
rect 6561 2601 6595 2635
rect 14381 2601 14415 2635
rect 17233 2601 17267 2635
rect 20913 2601 20947 2635
rect 27997 2601 28031 2635
rect 2421 2533 2455 2567
rect 23581 2533 23615 2567
rect 12725 2465 12759 2499
rect 18245 2465 18279 2499
rect 19533 2465 19567 2499
rect 25237 2465 25271 2499
rect 4261 2397 4295 2431
rect 6377 2397 6411 2431
rect 8953 2397 8987 2431
rect 10701 2397 10735 2431
rect 14933 2397 14967 2431
rect 19257 2397 19291 2431
rect 21005 2397 21039 2431
rect 21833 2397 21867 2431
rect 1593 2329 1627 2363
rect 2145 2329 2179 2363
rect 11897 2329 11931 2363
rect 12449 2329 12483 2363
rect 17141 2329 17175 2363
rect 22845 2329 22879 2363
rect 23397 2329 23431 2363
rect 24777 2329 24811 2363
rect 25421 2329 25455 2363
rect 27353 2329 27387 2363
rect 27905 2329 27939 2363
rect 4077 2261 4111 2295
rect 5825 2261 5859 2295
rect 9137 2261 9171 2295
rect 10517 2261 10551 2295
rect 15117 2261 15151 2295
rect 22017 2261 22051 2295
<< metal1 >>
rect 1104 30490 29600 30512
rect 1104 30438 8034 30490
rect 8086 30438 8098 30490
rect 8150 30438 8162 30490
rect 8214 30438 8226 30490
rect 8278 30438 8290 30490
rect 8342 30438 15118 30490
rect 15170 30438 15182 30490
rect 15234 30438 15246 30490
rect 15298 30438 15310 30490
rect 15362 30438 15374 30490
rect 15426 30438 22202 30490
rect 22254 30438 22266 30490
rect 22318 30438 22330 30490
rect 22382 30438 22394 30490
rect 22446 30438 22458 30490
rect 22510 30438 29286 30490
rect 29338 30438 29350 30490
rect 29402 30438 29414 30490
rect 29466 30438 29478 30490
rect 29530 30438 29542 30490
rect 29594 30438 29600 30490
rect 1104 30416 29600 30438
rect 658 30268 664 30320
rect 716 30308 722 30320
rect 1302 30308 1308 30320
rect 716 30280 1308 30308
rect 716 30268 722 30280
rect 1302 30268 1308 30280
rect 1360 30308 1366 30320
rect 1857 30311 1915 30317
rect 1857 30308 1869 30311
rect 1360 30280 1869 30308
rect 1360 30268 1366 30280
rect 1857 30277 1869 30280
rect 1903 30277 1915 30311
rect 1857 30271 1915 30277
rect 2590 30268 2596 30320
rect 2648 30308 2654 30320
rect 2777 30311 2835 30317
rect 2777 30308 2789 30311
rect 2648 30280 2789 30308
rect 2648 30268 2654 30280
rect 2777 30277 2789 30280
rect 2823 30277 2835 30311
rect 2777 30271 2835 30277
rect 7469 30311 7527 30317
rect 7469 30277 7481 30311
rect 7515 30308 7527 30311
rect 13538 30308 13544 30320
rect 7515 30280 12434 30308
rect 13499 30280 13544 30308
rect 7515 30277 7527 30280
rect 7469 30271 7527 30277
rect 5534 30240 5540 30252
rect 5495 30212 5540 30240
rect 5534 30200 5540 30212
rect 5592 30200 5598 30252
rect 6733 30243 6791 30249
rect 6733 30209 6745 30243
rect 6779 30240 6791 30243
rect 7098 30240 7104 30252
rect 6779 30212 7104 30240
rect 6779 30209 6791 30212
rect 6733 30203 6791 30209
rect 7098 30200 7104 30212
rect 7156 30240 7162 30252
rect 7193 30243 7251 30249
rect 7193 30240 7205 30243
rect 7156 30212 7205 30240
rect 7156 30200 7162 30212
rect 7193 30209 7205 30212
rect 7239 30209 7251 30243
rect 7193 30203 7251 30209
rect 7834 30200 7840 30252
rect 7892 30240 7898 30252
rect 9125 30243 9183 30249
rect 9125 30240 9137 30243
rect 7892 30212 9137 30240
rect 7892 30200 7898 30212
rect 9125 30209 9137 30212
rect 9171 30209 9183 30243
rect 9125 30203 9183 30209
rect 11330 30200 11336 30252
rect 11388 30240 11394 30252
rect 11701 30243 11759 30249
rect 11701 30240 11713 30243
rect 11388 30212 11713 30240
rect 11388 30200 11394 30212
rect 11701 30209 11713 30212
rect 11747 30209 11759 30243
rect 12406 30240 12434 30280
rect 13538 30268 13544 30280
rect 13596 30268 13602 30320
rect 15105 30311 15163 30317
rect 15105 30277 15117 30311
rect 15151 30308 15163 30311
rect 15470 30308 15476 30320
rect 15151 30280 15476 30308
rect 15151 30277 15163 30280
rect 15105 30271 15163 30277
rect 15470 30268 15476 30280
rect 15528 30308 15534 30320
rect 15657 30311 15715 30317
rect 15657 30308 15669 30311
rect 15528 30280 15669 30308
rect 15528 30268 15534 30280
rect 15657 30277 15669 30280
rect 15703 30277 15715 30311
rect 15657 30271 15715 30277
rect 13556 30240 13584 30268
rect 14093 30243 14151 30249
rect 14093 30240 14105 30243
rect 12406 30212 13400 30240
rect 13556 30212 14105 30240
rect 11701 30203 11759 30209
rect 13372 30172 13400 30212
rect 14093 30209 14105 30212
rect 14139 30209 14151 30243
rect 14093 30203 14151 30209
rect 18046 30200 18052 30252
rect 18104 30240 18110 30252
rect 18141 30243 18199 30249
rect 18141 30240 18153 30243
rect 18104 30212 18153 30240
rect 18104 30200 18110 30212
rect 18141 30209 18153 30212
rect 18187 30240 18199 30243
rect 19245 30243 19303 30249
rect 19245 30240 19257 30243
rect 18187 30212 19257 30240
rect 18187 30209 18199 30212
rect 18141 30203 18199 30209
rect 19245 30209 19257 30212
rect 19291 30209 19303 30243
rect 19245 30203 19303 30209
rect 19978 30200 19984 30252
rect 20036 30240 20042 30252
rect 20073 30243 20131 30249
rect 20073 30240 20085 30243
rect 20036 30212 20085 30240
rect 20036 30200 20042 30212
rect 20073 30209 20085 30212
rect 20119 30209 20131 30243
rect 20073 30203 20131 30209
rect 21269 30243 21327 30249
rect 21269 30209 21281 30243
rect 21315 30240 21327 30243
rect 21910 30240 21916 30252
rect 21315 30212 21916 30240
rect 21315 30209 21327 30212
rect 21269 30203 21327 30209
rect 21910 30200 21916 30212
rect 21968 30240 21974 30252
rect 22005 30243 22063 30249
rect 22005 30240 22017 30243
rect 21968 30212 22017 30240
rect 21968 30200 21974 30212
rect 22005 30209 22017 30212
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 24486 30200 24492 30252
rect 24544 30240 24550 30252
rect 24581 30243 24639 30249
rect 24581 30240 24593 30243
rect 24544 30212 24593 30240
rect 24544 30200 24550 30212
rect 24581 30209 24593 30212
rect 24627 30209 24639 30243
rect 24581 30203 24639 30209
rect 26326 30200 26332 30252
rect 26384 30240 26390 30252
rect 26973 30243 27031 30249
rect 26973 30240 26985 30243
rect 26384 30212 26985 30240
rect 26384 30200 26390 30212
rect 26973 30209 26985 30212
rect 27019 30209 27031 30243
rect 26973 30203 27031 30209
rect 27614 30200 27620 30252
rect 27672 30240 27678 30252
rect 27709 30243 27767 30249
rect 27709 30240 27721 30243
rect 27672 30212 27721 30240
rect 27672 30200 27678 30212
rect 27709 30209 27721 30212
rect 27755 30209 27767 30243
rect 27709 30203 27767 30209
rect 28258 30200 28264 30252
rect 28316 30240 28322 30252
rect 28445 30243 28503 30249
rect 28445 30240 28457 30243
rect 28316 30212 28457 30240
rect 28316 30200 28322 30212
rect 28445 30209 28457 30212
rect 28491 30209 28503 30243
rect 28445 30203 28503 30209
rect 13906 30172 13912 30184
rect 6886 30144 13308 30172
rect 13372 30144 13912 30172
rect 2038 30104 2044 30116
rect 1999 30076 2044 30104
rect 2038 30064 2044 30076
rect 2096 30064 2102 30116
rect 5166 30064 5172 30116
rect 5224 30104 5230 30116
rect 5353 30107 5411 30113
rect 5353 30104 5365 30107
rect 5224 30076 5365 30104
rect 5224 30064 5230 30076
rect 5353 30073 5365 30076
rect 5399 30073 5411 30107
rect 5353 30067 5411 30073
rect 3053 30039 3111 30045
rect 3053 30005 3065 30039
rect 3099 30036 3111 30039
rect 6886 30036 6914 30144
rect 9030 30064 9036 30116
rect 9088 30104 9094 30116
rect 9309 30107 9367 30113
rect 9309 30104 9321 30107
rect 9088 30076 9321 30104
rect 9088 30064 9094 30076
rect 9309 30073 9321 30076
rect 9355 30073 9367 30107
rect 9309 30067 9367 30073
rect 11606 30064 11612 30116
rect 11664 30104 11670 30116
rect 11885 30107 11943 30113
rect 11885 30104 11897 30107
rect 11664 30076 11897 30104
rect 11664 30064 11670 30076
rect 11885 30073 11897 30076
rect 11931 30073 11943 30107
rect 13078 30104 13084 30116
rect 11885 30067 11943 30073
rect 12406 30076 13084 30104
rect 3099 30008 6914 30036
rect 3099 30005 3111 30008
rect 3053 29999 3111 30005
rect 10962 29996 10968 30048
rect 11020 30036 11026 30048
rect 12406 30036 12434 30076
rect 13078 30064 13084 30076
rect 13136 30064 13142 30116
rect 11020 30008 12434 30036
rect 13280 30036 13308 30144
rect 13906 30132 13912 30144
rect 13964 30132 13970 30184
rect 13354 30064 13360 30116
rect 13412 30104 13418 30116
rect 14277 30107 14335 30113
rect 14277 30104 14289 30107
rect 13412 30076 14289 30104
rect 13412 30064 13418 30076
rect 14277 30073 14289 30076
rect 14323 30073 14335 30107
rect 17497 30107 17555 30113
rect 17497 30104 17509 30107
rect 14277 30067 14335 30073
rect 15856 30076 17509 30104
rect 15856 30036 15884 30076
rect 17497 30073 17509 30076
rect 17543 30104 17555 30107
rect 17954 30104 17960 30116
rect 17543 30076 17960 30104
rect 17543 30073 17555 30076
rect 17497 30067 17555 30073
rect 17954 30064 17960 30076
rect 18012 30064 18018 30116
rect 18325 30107 18383 30113
rect 18325 30073 18337 30107
rect 18371 30104 18383 30107
rect 22646 30104 22652 30116
rect 18371 30076 22652 30104
rect 18371 30073 18383 30076
rect 18325 30067 18383 30073
rect 22646 30064 22652 30076
rect 22704 30064 22710 30116
rect 26418 30064 26424 30116
rect 26476 30104 26482 30116
rect 27157 30107 27215 30113
rect 27157 30104 27169 30107
rect 26476 30076 27169 30104
rect 26476 30064 26482 30076
rect 27157 30073 27169 30076
rect 27203 30073 27215 30107
rect 27157 30067 27215 30073
rect 28350 30064 28356 30116
rect 28408 30104 28414 30116
rect 28629 30107 28687 30113
rect 28629 30104 28641 30107
rect 28408 30076 28641 30104
rect 28408 30064 28414 30076
rect 28629 30073 28641 30076
rect 28675 30073 28687 30107
rect 28629 30067 28687 30073
rect 13280 30008 15884 30036
rect 15933 30039 15991 30045
rect 11020 29996 11026 30008
rect 15933 30005 15945 30039
rect 15979 30036 15991 30039
rect 16022 30036 16028 30048
rect 15979 30008 16028 30036
rect 15979 30005 15991 30008
rect 15933 29999 15991 30005
rect 16022 29996 16028 30008
rect 16080 29996 16086 30048
rect 20070 29996 20076 30048
rect 20128 30036 20134 30048
rect 20257 30039 20315 30045
rect 20257 30036 20269 30039
rect 20128 30008 20269 30036
rect 20128 29996 20134 30008
rect 20257 30005 20269 30008
rect 20303 30005 20315 30039
rect 20257 29999 20315 30005
rect 22002 29996 22008 30048
rect 22060 30036 22066 30048
rect 22189 30039 22247 30045
rect 22189 30036 22201 30039
rect 22060 30008 22201 30036
rect 22060 29996 22066 30008
rect 22189 30005 22201 30008
rect 22235 30005 22247 30039
rect 22189 29999 22247 30005
rect 24394 29996 24400 30048
rect 24452 30036 24458 30048
rect 24765 30039 24823 30045
rect 24765 30036 24777 30039
rect 24452 30008 24777 30036
rect 24452 29996 24458 30008
rect 24765 30005 24777 30008
rect 24811 30005 24823 30039
rect 26326 30036 26332 30048
rect 26287 30008 26332 30036
rect 24765 29999 24823 30005
rect 26326 29996 26332 30008
rect 26384 29996 26390 30048
rect 27890 30036 27896 30048
rect 27851 30008 27896 30036
rect 27890 29996 27896 30008
rect 27948 29996 27954 30048
rect 1104 29946 29440 29968
rect 1104 29894 4492 29946
rect 4544 29894 4556 29946
rect 4608 29894 4620 29946
rect 4672 29894 4684 29946
rect 4736 29894 4748 29946
rect 4800 29894 11576 29946
rect 11628 29894 11640 29946
rect 11692 29894 11704 29946
rect 11756 29894 11768 29946
rect 11820 29894 11832 29946
rect 11884 29894 18660 29946
rect 18712 29894 18724 29946
rect 18776 29894 18788 29946
rect 18840 29894 18852 29946
rect 18904 29894 18916 29946
rect 18968 29894 25744 29946
rect 25796 29894 25808 29946
rect 25860 29894 25872 29946
rect 25924 29894 25936 29946
rect 25988 29894 26000 29946
rect 26052 29894 29440 29946
rect 1104 29872 29440 29894
rect 2590 29832 2596 29844
rect 2551 29804 2596 29832
rect 2590 29792 2596 29804
rect 2648 29792 2654 29844
rect 19978 29832 19984 29844
rect 19939 29804 19984 29832
rect 19978 29792 19984 29804
rect 20036 29792 20042 29844
rect 22094 29792 22100 29844
rect 22152 29832 22158 29844
rect 22373 29835 22431 29841
rect 22373 29832 22385 29835
rect 22152 29804 22385 29832
rect 22152 29792 22158 29804
rect 22373 29801 22385 29804
rect 22419 29801 22431 29835
rect 24486 29832 24492 29844
rect 24447 29804 24492 29832
rect 22373 29795 22431 29801
rect 24486 29792 24492 29804
rect 24544 29792 24550 29844
rect 1302 29724 1308 29776
rect 1360 29764 1366 29776
rect 3053 29767 3111 29773
rect 3053 29764 3065 29767
rect 1360 29736 3065 29764
rect 1360 29724 1366 29736
rect 3053 29733 3065 29736
rect 3099 29733 3111 29767
rect 13354 29764 13360 29776
rect 3053 29727 3111 29733
rect 12544 29736 13360 29764
rect 12544 29705 12572 29736
rect 13354 29724 13360 29736
rect 13412 29724 13418 29776
rect 15654 29724 15660 29776
rect 15712 29764 15718 29776
rect 16301 29767 16359 29773
rect 16301 29764 16313 29767
rect 15712 29736 16313 29764
rect 15712 29724 15718 29736
rect 16301 29733 16313 29736
rect 16347 29733 16359 29767
rect 16301 29727 16359 29733
rect 12529 29699 12587 29705
rect 12529 29665 12541 29699
rect 12575 29665 12587 29699
rect 12529 29659 12587 29665
rect 12805 29699 12863 29705
rect 12805 29665 12817 29699
rect 12851 29696 12863 29699
rect 12986 29696 12992 29708
rect 12851 29668 12992 29696
rect 12851 29665 12863 29668
rect 12805 29659 12863 29665
rect 12986 29656 12992 29668
rect 13044 29656 13050 29708
rect 17129 29699 17187 29705
rect 17129 29696 17141 29699
rect 16500 29668 17141 29696
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29628 1731 29631
rect 2130 29628 2136 29640
rect 1719 29600 2136 29628
rect 1719 29597 1731 29600
rect 1673 29591 1731 29597
rect 2130 29588 2136 29600
rect 2188 29588 2194 29640
rect 12437 29631 12495 29637
rect 12437 29597 12449 29631
rect 12483 29628 12495 29631
rect 12894 29628 12900 29640
rect 12483 29600 12900 29628
rect 12483 29597 12495 29600
rect 12437 29591 12495 29597
rect 12894 29588 12900 29600
rect 12952 29588 12958 29640
rect 16500 29637 16528 29668
rect 17129 29665 17141 29668
rect 17175 29696 17187 29699
rect 18230 29696 18236 29708
rect 17175 29668 18236 29696
rect 17175 29665 17187 29668
rect 17129 29659 17187 29665
rect 18230 29656 18236 29668
rect 18288 29656 18294 29708
rect 21361 29699 21419 29705
rect 21361 29665 21373 29699
rect 21407 29696 21419 29699
rect 22097 29699 22155 29705
rect 22097 29696 22109 29699
rect 21407 29668 22109 29696
rect 21407 29665 21419 29668
rect 21361 29659 21419 29665
rect 22097 29665 22109 29668
rect 22143 29696 22155 29699
rect 22830 29696 22836 29708
rect 22143 29668 22836 29696
rect 22143 29665 22155 29668
rect 22097 29659 22155 29665
rect 22830 29656 22836 29668
rect 22888 29656 22894 29708
rect 16485 29631 16543 29637
rect 16485 29597 16497 29631
rect 16531 29597 16543 29631
rect 16485 29591 16543 29597
rect 16577 29631 16635 29637
rect 16577 29597 16589 29631
rect 16623 29628 16635 29631
rect 16850 29628 16856 29640
rect 16623 29600 16856 29628
rect 16623 29597 16635 29600
rect 16577 29591 16635 29597
rect 16850 29588 16856 29600
rect 16908 29588 16914 29640
rect 17862 29628 17868 29640
rect 17823 29600 17868 29628
rect 17862 29588 17868 29600
rect 17920 29588 17926 29640
rect 17954 29588 17960 29640
rect 18012 29628 18018 29640
rect 18509 29631 18567 29637
rect 18509 29628 18521 29631
rect 18012 29600 18521 29628
rect 18012 29588 18018 29600
rect 18509 29597 18521 29600
rect 18555 29628 18567 29631
rect 20162 29628 20168 29640
rect 18555 29600 20168 29628
rect 18555 29597 18567 29600
rect 18509 29591 18567 29597
rect 20162 29588 20168 29600
rect 20220 29588 20226 29640
rect 22005 29631 22063 29637
rect 22005 29597 22017 29631
rect 22051 29628 22063 29631
rect 22646 29628 22652 29640
rect 22051 29600 22652 29628
rect 22051 29597 22063 29600
rect 22005 29591 22063 29597
rect 22646 29588 22652 29600
rect 22704 29588 22710 29640
rect 27065 29631 27123 29637
rect 27065 29597 27077 29631
rect 27111 29628 27123 29631
rect 28721 29631 28779 29637
rect 28721 29628 28733 29631
rect 27111 29600 28733 29628
rect 27111 29597 27123 29600
rect 27065 29591 27123 29597
rect 28721 29597 28733 29600
rect 28767 29628 28779 29631
rect 30282 29628 30288 29640
rect 28767 29600 30288 29628
rect 28767 29597 28779 29600
rect 28721 29591 28779 29597
rect 30282 29588 30288 29600
rect 30340 29588 30346 29640
rect 16301 29563 16359 29569
rect 16301 29529 16313 29563
rect 16347 29560 16359 29563
rect 16347 29532 17264 29560
rect 16347 29529 16359 29532
rect 16301 29523 16359 29529
rect 17236 29504 17264 29532
rect 1486 29492 1492 29504
rect 1447 29464 1492 29492
rect 1486 29452 1492 29464
rect 1544 29452 1550 29504
rect 8754 29452 8760 29504
rect 8812 29492 8818 29504
rect 9217 29495 9275 29501
rect 9217 29492 9229 29495
rect 8812 29464 9229 29492
rect 8812 29452 8818 29464
rect 9217 29461 9229 29464
rect 9263 29492 9275 29495
rect 9398 29492 9404 29504
rect 9263 29464 9404 29492
rect 9263 29461 9275 29464
rect 9217 29455 9275 29461
rect 9398 29452 9404 29464
rect 9456 29452 9462 29504
rect 11330 29452 11336 29504
rect 11388 29492 11394 29504
rect 11517 29495 11575 29501
rect 11517 29492 11529 29495
rect 11388 29464 11529 29492
rect 11388 29452 11394 29464
rect 11517 29461 11529 29464
rect 11563 29461 11575 29495
rect 11517 29455 11575 29461
rect 17218 29452 17224 29504
rect 17276 29492 17282 29504
rect 17681 29495 17739 29501
rect 17681 29492 17693 29495
rect 17276 29464 17693 29492
rect 17276 29452 17282 29464
rect 17681 29461 17693 29464
rect 17727 29461 17739 29495
rect 27614 29492 27620 29504
rect 27575 29464 27620 29492
rect 17681 29455 17739 29461
rect 27614 29452 27620 29464
rect 27672 29452 27678 29504
rect 28537 29495 28595 29501
rect 28537 29461 28549 29495
rect 28583 29492 28595 29495
rect 28810 29492 28816 29504
rect 28583 29464 28816 29492
rect 28583 29461 28595 29464
rect 28537 29455 28595 29461
rect 28810 29452 28816 29464
rect 28868 29452 28874 29504
rect 1104 29402 29600 29424
rect 1104 29350 8034 29402
rect 8086 29350 8098 29402
rect 8150 29350 8162 29402
rect 8214 29350 8226 29402
rect 8278 29350 8290 29402
rect 8342 29350 15118 29402
rect 15170 29350 15182 29402
rect 15234 29350 15246 29402
rect 15298 29350 15310 29402
rect 15362 29350 15374 29402
rect 15426 29350 22202 29402
rect 22254 29350 22266 29402
rect 22318 29350 22330 29402
rect 22382 29350 22394 29402
rect 22446 29350 22458 29402
rect 22510 29350 29286 29402
rect 29338 29350 29350 29402
rect 29402 29350 29414 29402
rect 29466 29350 29478 29402
rect 29530 29350 29542 29402
rect 29594 29350 29600 29402
rect 1104 29328 29600 29350
rect 12986 29288 12992 29300
rect 12947 29260 12992 29288
rect 12986 29248 12992 29260
rect 13044 29248 13050 29300
rect 16850 29248 16856 29300
rect 16908 29288 16914 29300
rect 16908 29260 19012 29288
rect 16908 29248 16914 29260
rect 1854 29220 1860 29232
rect 1815 29192 1860 29220
rect 1854 29180 1860 29192
rect 1912 29180 1918 29232
rect 8662 29220 8668 29232
rect 6886 29192 8668 29220
rect 6730 29152 6736 29164
rect 6691 29124 6736 29152
rect 6730 29112 6736 29124
rect 6788 29112 6794 29164
rect 6886 29152 6914 29192
rect 8662 29180 8668 29192
rect 8720 29180 8726 29232
rect 12894 29220 12900 29232
rect 12855 29192 12900 29220
rect 12894 29180 12900 29192
rect 12952 29180 12958 29232
rect 16574 29220 16580 29232
rect 15580 29192 16580 29220
rect 6840 29124 6914 29152
rect 7745 29155 7803 29161
rect 2130 29044 2136 29096
rect 2188 29084 2194 29096
rect 6840 29093 6868 29124
rect 7745 29121 7757 29155
rect 7791 29152 7803 29155
rect 8294 29152 8300 29164
rect 7791 29124 8300 29152
rect 7791 29121 7803 29124
rect 7745 29115 7803 29121
rect 8294 29112 8300 29124
rect 8352 29112 8358 29164
rect 8754 29152 8760 29164
rect 8715 29124 8760 29152
rect 8754 29112 8760 29124
rect 8812 29112 8818 29164
rect 15580 29161 15608 29192
rect 16574 29180 16580 29192
rect 16632 29220 16638 29232
rect 18984 29229 19012 29260
rect 18969 29223 19027 29229
rect 16632 29192 17172 29220
rect 16632 29180 16638 29192
rect 15565 29155 15623 29161
rect 15565 29121 15577 29155
rect 15611 29121 15623 29155
rect 16850 29152 16856 29164
rect 16811 29124 16856 29152
rect 15565 29115 15623 29121
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 16942 29112 16948 29164
rect 17000 29152 17006 29164
rect 17144 29161 17172 29192
rect 18969 29189 18981 29223
rect 19015 29189 19027 29223
rect 18969 29183 19027 29189
rect 17129 29155 17187 29161
rect 17000 29124 17045 29152
rect 17000 29112 17006 29124
rect 17129 29121 17141 29155
rect 17175 29121 17187 29155
rect 17129 29115 17187 29121
rect 17218 29112 17224 29164
rect 17276 29152 17282 29164
rect 17276 29124 17321 29152
rect 17276 29112 17282 29124
rect 17954 29112 17960 29164
rect 18012 29152 18018 29164
rect 18233 29155 18291 29161
rect 18233 29152 18245 29155
rect 18012 29124 18245 29152
rect 18012 29112 18018 29124
rect 18233 29121 18245 29124
rect 18279 29121 18291 29155
rect 18984 29152 19012 29183
rect 19150 29180 19156 29232
rect 19208 29220 19214 29232
rect 19208 29192 19932 29220
rect 19208 29180 19214 29192
rect 19610 29152 19616 29164
rect 18233 29115 18291 29121
rect 2501 29087 2559 29093
rect 2501 29084 2513 29087
rect 2188 29056 2513 29084
rect 2188 29044 2194 29056
rect 2501 29053 2513 29056
rect 2547 29053 2559 29087
rect 2501 29047 2559 29053
rect 6825 29087 6883 29093
rect 6825 29053 6837 29087
rect 6871 29053 6883 29087
rect 6825 29047 6883 29053
rect 7837 29087 7895 29093
rect 7837 29053 7849 29087
rect 7883 29084 7895 29087
rect 8386 29084 8392 29096
rect 7883 29056 8392 29084
rect 7883 29053 7895 29056
rect 7837 29047 7895 29053
rect 8386 29044 8392 29056
rect 8444 29044 8450 29096
rect 8665 29087 8723 29093
rect 8665 29053 8677 29087
rect 8711 29084 8723 29087
rect 9677 29087 9735 29093
rect 9677 29084 9689 29087
rect 8711 29056 9689 29084
rect 8711 29053 8723 29056
rect 8665 29047 8723 29053
rect 9677 29053 9689 29056
rect 9723 29084 9735 29087
rect 10134 29084 10140 29096
rect 9723 29056 10140 29084
rect 9723 29053 9735 29056
rect 9677 29047 9735 29053
rect 10134 29044 10140 29056
rect 10192 29044 10198 29096
rect 12986 29044 12992 29096
rect 13044 29084 13050 29096
rect 13173 29087 13231 29093
rect 13173 29084 13185 29087
rect 13044 29056 13185 29084
rect 13044 29044 13050 29056
rect 13173 29053 13185 29056
rect 13219 29084 13231 29087
rect 15654 29084 15660 29096
rect 13219 29056 13768 29084
rect 15615 29056 15660 29084
rect 13219 29053 13231 29056
rect 13173 29047 13231 29053
rect 2041 29019 2099 29025
rect 2041 28985 2053 29019
rect 2087 29016 2099 29019
rect 4982 29016 4988 29028
rect 2087 28988 4988 29016
rect 2087 28985 2099 28988
rect 2041 28979 2099 28985
rect 4982 28976 4988 28988
rect 5040 28976 5046 29028
rect 5810 28976 5816 29028
rect 5868 29016 5874 29028
rect 6365 29019 6423 29025
rect 6365 29016 6377 29019
rect 5868 28988 6377 29016
rect 5868 28976 5874 28988
rect 6365 28985 6377 28988
rect 6411 28985 6423 29019
rect 6365 28979 6423 28985
rect 8113 29019 8171 29025
rect 8113 28985 8125 29019
rect 8159 29016 8171 29019
rect 9306 29016 9312 29028
rect 8159 28988 9312 29016
rect 8159 28985 8171 28988
rect 8113 28979 8171 28985
rect 9306 28976 9312 28988
rect 9364 28976 9370 29028
rect 12529 29019 12587 29025
rect 12529 28985 12541 29019
rect 12575 29016 12587 29019
rect 12618 29016 12624 29028
rect 12575 28988 12624 29016
rect 12575 28985 12587 28988
rect 12529 28979 12587 28985
rect 12618 28976 12624 28988
rect 12676 28976 12682 29028
rect 9122 28948 9128 28960
rect 9083 28920 9128 28948
rect 9122 28908 9128 28920
rect 9180 28908 9186 28960
rect 10226 28948 10232 28960
rect 10139 28920 10232 28948
rect 10226 28908 10232 28920
rect 10284 28948 10290 28960
rect 13630 28948 13636 28960
rect 10284 28920 13636 28948
rect 10284 28908 10290 28920
rect 13630 28908 13636 28920
rect 13688 28908 13694 28960
rect 13740 28948 13768 29056
rect 15654 29044 15660 29056
rect 15712 29044 15718 29096
rect 17862 29044 17868 29096
rect 17920 29084 17926 29096
rect 18800 29084 18828 29138
rect 18984 29124 19616 29152
rect 19610 29112 19616 29124
rect 19668 29152 19674 29164
rect 19904 29161 19932 29192
rect 19705 29155 19763 29161
rect 19705 29152 19717 29155
rect 19668 29124 19717 29152
rect 19668 29112 19674 29124
rect 19705 29121 19717 29124
rect 19751 29121 19763 29155
rect 19705 29115 19763 29121
rect 19889 29155 19947 29161
rect 19889 29121 19901 29155
rect 19935 29152 19947 29155
rect 20349 29155 20407 29161
rect 20349 29152 20361 29155
rect 19935 29124 20361 29152
rect 19935 29121 19947 29124
rect 19889 29115 19947 29121
rect 20349 29121 20361 29124
rect 20395 29121 20407 29155
rect 20349 29115 20407 29121
rect 21450 29112 21456 29164
rect 21508 29152 21514 29164
rect 22002 29152 22008 29164
rect 21508 29124 22008 29152
rect 21508 29112 21514 29124
rect 22002 29112 22008 29124
rect 22060 29152 22066 29164
rect 22097 29155 22155 29161
rect 22097 29152 22109 29155
rect 22060 29124 22109 29152
rect 22060 29112 22066 29124
rect 22097 29121 22109 29124
rect 22143 29121 22155 29155
rect 22097 29115 22155 29121
rect 22646 29112 22652 29164
rect 22704 29152 22710 29164
rect 22833 29155 22891 29161
rect 22833 29152 22845 29155
rect 22704 29124 22845 29152
rect 22704 29112 22710 29124
rect 22833 29121 22845 29124
rect 22879 29121 22891 29155
rect 22833 29115 22891 29121
rect 17920 29056 18828 29084
rect 17920 29044 17926 29056
rect 18800 29016 18828 29056
rect 19242 29016 19248 29028
rect 15212 28988 15608 29016
rect 18800 28988 19248 29016
rect 15212 28948 15240 28988
rect 13740 28920 15240 28948
rect 15289 28951 15347 28957
rect 15289 28917 15301 28951
rect 15335 28948 15347 28951
rect 15470 28948 15476 28960
rect 15335 28920 15476 28948
rect 15335 28917 15347 28920
rect 15289 28911 15347 28917
rect 15470 28908 15476 28920
rect 15528 28908 15534 28960
rect 15580 28948 15608 28988
rect 19242 28976 19248 28988
rect 19300 28976 19306 29028
rect 19978 28976 19984 29028
rect 20036 29016 20042 29028
rect 21913 29019 21971 29025
rect 21913 29016 21925 29019
rect 20036 28988 21925 29016
rect 20036 28976 20042 28988
rect 21913 28985 21925 28988
rect 21959 28985 21971 29019
rect 28258 29016 28264 29028
rect 28219 28988 28264 29016
rect 21913 28979 21971 28985
rect 28258 28976 28264 28988
rect 28316 28976 28322 29028
rect 16669 28951 16727 28957
rect 16669 28948 16681 28951
rect 15580 28920 16681 28948
rect 16669 28917 16681 28920
rect 16715 28917 16727 28951
rect 19794 28948 19800 28960
rect 19755 28920 19800 28948
rect 16669 28911 16727 28917
rect 19794 28908 19800 28920
rect 19852 28908 19858 28960
rect 21266 28948 21272 28960
rect 21227 28920 21272 28948
rect 21266 28908 21272 28920
rect 21324 28908 21330 28960
rect 22830 28908 22836 28960
rect 22888 28948 22894 28960
rect 22925 28951 22983 28957
rect 22925 28948 22937 28951
rect 22888 28920 22937 28948
rect 22888 28908 22894 28920
rect 22925 28917 22937 28920
rect 22971 28917 22983 28951
rect 22925 28911 22983 28917
rect 23014 28908 23020 28960
rect 23072 28948 23078 28960
rect 23293 28951 23351 28957
rect 23293 28948 23305 28951
rect 23072 28920 23305 28948
rect 23072 28908 23078 28920
rect 23293 28917 23305 28920
rect 23339 28917 23351 28951
rect 23750 28948 23756 28960
rect 23711 28920 23756 28948
rect 23293 28911 23351 28917
rect 23750 28908 23756 28920
rect 23808 28908 23814 28960
rect 1104 28858 29440 28880
rect 1104 28806 4492 28858
rect 4544 28806 4556 28858
rect 4608 28806 4620 28858
rect 4672 28806 4684 28858
rect 4736 28806 4748 28858
rect 4800 28806 11576 28858
rect 11628 28806 11640 28858
rect 11692 28806 11704 28858
rect 11756 28806 11768 28858
rect 11820 28806 11832 28858
rect 11884 28806 18660 28858
rect 18712 28806 18724 28858
rect 18776 28806 18788 28858
rect 18840 28806 18852 28858
rect 18904 28806 18916 28858
rect 18968 28806 25744 28858
rect 25796 28806 25808 28858
rect 25860 28806 25872 28858
rect 25924 28806 25936 28858
rect 25988 28806 26000 28858
rect 26052 28806 29440 28858
rect 1104 28784 29440 28806
rect 1673 28747 1731 28753
rect 1673 28713 1685 28747
rect 1719 28744 1731 28747
rect 1854 28744 1860 28756
rect 1719 28716 1860 28744
rect 1719 28713 1731 28716
rect 1673 28707 1731 28713
rect 1854 28704 1860 28716
rect 1912 28704 1918 28756
rect 6365 28747 6423 28753
rect 6365 28713 6377 28747
rect 6411 28744 6423 28747
rect 6730 28744 6736 28756
rect 6411 28716 6736 28744
rect 6411 28713 6423 28716
rect 6365 28707 6423 28713
rect 6730 28704 6736 28716
rect 6788 28704 6794 28756
rect 7193 28747 7251 28753
rect 7193 28713 7205 28747
rect 7239 28744 7251 28747
rect 7834 28744 7840 28756
rect 7239 28716 7840 28744
rect 7239 28713 7251 28716
rect 7193 28707 7251 28713
rect 7208 28676 7236 28707
rect 7834 28704 7840 28716
rect 7892 28704 7898 28756
rect 8386 28704 8392 28756
rect 8444 28744 8450 28756
rect 10226 28744 10232 28756
rect 8444 28716 10232 28744
rect 8444 28704 8450 28716
rect 10226 28704 10232 28716
rect 10284 28704 10290 28756
rect 19610 28744 19616 28756
rect 19571 28716 19616 28744
rect 19610 28704 19616 28716
rect 19668 28704 19674 28756
rect 6104 28648 7236 28676
rect 6104 28617 6132 28648
rect 8662 28636 8668 28688
rect 8720 28676 8726 28688
rect 8941 28679 8999 28685
rect 8941 28676 8953 28679
rect 8720 28648 8953 28676
rect 8720 28636 8726 28648
rect 8941 28645 8953 28648
rect 8987 28645 8999 28679
rect 16206 28676 16212 28688
rect 16167 28648 16212 28676
rect 8941 28639 8999 28645
rect 16206 28636 16212 28648
rect 16264 28636 16270 28688
rect 19242 28636 19248 28688
rect 19300 28676 19306 28688
rect 22097 28679 22155 28685
rect 22097 28676 22109 28679
rect 19300 28648 22109 28676
rect 19300 28636 19306 28648
rect 22097 28645 22109 28648
rect 22143 28645 22155 28679
rect 22097 28639 22155 28645
rect 6089 28611 6147 28617
rect 6089 28577 6101 28611
rect 6135 28577 6147 28611
rect 6089 28571 6147 28577
rect 9122 28568 9128 28620
rect 9180 28608 9186 28620
rect 9217 28611 9275 28617
rect 9217 28608 9229 28611
rect 9180 28580 9229 28608
rect 9180 28568 9186 28580
rect 9217 28577 9229 28580
rect 9263 28577 9275 28611
rect 9217 28571 9275 28577
rect 11885 28611 11943 28617
rect 11885 28577 11897 28611
rect 11931 28608 11943 28611
rect 12434 28608 12440 28620
rect 11931 28580 12440 28608
rect 11931 28577 11943 28580
rect 11885 28571 11943 28577
rect 12434 28568 12440 28580
rect 12492 28568 12498 28620
rect 13814 28568 13820 28620
rect 13872 28608 13878 28620
rect 14826 28608 14832 28620
rect 13872 28580 14832 28608
rect 13872 28568 13878 28580
rect 14826 28568 14832 28580
rect 14884 28568 14890 28620
rect 18230 28608 18236 28620
rect 18143 28580 18236 28608
rect 18230 28568 18236 28580
rect 18288 28608 18294 28620
rect 19150 28608 19156 28620
rect 18288 28580 19156 28608
rect 18288 28568 18294 28580
rect 19150 28568 19156 28580
rect 19208 28608 19214 28620
rect 19705 28611 19763 28617
rect 19705 28608 19717 28611
rect 19208 28580 19717 28608
rect 19208 28568 19214 28580
rect 19705 28577 19717 28580
rect 19751 28608 19763 28611
rect 20717 28611 20775 28617
rect 20717 28608 20729 28611
rect 19751 28580 20729 28608
rect 19751 28577 19763 28580
rect 19705 28571 19763 28577
rect 20717 28577 20729 28580
rect 20763 28577 20775 28611
rect 20717 28571 20775 28577
rect 21266 28568 21272 28620
rect 21324 28608 21330 28620
rect 21818 28608 21824 28620
rect 21324 28580 21824 28608
rect 21324 28568 21330 28580
rect 21818 28568 21824 28580
rect 21876 28608 21882 28620
rect 21913 28611 21971 28617
rect 21913 28608 21925 28611
rect 21876 28580 21925 28608
rect 21876 28568 21882 28580
rect 21913 28577 21925 28580
rect 21959 28577 21971 28611
rect 21913 28571 21971 28577
rect 22112 28580 23428 28608
rect 22112 28552 22140 28580
rect 5534 28500 5540 28552
rect 5592 28540 5598 28552
rect 5997 28543 6055 28549
rect 5997 28540 6009 28543
rect 5592 28512 6009 28540
rect 5592 28500 5598 28512
rect 5997 28509 6009 28512
rect 6043 28540 6055 28543
rect 7098 28540 7104 28552
rect 6043 28512 7104 28540
rect 6043 28509 6055 28512
rect 5997 28503 6055 28509
rect 7098 28500 7104 28512
rect 7156 28500 7162 28552
rect 7193 28543 7251 28549
rect 7193 28509 7205 28543
rect 7239 28540 7251 28543
rect 8938 28540 8944 28552
rect 7239 28512 8944 28540
rect 7239 28509 7251 28512
rect 7193 28503 7251 28509
rect 8938 28500 8944 28512
rect 8996 28500 9002 28552
rect 9306 28540 9312 28552
rect 9267 28512 9312 28540
rect 9306 28500 9312 28512
rect 9364 28500 9370 28552
rect 11790 28540 11796 28552
rect 11751 28512 11796 28540
rect 11790 28500 11796 28512
rect 11848 28540 11854 28552
rect 12805 28543 12863 28549
rect 12805 28540 12817 28543
rect 11848 28512 12817 28540
rect 11848 28500 11854 28512
rect 12805 28509 12817 28512
rect 12851 28540 12863 28543
rect 12894 28540 12900 28552
rect 12851 28512 12900 28540
rect 12851 28509 12863 28512
rect 12805 28503 12863 28509
rect 12894 28500 12900 28512
rect 12952 28500 12958 28552
rect 13081 28543 13139 28549
rect 13081 28509 13093 28543
rect 13127 28540 13139 28543
rect 13354 28540 13360 28552
rect 13127 28512 13360 28540
rect 13127 28509 13139 28512
rect 13081 28503 13139 28509
rect 13354 28500 13360 28512
rect 13412 28500 13418 28552
rect 14550 28540 14556 28552
rect 14511 28512 14556 28540
rect 14550 28500 14556 28512
rect 14608 28500 14614 28552
rect 15838 28500 15844 28552
rect 15896 28540 15902 28552
rect 16025 28543 16083 28549
rect 16025 28540 16037 28543
rect 15896 28512 16037 28540
rect 15896 28500 15902 28512
rect 16025 28509 16037 28512
rect 16071 28509 16083 28543
rect 16298 28540 16304 28552
rect 16259 28512 16304 28540
rect 16025 28503 16083 28509
rect 16298 28500 16304 28512
rect 16356 28500 16362 28552
rect 19429 28543 19487 28549
rect 19429 28509 19441 28543
rect 19475 28509 19487 28543
rect 19429 28503 19487 28509
rect 8294 28472 8300 28484
rect 8207 28444 8300 28472
rect 8294 28432 8300 28444
rect 8352 28472 8358 28484
rect 9214 28472 9220 28484
rect 8352 28444 9220 28472
rect 8352 28432 8358 28444
rect 9214 28432 9220 28444
rect 9272 28472 9278 28484
rect 10045 28475 10103 28481
rect 10045 28472 10057 28475
rect 9272 28444 10057 28472
rect 9272 28432 9278 28444
rect 10045 28441 10057 28444
rect 10091 28472 10103 28475
rect 16206 28472 16212 28484
rect 10091 28444 16212 28472
rect 10091 28441 10103 28444
rect 10045 28435 10103 28441
rect 16206 28432 16212 28444
rect 16264 28432 16270 28484
rect 16942 28432 16948 28484
rect 17000 28472 17006 28484
rect 17405 28475 17463 28481
rect 17405 28472 17417 28475
rect 17000 28444 17417 28472
rect 17000 28432 17006 28444
rect 17405 28441 17417 28444
rect 17451 28472 17463 28475
rect 17957 28475 18015 28481
rect 17957 28472 17969 28475
rect 17451 28444 17969 28472
rect 17451 28441 17463 28444
rect 17405 28435 17463 28441
rect 17957 28441 17969 28444
rect 18003 28472 18015 28475
rect 19444 28472 19472 28503
rect 22094 28500 22100 28552
rect 22152 28540 22158 28552
rect 22465 28543 22523 28549
rect 22152 28512 22197 28540
rect 22152 28500 22158 28512
rect 22465 28509 22477 28543
rect 22511 28540 22523 28543
rect 23014 28540 23020 28552
rect 22511 28512 23020 28540
rect 22511 28509 22523 28512
rect 22465 28503 22523 28509
rect 23014 28500 23020 28512
rect 23072 28500 23078 28552
rect 23400 28549 23428 28580
rect 23109 28543 23167 28549
rect 23109 28509 23121 28543
rect 23155 28540 23167 28543
rect 23385 28543 23443 28549
rect 23155 28512 23336 28540
rect 23155 28509 23167 28512
rect 23109 28503 23167 28509
rect 23198 28472 23204 28484
rect 18003 28444 19380 28472
rect 19444 28444 23204 28472
rect 18003 28441 18015 28444
rect 17957 28435 18015 28441
rect 6638 28364 6644 28416
rect 6696 28404 6702 28416
rect 6825 28407 6883 28413
rect 6825 28404 6837 28407
rect 6696 28376 6837 28404
rect 6696 28364 6702 28376
rect 6825 28373 6837 28376
rect 6871 28373 6883 28407
rect 6825 28367 6883 28373
rect 10134 28364 10140 28416
rect 10192 28404 10198 28416
rect 10505 28407 10563 28413
rect 10505 28404 10517 28407
rect 10192 28376 10517 28404
rect 10192 28364 10198 28376
rect 10505 28373 10517 28376
rect 10551 28373 10563 28407
rect 11146 28404 11152 28416
rect 11107 28376 11152 28404
rect 10505 28367 10563 28373
rect 11146 28364 11152 28376
rect 11204 28364 11210 28416
rect 12158 28404 12164 28416
rect 12119 28376 12164 28404
rect 12158 28364 12164 28376
rect 12216 28364 12222 28416
rect 12526 28364 12532 28416
rect 12584 28404 12590 28416
rect 12621 28407 12679 28413
rect 12621 28404 12633 28407
rect 12584 28376 12633 28404
rect 12584 28364 12590 28376
rect 12621 28373 12633 28376
rect 12667 28373 12679 28407
rect 12986 28404 12992 28416
rect 12947 28376 12992 28404
rect 12621 28367 12679 28373
rect 12986 28364 12992 28376
rect 13044 28364 13050 28416
rect 19150 28364 19156 28416
rect 19208 28404 19214 28416
rect 19245 28407 19303 28413
rect 19245 28404 19257 28407
rect 19208 28376 19257 28404
rect 19208 28364 19214 28376
rect 19245 28373 19257 28376
rect 19291 28373 19303 28407
rect 19352 28404 19380 28444
rect 23198 28432 23204 28444
rect 23256 28432 23262 28484
rect 23308 28472 23336 28512
rect 23385 28509 23397 28543
rect 23431 28540 23443 28543
rect 24397 28543 24455 28549
rect 24397 28540 24409 28543
rect 23431 28512 24409 28540
rect 23431 28509 23443 28512
rect 23385 28503 23443 28509
rect 24397 28509 24409 28512
rect 24443 28509 24455 28543
rect 24397 28503 24455 28509
rect 24581 28543 24639 28549
rect 24581 28509 24593 28543
rect 24627 28540 24639 28543
rect 24627 28512 24661 28540
rect 24627 28509 24639 28512
rect 24581 28503 24639 28509
rect 23658 28472 23664 28484
rect 23308 28444 23664 28472
rect 23658 28432 23664 28444
rect 23716 28432 23722 28484
rect 24596 28472 24624 28503
rect 25041 28475 25099 28481
rect 25041 28472 25053 28475
rect 23768 28444 25053 28472
rect 23768 28416 23796 28444
rect 25041 28441 25053 28444
rect 25087 28441 25099 28475
rect 25041 28435 25099 28441
rect 19978 28404 19984 28416
rect 19352 28376 19984 28404
rect 19245 28367 19303 28373
rect 19978 28364 19984 28376
rect 20036 28404 20042 28416
rect 20165 28407 20223 28413
rect 20165 28404 20177 28407
rect 20036 28376 20177 28404
rect 20036 28364 20042 28376
rect 20165 28373 20177 28376
rect 20211 28373 20223 28407
rect 21266 28404 21272 28416
rect 21227 28376 21272 28404
rect 20165 28367 20223 28373
rect 21266 28364 21272 28376
rect 21324 28364 21330 28416
rect 22554 28364 22560 28416
rect 22612 28404 22618 28416
rect 22925 28407 22983 28413
rect 22925 28404 22937 28407
rect 22612 28376 22937 28404
rect 22612 28364 22618 28376
rect 22925 28373 22937 28376
rect 22971 28373 22983 28407
rect 22925 28367 22983 28373
rect 23293 28407 23351 28413
rect 23293 28373 23305 28407
rect 23339 28404 23351 28407
rect 23750 28404 23756 28416
rect 23339 28376 23756 28404
rect 23339 28373 23351 28376
rect 23293 28367 23351 28373
rect 23750 28364 23756 28376
rect 23808 28364 23814 28416
rect 24486 28404 24492 28416
rect 24447 28376 24492 28404
rect 24486 28364 24492 28376
rect 24544 28364 24550 28416
rect 1104 28314 29600 28336
rect 1104 28262 8034 28314
rect 8086 28262 8098 28314
rect 8150 28262 8162 28314
rect 8214 28262 8226 28314
rect 8278 28262 8290 28314
rect 8342 28262 15118 28314
rect 15170 28262 15182 28314
rect 15234 28262 15246 28314
rect 15298 28262 15310 28314
rect 15362 28262 15374 28314
rect 15426 28262 22202 28314
rect 22254 28262 22266 28314
rect 22318 28262 22330 28314
rect 22382 28262 22394 28314
rect 22446 28262 22458 28314
rect 22510 28262 29286 28314
rect 29338 28262 29350 28314
rect 29402 28262 29414 28314
rect 29466 28262 29478 28314
rect 29530 28262 29542 28314
rect 29594 28262 29600 28314
rect 1104 28240 29600 28262
rect 7834 28200 7840 28212
rect 7795 28172 7840 28200
rect 7834 28160 7840 28172
rect 7892 28160 7898 28212
rect 8938 28200 8944 28212
rect 8899 28172 8944 28200
rect 8938 28160 8944 28172
rect 8996 28160 9002 28212
rect 10137 28203 10195 28209
rect 10137 28169 10149 28203
rect 10183 28200 10195 28203
rect 10226 28200 10232 28212
rect 10183 28172 10232 28200
rect 10183 28169 10195 28172
rect 10137 28163 10195 28169
rect 9401 28135 9459 28141
rect 9401 28101 9413 28135
rect 9447 28132 9459 28135
rect 10152 28132 10180 28163
rect 10226 28160 10232 28172
rect 10284 28160 10290 28212
rect 15470 28160 15476 28212
rect 15528 28160 15534 28212
rect 15838 28200 15844 28212
rect 15799 28172 15844 28200
rect 15838 28160 15844 28172
rect 15896 28160 15902 28212
rect 19061 28203 19119 28209
rect 19061 28169 19073 28203
rect 19107 28200 19119 28203
rect 19794 28200 19800 28212
rect 19107 28172 19800 28200
rect 19107 28169 19119 28172
rect 19061 28163 19119 28169
rect 19794 28160 19800 28172
rect 19852 28160 19858 28212
rect 20714 28160 20720 28212
rect 20772 28200 20778 28212
rect 21913 28203 21971 28209
rect 21913 28200 21925 28203
rect 20772 28172 21925 28200
rect 20772 28160 20778 28172
rect 21913 28169 21925 28172
rect 21959 28169 21971 28203
rect 21913 28163 21971 28169
rect 22097 28203 22155 28209
rect 22097 28169 22109 28203
rect 22143 28200 22155 28203
rect 22143 28172 22779 28200
rect 22143 28169 22155 28172
rect 22097 28163 22155 28169
rect 9447 28104 10180 28132
rect 9447 28101 9459 28104
rect 9401 28095 9459 28101
rect 12158 28092 12164 28144
rect 12216 28132 12222 28144
rect 12216 28104 13308 28132
rect 12216 28092 12222 28104
rect 7650 28064 7656 28076
rect 7611 28036 7656 28064
rect 7650 28024 7656 28036
rect 7708 28024 7714 28076
rect 9125 28067 9183 28073
rect 9125 28033 9137 28067
rect 9171 28064 9183 28067
rect 9306 28064 9312 28076
rect 9171 28036 9312 28064
rect 9171 28033 9183 28036
rect 9125 28027 9183 28033
rect 9306 28024 9312 28036
rect 9364 28024 9370 28076
rect 11790 28024 11796 28076
rect 11848 28064 11854 28076
rect 11885 28067 11943 28073
rect 11885 28064 11897 28067
rect 11848 28036 11897 28064
rect 11848 28024 11854 28036
rect 11885 28033 11897 28036
rect 11931 28033 11943 28067
rect 12894 28064 12900 28076
rect 12855 28036 12900 28064
rect 11885 28027 11943 28033
rect 12894 28024 12900 28036
rect 12952 28024 12958 28076
rect 12986 28024 12992 28076
rect 13044 28064 13050 28076
rect 13280 28073 13308 28104
rect 14826 28092 14832 28144
rect 14884 28132 14890 28144
rect 14884 28104 15332 28132
rect 14884 28092 14890 28104
rect 13173 28067 13231 28073
rect 13044 28036 13089 28064
rect 13044 28024 13050 28036
rect 13173 28033 13185 28067
rect 13219 28033 13231 28067
rect 13173 28027 13231 28033
rect 13265 28067 13323 28073
rect 13265 28033 13277 28067
rect 13311 28033 13323 28067
rect 13265 28027 13323 28033
rect 9214 27996 9220 28008
rect 9175 27968 9220 27996
rect 9214 27956 9220 27968
rect 9272 27956 9278 28008
rect 10686 27956 10692 28008
rect 10744 27996 10750 28008
rect 11609 27999 11667 28005
rect 11609 27996 11621 27999
rect 10744 27968 11621 27996
rect 10744 27956 10750 27968
rect 11609 27965 11621 27968
rect 11655 27965 11667 27999
rect 11609 27959 11667 27965
rect 13188 27996 13216 28027
rect 13722 28024 13728 28076
rect 13780 28064 13786 28076
rect 14461 28067 14519 28073
rect 14461 28064 14473 28067
rect 13780 28036 14473 28064
rect 13780 28024 13786 28036
rect 14461 28033 14473 28036
rect 14507 28033 14519 28067
rect 14461 28027 14519 28033
rect 14476 27996 14504 28027
rect 14918 28024 14924 28076
rect 14976 28064 14982 28076
rect 15197 28067 15255 28073
rect 15197 28064 15209 28067
rect 14976 28036 15209 28064
rect 14976 28024 14982 28036
rect 15197 28033 15209 28036
rect 15243 28033 15255 28067
rect 15304 28070 15332 28104
rect 15360 28073 15418 28079
rect 15488 28076 15516 28160
rect 19981 28135 20039 28141
rect 19981 28101 19993 28135
rect 20027 28132 20039 28135
rect 21358 28132 21364 28144
rect 20027 28104 21364 28132
rect 20027 28101 20039 28104
rect 19981 28095 20039 28101
rect 21358 28092 21364 28104
rect 21416 28092 21422 28144
rect 21542 28092 21548 28144
rect 21600 28132 21606 28144
rect 22112 28132 22140 28163
rect 22646 28132 22652 28144
rect 21600 28104 22140 28132
rect 22388 28104 22652 28132
rect 21600 28092 21606 28104
rect 15360 28070 15372 28073
rect 15304 28042 15372 28070
rect 15360 28039 15372 28042
rect 15406 28039 15418 28073
rect 15360 28033 15418 28039
rect 15460 28070 15518 28076
rect 15460 28036 15472 28070
rect 15506 28036 15518 28070
rect 15197 28027 15255 28033
rect 15460 28030 15518 28036
rect 15565 28067 15623 28073
rect 15565 28033 15577 28067
rect 15611 28033 15623 28067
rect 15565 28027 15623 28033
rect 18877 28067 18935 28073
rect 18877 28033 18889 28067
rect 18923 28033 18935 28067
rect 18877 28027 18935 28033
rect 15579 27996 15607 28027
rect 16666 27996 16672 28008
rect 13188 27968 14044 27996
rect 14476 27968 16672 27996
rect 7742 27888 7748 27940
rect 7800 27928 7806 27940
rect 13188 27928 13216 27968
rect 14016 27937 14044 27968
rect 16666 27956 16672 27968
rect 16724 27956 16730 28008
rect 18892 27996 18920 28027
rect 19150 28024 19156 28076
rect 19208 28064 19214 28076
rect 20162 28064 20168 28076
rect 19208 28036 19253 28064
rect 20123 28036 20168 28064
rect 19208 28024 19214 28036
rect 20162 28024 20168 28036
rect 20220 28064 20226 28076
rect 21177 28067 21235 28073
rect 21177 28064 21189 28067
rect 20220 28036 21189 28064
rect 20220 28024 20226 28036
rect 21177 28033 21189 28036
rect 21223 28064 21235 28067
rect 21266 28064 21272 28076
rect 21223 28036 21272 28064
rect 21223 28033 21235 28036
rect 21177 28027 21235 28033
rect 21266 28024 21272 28036
rect 21324 28024 21330 28076
rect 22094 28024 22100 28076
rect 22152 28064 22158 28076
rect 22388 28064 22416 28104
rect 22646 28092 22652 28104
rect 22704 28092 22710 28144
rect 22751 28132 22779 28172
rect 23198 28160 23204 28212
rect 23256 28200 23262 28212
rect 24213 28203 24271 28209
rect 24213 28200 24225 28203
rect 23256 28172 24225 28200
rect 23256 28160 23262 28172
rect 24213 28169 24225 28172
rect 24259 28169 24271 28203
rect 24213 28163 24271 28169
rect 24381 28203 24439 28209
rect 24381 28169 24393 28203
rect 24427 28200 24439 28203
rect 24670 28200 24676 28212
rect 24427 28172 24676 28200
rect 24427 28169 24439 28172
rect 24381 28163 24439 28169
rect 24670 28160 24676 28172
rect 24728 28160 24734 28212
rect 23106 28132 23112 28144
rect 22751 28104 23112 28132
rect 23106 28092 23112 28104
rect 23164 28132 23170 28144
rect 24578 28132 24584 28144
rect 23164 28104 23796 28132
rect 24539 28104 24584 28132
rect 23164 28092 23170 28104
rect 22554 28064 22560 28076
rect 22152 28036 22416 28064
rect 22515 28036 22560 28064
rect 22152 28024 22158 28036
rect 22554 28024 22560 28036
rect 22612 28024 22618 28076
rect 23385 28067 23443 28073
rect 23385 28033 23397 28067
rect 23431 28064 23443 28067
rect 23474 28064 23480 28076
rect 23431 28036 23480 28064
rect 23431 28033 23443 28036
rect 23385 28027 23443 28033
rect 23474 28024 23480 28036
rect 23532 28024 23538 28076
rect 23569 28067 23627 28073
rect 23569 28033 23581 28067
rect 23615 28064 23627 28067
rect 23658 28064 23664 28076
rect 23615 28036 23664 28064
rect 23615 28033 23627 28036
rect 23569 28027 23627 28033
rect 23658 28024 23664 28036
rect 23716 28024 23722 28076
rect 23768 28064 23796 28104
rect 24578 28092 24584 28104
rect 24636 28092 24642 28144
rect 25041 28067 25099 28073
rect 25041 28064 25053 28067
rect 23768 28036 25053 28064
rect 25041 28033 25053 28036
rect 25087 28033 25099 28067
rect 25041 28027 25099 28033
rect 27985 28067 28043 28073
rect 27985 28033 27997 28067
rect 28031 28064 28043 28067
rect 28626 28064 28632 28076
rect 28031 28036 28632 28064
rect 28031 28033 28043 28036
rect 27985 28027 28043 28033
rect 28626 28024 28632 28036
rect 28684 28024 28690 28076
rect 19610 27996 19616 28008
rect 18892 27968 19616 27996
rect 19610 27956 19616 27968
rect 19668 27956 19674 28008
rect 22465 27999 22523 28005
rect 22465 27965 22477 27999
rect 22511 27996 22523 27999
rect 24486 27996 24492 28008
rect 22511 27968 24492 27996
rect 22511 27965 22523 27968
rect 22465 27959 22523 27965
rect 24486 27956 24492 27968
rect 24544 27956 24550 28008
rect 7800 27900 13216 27928
rect 14001 27931 14059 27937
rect 7800 27888 7806 27900
rect 14001 27897 14013 27931
rect 14047 27928 14059 27931
rect 21726 27928 21732 27940
rect 14047 27900 21732 27928
rect 14047 27897 14059 27900
rect 14001 27891 14059 27897
rect 21726 27888 21732 27900
rect 21784 27888 21790 27940
rect 23934 27928 23940 27940
rect 21836 27900 23940 27928
rect 9401 27863 9459 27869
rect 9401 27829 9413 27863
rect 9447 27860 9459 27863
rect 10134 27860 10140 27872
rect 9447 27832 10140 27860
rect 9447 27829 9459 27832
rect 9401 27823 9459 27829
rect 10134 27820 10140 27832
rect 10192 27820 10198 27872
rect 10965 27863 11023 27869
rect 10965 27829 10977 27863
rect 11011 27860 11023 27863
rect 11054 27860 11060 27872
rect 11011 27832 11060 27860
rect 11011 27829 11023 27832
rect 10965 27823 11023 27829
rect 11054 27820 11060 27832
rect 11112 27820 11118 27872
rect 13449 27863 13507 27869
rect 13449 27829 13461 27863
rect 13495 27860 13507 27863
rect 13814 27860 13820 27872
rect 13495 27832 13820 27860
rect 13495 27829 13507 27832
rect 13449 27823 13507 27829
rect 13814 27820 13820 27832
rect 13872 27820 13878 27872
rect 18506 27820 18512 27872
rect 18564 27860 18570 27872
rect 18877 27863 18935 27869
rect 18877 27860 18889 27863
rect 18564 27832 18889 27860
rect 18564 27820 18570 27832
rect 18877 27829 18889 27832
rect 18923 27829 18935 27863
rect 18877 27823 18935 27829
rect 19797 27863 19855 27869
rect 19797 27829 19809 27863
rect 19843 27860 19855 27863
rect 19886 27860 19892 27872
rect 19843 27832 19892 27860
rect 19843 27829 19855 27832
rect 19797 27823 19855 27829
rect 19886 27820 19892 27832
rect 19944 27820 19950 27872
rect 20162 27820 20168 27872
rect 20220 27860 20226 27872
rect 20717 27863 20775 27869
rect 20717 27860 20729 27863
rect 20220 27832 20729 27860
rect 20220 27820 20226 27832
rect 20717 27829 20729 27832
rect 20763 27860 20775 27863
rect 21836 27860 21864 27900
rect 23934 27888 23940 27900
rect 23992 27888 23998 27940
rect 26142 27888 26148 27940
rect 26200 27928 26206 27940
rect 28445 27931 28503 27937
rect 28445 27928 28457 27931
rect 26200 27900 28457 27928
rect 26200 27888 26206 27900
rect 28445 27897 28457 27900
rect 28491 27897 28503 27931
rect 28445 27891 28503 27897
rect 20763 27832 21864 27860
rect 20763 27829 20775 27832
rect 20717 27823 20775 27829
rect 22738 27820 22744 27872
rect 22796 27860 22802 27872
rect 23201 27863 23259 27869
rect 23201 27860 23213 27863
rect 22796 27832 23213 27860
rect 22796 27820 22802 27832
rect 23201 27829 23213 27832
rect 23247 27829 23259 27863
rect 23201 27823 23259 27829
rect 23474 27820 23480 27872
rect 23532 27860 23538 27872
rect 24302 27860 24308 27872
rect 23532 27832 24308 27860
rect 23532 27820 23538 27832
rect 24302 27820 24308 27832
rect 24360 27860 24366 27872
rect 24397 27863 24455 27869
rect 24397 27860 24409 27863
rect 24360 27832 24409 27860
rect 24360 27820 24366 27832
rect 24397 27829 24409 27832
rect 24443 27829 24455 27863
rect 24397 27823 24455 27829
rect 1104 27770 29440 27792
rect 1104 27718 4492 27770
rect 4544 27718 4556 27770
rect 4608 27718 4620 27770
rect 4672 27718 4684 27770
rect 4736 27718 4748 27770
rect 4800 27718 11576 27770
rect 11628 27718 11640 27770
rect 11692 27718 11704 27770
rect 11756 27718 11768 27770
rect 11820 27718 11832 27770
rect 11884 27718 18660 27770
rect 18712 27718 18724 27770
rect 18776 27718 18788 27770
rect 18840 27718 18852 27770
rect 18904 27718 18916 27770
rect 18968 27718 25744 27770
rect 25796 27718 25808 27770
rect 25860 27718 25872 27770
rect 25924 27718 25936 27770
rect 25988 27718 26000 27770
rect 26052 27718 29440 27770
rect 1104 27696 29440 27718
rect 12621 27659 12679 27665
rect 12621 27625 12633 27659
rect 12667 27656 12679 27659
rect 12894 27656 12900 27668
rect 12667 27628 12900 27656
rect 12667 27625 12679 27628
rect 12621 27619 12679 27625
rect 12894 27616 12900 27628
rect 12952 27616 12958 27668
rect 14461 27659 14519 27665
rect 14461 27625 14473 27659
rect 14507 27656 14519 27659
rect 14550 27656 14556 27668
rect 14507 27628 14556 27656
rect 14507 27625 14519 27628
rect 14461 27619 14519 27625
rect 14550 27616 14556 27628
rect 14608 27616 14614 27668
rect 14642 27616 14648 27668
rect 14700 27656 14706 27668
rect 19610 27656 19616 27668
rect 14700 27628 14745 27656
rect 19571 27628 19616 27656
rect 14700 27616 14706 27628
rect 19610 27616 19616 27628
rect 19668 27616 19674 27668
rect 20993 27659 21051 27665
rect 20993 27625 21005 27659
rect 21039 27656 21051 27659
rect 25498 27656 25504 27668
rect 21039 27628 22094 27656
rect 25459 27628 25504 27656
rect 21039 27625 21051 27628
rect 20993 27619 21051 27625
rect 10686 27588 10692 27600
rect 10647 27560 10692 27588
rect 10686 27548 10692 27560
rect 10744 27548 10750 27600
rect 15654 27548 15660 27600
rect 15712 27588 15718 27600
rect 16853 27591 16911 27597
rect 16853 27588 16865 27591
rect 15712 27560 16865 27588
rect 15712 27548 15718 27560
rect 16853 27557 16865 27560
rect 16899 27588 16911 27591
rect 19702 27588 19708 27600
rect 16899 27560 19708 27588
rect 16899 27557 16911 27560
rect 16853 27551 16911 27557
rect 19702 27548 19708 27560
rect 19760 27588 19766 27600
rect 21542 27588 21548 27600
rect 19760 27560 21548 27588
rect 19760 27548 19766 27560
rect 21542 27548 21548 27560
rect 21600 27548 21606 27600
rect 21726 27588 21732 27600
rect 21687 27560 21732 27588
rect 21726 27548 21732 27560
rect 21784 27548 21790 27600
rect 10042 27480 10048 27532
rect 10100 27520 10106 27532
rect 13722 27520 13728 27532
rect 10100 27492 13728 27520
rect 10100 27480 10106 27492
rect 10413 27455 10471 27461
rect 10413 27421 10425 27455
rect 10459 27421 10471 27455
rect 10413 27415 10471 27421
rect 10505 27455 10563 27461
rect 10505 27421 10517 27455
rect 10551 27452 10563 27455
rect 11149 27455 11207 27461
rect 11149 27452 11161 27455
rect 10551 27424 11161 27452
rect 10551 27421 10563 27424
rect 10505 27415 10563 27421
rect 11149 27421 11161 27424
rect 11195 27452 11207 27455
rect 11238 27452 11244 27464
rect 11195 27424 11244 27452
rect 11195 27421 11207 27424
rect 11149 27415 11207 27421
rect 10428 27384 10456 27415
rect 11238 27412 11244 27424
rect 11296 27412 11302 27464
rect 12452 27461 12480 27492
rect 13722 27480 13728 27492
rect 13780 27480 13786 27532
rect 19242 27480 19248 27532
rect 19300 27520 19306 27532
rect 20625 27523 20683 27529
rect 20625 27520 20637 27523
rect 19300 27492 20637 27520
rect 19300 27480 19306 27492
rect 20625 27489 20637 27492
rect 20671 27489 20683 27523
rect 22066 27520 22094 27628
rect 25498 27616 25504 27628
rect 25556 27616 25562 27668
rect 23753 27523 23811 27529
rect 23753 27520 23765 27523
rect 20625 27483 20683 27489
rect 22020 27492 23765 27520
rect 12437 27455 12495 27461
rect 12437 27421 12449 27455
rect 12483 27421 12495 27455
rect 12618 27452 12624 27464
rect 12579 27424 12624 27452
rect 12437 27415 12495 27421
rect 12618 27412 12624 27424
rect 12676 27412 12682 27464
rect 13814 27412 13820 27464
rect 13872 27452 13878 27464
rect 14645 27455 14703 27461
rect 14645 27452 14657 27455
rect 13872 27424 14657 27452
rect 13872 27412 13878 27424
rect 14645 27421 14657 27424
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 15013 27455 15071 27461
rect 15013 27421 15025 27455
rect 15059 27452 15071 27455
rect 16114 27452 16120 27464
rect 15059 27424 16120 27452
rect 15059 27421 15071 27424
rect 15013 27415 15071 27421
rect 16114 27412 16120 27424
rect 16172 27412 16178 27464
rect 19794 27452 19800 27464
rect 19755 27424 19800 27452
rect 19794 27412 19800 27424
rect 19852 27412 19858 27464
rect 19886 27412 19892 27464
rect 19944 27452 19950 27464
rect 20073 27455 20131 27461
rect 19944 27424 19989 27452
rect 19944 27412 19950 27424
rect 20073 27421 20085 27455
rect 20119 27421 20131 27455
rect 20073 27415 20131 27421
rect 20165 27455 20223 27461
rect 20165 27421 20177 27455
rect 20211 27452 20223 27455
rect 20438 27452 20444 27464
rect 20211 27424 20444 27452
rect 20211 27421 20223 27424
rect 20165 27415 20223 27421
rect 10870 27384 10876 27396
rect 10428 27356 10876 27384
rect 10870 27344 10876 27356
rect 10928 27344 10934 27396
rect 11054 27344 11060 27396
rect 11112 27384 11118 27396
rect 11333 27387 11391 27393
rect 11333 27384 11345 27387
rect 11112 27356 11345 27384
rect 11112 27344 11118 27356
rect 11333 27353 11345 27356
rect 11379 27353 11391 27387
rect 11333 27347 11391 27353
rect 11517 27387 11575 27393
rect 11517 27353 11529 27387
rect 11563 27384 11575 27387
rect 12066 27384 12072 27396
rect 11563 27356 12072 27384
rect 11563 27353 11575 27356
rect 11517 27347 11575 27353
rect 12066 27344 12072 27356
rect 12124 27384 12130 27396
rect 13081 27387 13139 27393
rect 13081 27384 13093 27387
rect 12124 27356 13093 27384
rect 12124 27344 12130 27356
rect 13081 27353 13093 27356
rect 13127 27353 13139 27387
rect 20088 27384 20116 27415
rect 20438 27412 20444 27424
rect 20496 27412 20502 27464
rect 22020 27461 22048 27492
rect 23753 27489 23765 27492
rect 23799 27489 23811 27523
rect 23753 27483 23811 27489
rect 24670 27480 24676 27532
rect 24728 27520 24734 27532
rect 24728 27492 25636 27520
rect 24728 27480 24734 27492
rect 25608 27464 25636 27492
rect 22005 27455 22063 27461
rect 22005 27421 22017 27455
rect 22051 27421 22063 27455
rect 23198 27452 23204 27464
rect 23159 27424 23204 27452
rect 22005 27415 22063 27421
rect 23198 27412 23204 27424
rect 23256 27412 23262 27464
rect 23658 27452 23664 27464
rect 23619 27424 23664 27452
rect 23658 27412 23664 27424
rect 23716 27412 23722 27464
rect 23845 27455 23903 27461
rect 23845 27421 23857 27455
rect 23891 27452 23903 27455
rect 24302 27452 24308 27464
rect 23891 27424 24308 27452
rect 23891 27421 23903 27424
rect 23845 27415 23903 27421
rect 24302 27412 24308 27424
rect 24360 27412 24366 27464
rect 24578 27452 24584 27464
rect 24539 27424 24584 27452
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 25130 27452 25136 27464
rect 25091 27424 25136 27452
rect 25130 27412 25136 27424
rect 25188 27412 25194 27464
rect 25590 27452 25596 27464
rect 25551 27424 25596 27452
rect 25590 27412 25596 27424
rect 25648 27412 25654 27464
rect 20088 27356 21220 27384
rect 13081 27347 13139 27353
rect 8021 27319 8079 27325
rect 8021 27285 8033 27319
rect 8067 27316 8079 27319
rect 8386 27316 8392 27328
rect 8067 27288 8392 27316
rect 8067 27285 8079 27288
rect 8021 27279 8079 27285
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 9309 27319 9367 27325
rect 9309 27285 9321 27319
rect 9355 27316 9367 27319
rect 9398 27316 9404 27328
rect 9355 27288 9404 27316
rect 9355 27285 9367 27288
rect 9309 27279 9367 27285
rect 9398 27276 9404 27288
rect 9456 27276 9462 27328
rect 9861 27319 9919 27325
rect 9861 27285 9873 27319
rect 9907 27316 9919 27319
rect 11146 27316 11152 27328
rect 9907 27288 11152 27316
rect 9907 27285 9919 27288
rect 9861 27279 9919 27285
rect 11146 27276 11152 27288
rect 11204 27276 11210 27328
rect 15749 27319 15807 27325
rect 15749 27285 15761 27319
rect 15795 27316 15807 27319
rect 15838 27316 15844 27328
rect 15795 27288 15844 27316
rect 15795 27285 15807 27288
rect 15749 27279 15807 27285
rect 15838 27276 15844 27288
rect 15896 27276 15902 27328
rect 16206 27316 16212 27328
rect 16167 27288 16212 27316
rect 16206 27276 16212 27288
rect 16264 27276 16270 27328
rect 19610 27276 19616 27328
rect 19668 27316 19674 27328
rect 20162 27316 20168 27328
rect 19668 27288 20168 27316
rect 19668 27276 19674 27288
rect 20162 27276 20168 27288
rect 20220 27276 20226 27328
rect 20990 27316 20996 27328
rect 20951 27288 20996 27316
rect 20990 27276 20996 27288
rect 21048 27276 21054 27328
rect 21192 27325 21220 27356
rect 22646 27344 22652 27396
rect 22704 27384 22710 27396
rect 22925 27387 22983 27393
rect 22925 27384 22937 27387
rect 22704 27356 22937 27384
rect 22704 27344 22710 27356
rect 22925 27353 22937 27356
rect 22971 27353 22983 27387
rect 22925 27347 22983 27353
rect 21177 27319 21235 27325
rect 21177 27285 21189 27319
rect 21223 27285 21235 27319
rect 21177 27279 21235 27285
rect 1104 27226 29600 27248
rect 1104 27174 8034 27226
rect 8086 27174 8098 27226
rect 8150 27174 8162 27226
rect 8214 27174 8226 27226
rect 8278 27174 8290 27226
rect 8342 27174 15118 27226
rect 15170 27174 15182 27226
rect 15234 27174 15246 27226
rect 15298 27174 15310 27226
rect 15362 27174 15374 27226
rect 15426 27174 22202 27226
rect 22254 27174 22266 27226
rect 22318 27174 22330 27226
rect 22382 27174 22394 27226
rect 22446 27174 22458 27226
rect 22510 27174 29286 27226
rect 29338 27174 29350 27226
rect 29402 27174 29414 27226
rect 29466 27174 29478 27226
rect 29530 27174 29542 27226
rect 29594 27174 29600 27226
rect 1104 27152 29600 27174
rect 7377 27115 7435 27121
rect 7377 27081 7389 27115
rect 7423 27112 7435 27115
rect 7650 27112 7656 27124
rect 7423 27084 7656 27112
rect 7423 27081 7435 27084
rect 7377 27075 7435 27081
rect 7650 27072 7656 27084
rect 7708 27072 7714 27124
rect 11146 27112 11152 27124
rect 10980 27084 11152 27112
rect 1578 26936 1584 26988
rect 1636 26976 1642 26988
rect 1857 26979 1915 26985
rect 1857 26976 1869 26979
rect 1636 26948 1869 26976
rect 1636 26936 1642 26948
rect 1857 26945 1869 26948
rect 1903 26945 1915 26979
rect 1857 26939 1915 26945
rect 5534 26936 5540 26988
rect 5592 26976 5598 26988
rect 7561 26979 7619 26985
rect 7561 26976 7573 26979
rect 5592 26948 7573 26976
rect 5592 26936 5598 26948
rect 7561 26945 7573 26948
rect 7607 26945 7619 26979
rect 7561 26939 7619 26945
rect 7837 26979 7895 26985
rect 7837 26945 7849 26979
rect 7883 26976 7895 26979
rect 8938 26976 8944 26988
rect 7883 26948 8944 26976
rect 7883 26945 7895 26948
rect 7837 26939 7895 26945
rect 8938 26936 8944 26948
rect 8996 26936 9002 26988
rect 9769 26979 9827 26985
rect 9769 26945 9781 26979
rect 9815 26976 9827 26979
rect 10226 26976 10232 26988
rect 9815 26948 10232 26976
rect 9815 26945 9827 26948
rect 9769 26939 9827 26945
rect 10226 26936 10232 26948
rect 10284 26976 10290 26988
rect 10980 26985 11008 27084
rect 11146 27072 11152 27084
rect 11204 27112 11210 27124
rect 12069 27115 12127 27121
rect 11204 27084 11836 27112
rect 11204 27072 11210 27084
rect 11238 27004 11244 27056
rect 11296 27044 11302 27056
rect 11808 27053 11836 27084
rect 12069 27081 12081 27115
rect 12115 27112 12127 27115
rect 12986 27112 12992 27124
rect 12115 27084 12992 27112
rect 12115 27081 12127 27084
rect 12069 27075 12127 27081
rect 12986 27072 12992 27084
rect 13044 27072 13050 27124
rect 15654 27112 15660 27124
rect 14292 27084 15660 27112
rect 11701 27047 11759 27053
rect 11701 27044 11713 27047
rect 11296 27016 11713 27044
rect 11296 27004 11302 27016
rect 11701 27013 11713 27016
rect 11747 27013 11759 27047
rect 11701 27007 11759 27013
rect 11793 27047 11851 27053
rect 11793 27013 11805 27047
rect 11839 27044 11851 27047
rect 11974 27044 11980 27056
rect 11839 27016 11980 27044
rect 11839 27013 11851 27016
rect 11793 27007 11851 27013
rect 11974 27004 11980 27016
rect 12032 27004 12038 27056
rect 12434 27004 12440 27056
rect 12492 27044 12498 27056
rect 12621 27047 12679 27053
rect 12621 27044 12633 27047
rect 12492 27016 12633 27044
rect 12492 27004 12498 27016
rect 12621 27013 12633 27016
rect 12667 27013 12679 27047
rect 12621 27007 12679 27013
rect 10781 26979 10839 26985
rect 10781 26976 10793 26979
rect 10284 26948 10793 26976
rect 10284 26936 10290 26948
rect 10781 26945 10793 26948
rect 10827 26945 10839 26979
rect 10781 26939 10839 26945
rect 10965 26979 11023 26985
rect 10965 26945 10977 26979
rect 11011 26945 11023 26979
rect 10965 26939 11023 26945
rect 11517 26979 11575 26985
rect 11517 26945 11529 26979
rect 11563 26945 11575 26979
rect 11517 26939 11575 26945
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26976 11943 26979
rect 11931 26948 12296 26976
rect 11931 26945 11943 26948
rect 11885 26939 11943 26945
rect 7190 26868 7196 26920
rect 7248 26908 7254 26920
rect 7653 26911 7711 26917
rect 7653 26908 7665 26911
rect 7248 26880 7665 26908
rect 7248 26868 7254 26880
rect 7653 26877 7665 26880
rect 7699 26877 7711 26911
rect 10796 26908 10824 26939
rect 11054 26908 11060 26920
rect 10796 26880 11060 26908
rect 7653 26871 7711 26877
rect 11054 26868 11060 26880
rect 11112 26868 11118 26920
rect 11532 26908 11560 26939
rect 11974 26908 11980 26920
rect 11532 26880 11980 26908
rect 11974 26868 11980 26880
rect 12032 26868 12038 26920
rect 12268 26908 12296 26948
rect 12342 26936 12348 26988
rect 12400 26976 12406 26988
rect 12529 26979 12587 26985
rect 12529 26976 12541 26979
rect 12400 26948 12541 26976
rect 12400 26936 12406 26948
rect 12529 26945 12541 26948
rect 12575 26945 12587 26979
rect 12710 26976 12716 26988
rect 12671 26948 12716 26976
rect 12529 26939 12587 26945
rect 12710 26936 12716 26948
rect 12768 26936 12774 26988
rect 14292 26908 14320 27084
rect 15654 27072 15660 27084
rect 15712 27072 15718 27124
rect 15838 27072 15844 27124
rect 15896 27112 15902 27124
rect 19610 27112 19616 27124
rect 15896 27084 19616 27112
rect 15896 27072 15902 27084
rect 19610 27072 19616 27084
rect 19668 27112 19674 27124
rect 20438 27112 20444 27124
rect 19668 27084 20116 27112
rect 20399 27084 20444 27112
rect 19668 27072 19674 27084
rect 14366 27004 14372 27056
rect 14424 27044 14430 27056
rect 14737 27047 14795 27053
rect 14737 27044 14749 27047
rect 14424 27016 14749 27044
rect 14424 27004 14430 27016
rect 14737 27013 14749 27016
rect 14783 27013 14795 27047
rect 14737 27007 14795 27013
rect 15749 27047 15807 27053
rect 15749 27013 15761 27047
rect 15795 27044 15807 27047
rect 16574 27044 16580 27056
rect 15795 27016 16580 27044
rect 15795 27013 15807 27016
rect 15749 27007 15807 27013
rect 16574 27004 16580 27016
rect 16632 27004 16638 27056
rect 16666 27004 16672 27056
rect 16724 27044 16730 27056
rect 17681 27047 17739 27053
rect 17681 27044 17693 27047
rect 16724 27016 17693 27044
rect 16724 27004 16730 27016
rect 17681 27013 17693 27016
rect 17727 27013 17739 27047
rect 17681 27007 17739 27013
rect 19153 27047 19211 27053
rect 19153 27013 19165 27047
rect 19199 27044 19211 27047
rect 19426 27044 19432 27056
rect 19199 27016 19432 27044
rect 19199 27013 19211 27016
rect 19153 27007 19211 27013
rect 19426 27004 19432 27016
rect 19484 27004 19490 27056
rect 20088 27053 20116 27084
rect 20438 27072 20444 27084
rect 20496 27072 20502 27124
rect 23468 27115 23526 27121
rect 23468 27081 23480 27115
rect 23514 27112 23526 27115
rect 24670 27112 24676 27124
rect 23514 27084 24676 27112
rect 23514 27081 23526 27084
rect 23468 27075 23526 27081
rect 24670 27072 24676 27084
rect 24728 27072 24734 27124
rect 25130 27072 25136 27124
rect 25188 27112 25194 27124
rect 26237 27115 26295 27121
rect 26237 27112 26249 27115
rect 25188 27084 26249 27112
rect 25188 27072 25194 27084
rect 26237 27081 26249 27084
rect 26283 27081 26295 27115
rect 26237 27075 26295 27081
rect 20073 27047 20131 27053
rect 20073 27013 20085 27047
rect 20119 27013 20131 27047
rect 20073 27007 20131 27013
rect 20346 27004 20352 27056
rect 20404 27044 20410 27056
rect 20901 27047 20959 27053
rect 20901 27044 20913 27047
rect 20404 27016 20913 27044
rect 20404 27004 20410 27016
rect 20901 27013 20913 27016
rect 20947 27013 20959 27047
rect 20901 27007 20959 27013
rect 21266 27004 21272 27056
rect 21324 27004 21330 27056
rect 23934 27004 23940 27056
rect 23992 27044 23998 27056
rect 24489 27047 24547 27053
rect 24489 27044 24501 27047
rect 23992 27016 24501 27044
rect 23992 27004 23998 27016
rect 24489 27013 24501 27016
rect 24535 27013 24547 27047
rect 25038 27044 25044 27056
rect 24999 27016 25044 27044
rect 24489 27007 24547 27013
rect 25038 27004 25044 27016
rect 25096 27044 25102 27056
rect 26329 27047 26387 27053
rect 26329 27044 26341 27047
rect 25096 27016 26341 27044
rect 25096 27004 25102 27016
rect 26329 27013 26341 27016
rect 26375 27013 26387 27047
rect 26329 27007 26387 27013
rect 14645 26979 14703 26985
rect 14645 26945 14657 26979
rect 14691 26945 14703 26979
rect 14645 26939 14703 26945
rect 14921 26979 14979 26985
rect 14921 26945 14933 26979
rect 14967 26976 14979 26979
rect 15194 26976 15200 26988
rect 14967 26948 15200 26976
rect 14967 26945 14979 26948
rect 14921 26939 14979 26945
rect 12268 26880 14320 26908
rect 14660 26908 14688 26939
rect 15194 26936 15200 26948
rect 15252 26936 15258 26988
rect 15378 26976 15384 26988
rect 15339 26948 15384 26976
rect 15378 26936 15384 26948
rect 15436 26936 15442 26988
rect 15562 26976 15568 26988
rect 15523 26948 15568 26976
rect 15562 26936 15568 26948
rect 15620 26936 15626 26988
rect 16592 26976 16620 27004
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16592 26948 16865 26976
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 19242 26936 19248 26988
rect 19300 26976 19306 26988
rect 19337 26979 19395 26985
rect 19337 26976 19349 26979
rect 19300 26948 19349 26976
rect 19300 26936 19306 26948
rect 19337 26945 19349 26948
rect 19383 26945 19395 26979
rect 19337 26939 19395 26945
rect 19702 26936 19708 26988
rect 19760 26976 19766 26988
rect 19955 26979 20013 26985
rect 19955 26976 19967 26979
rect 19760 26948 19967 26976
rect 19760 26936 19766 26948
rect 19955 26945 19967 26948
rect 20001 26945 20013 26979
rect 20162 26976 20168 26988
rect 20123 26948 20168 26976
rect 19955 26939 20013 26945
rect 20162 26936 20168 26948
rect 20220 26936 20226 26988
rect 20254 26936 20260 26988
rect 20312 26976 20318 26988
rect 21085 26979 21143 26985
rect 20312 26948 20356 26976
rect 20312 26936 20318 26948
rect 21085 26945 21097 26979
rect 21131 26976 21143 26979
rect 21284 26976 21312 27004
rect 21821 26979 21879 26985
rect 21821 26976 21833 26979
rect 21131 26948 21833 26976
rect 21131 26945 21143 26948
rect 21085 26939 21143 26945
rect 21821 26945 21833 26948
rect 21867 26945 21879 26979
rect 22738 26976 22744 26988
rect 22699 26948 22744 26976
rect 21821 26939 21879 26945
rect 15010 26908 15016 26920
rect 14660 26880 15016 26908
rect 8754 26840 8760 26852
rect 7852 26812 8760 26840
rect 1854 26732 1860 26784
rect 1912 26772 1918 26784
rect 1949 26775 2007 26781
rect 1949 26772 1961 26775
rect 1912 26744 1961 26772
rect 1912 26732 1918 26744
rect 1949 26741 1961 26744
rect 1995 26741 2007 26775
rect 1949 26735 2007 26741
rect 5261 26775 5319 26781
rect 5261 26741 5273 26775
rect 5307 26772 5319 26775
rect 5350 26772 5356 26784
rect 5307 26744 5356 26772
rect 5307 26741 5319 26744
rect 5261 26735 5319 26741
rect 5350 26732 5356 26744
rect 5408 26732 5414 26784
rect 7852 26781 7880 26812
rect 8754 26800 8760 26812
rect 8812 26800 8818 26852
rect 10318 26840 10324 26852
rect 10231 26812 10324 26840
rect 10318 26800 10324 26812
rect 10376 26840 10382 26852
rect 12268 26840 12296 26880
rect 15010 26868 15016 26880
rect 15068 26868 15074 26920
rect 16945 26911 17003 26917
rect 16945 26877 16957 26911
rect 16991 26908 17003 26911
rect 18969 26911 19027 26917
rect 18969 26908 18981 26911
rect 16991 26880 18981 26908
rect 16991 26877 17003 26880
rect 16945 26871 17003 26877
rect 18969 26877 18981 26880
rect 19015 26877 19027 26911
rect 18969 26871 19027 26877
rect 19797 26911 19855 26917
rect 19797 26877 19809 26911
rect 19843 26908 19855 26911
rect 20898 26908 20904 26920
rect 19843 26880 20904 26908
rect 19843 26877 19855 26880
rect 19797 26871 19855 26877
rect 20898 26868 20904 26880
rect 20956 26908 20962 26920
rect 21100 26908 21128 26939
rect 22738 26936 22744 26948
rect 22796 26936 22802 26988
rect 23845 26979 23903 26985
rect 23845 26945 23857 26979
rect 23891 26976 23903 26979
rect 24854 26976 24860 26988
rect 23891 26948 24424 26976
rect 24815 26948 24860 26976
rect 23891 26945 23903 26948
rect 23845 26939 23903 26945
rect 21266 26908 21272 26920
rect 20956 26880 21128 26908
rect 21227 26880 21272 26908
rect 20956 26868 20962 26880
rect 21266 26868 21272 26880
rect 21324 26868 21330 26920
rect 24302 26908 24308 26920
rect 24263 26880 24308 26908
rect 24302 26868 24308 26880
rect 24360 26868 24366 26920
rect 24396 26908 24424 26948
rect 24854 26936 24860 26948
rect 24912 26936 24918 26988
rect 24949 26979 25007 26985
rect 24949 26945 24961 26979
rect 24995 26976 25007 26979
rect 26142 26976 26148 26988
rect 24995 26948 25029 26976
rect 26103 26948 26148 26976
rect 24995 26945 25007 26948
rect 24949 26939 25007 26945
rect 24578 26908 24584 26920
rect 24396 26880 24584 26908
rect 24578 26868 24584 26880
rect 24636 26908 24642 26920
rect 24964 26908 24992 26939
rect 26142 26936 26148 26948
rect 26200 26936 26206 26988
rect 25593 26911 25651 26917
rect 25593 26908 25605 26911
rect 24636 26880 25605 26908
rect 24636 26868 24642 26880
rect 25593 26877 25605 26880
rect 25639 26877 25651 26911
rect 25593 26871 25651 26877
rect 25777 26911 25835 26917
rect 25777 26877 25789 26911
rect 25823 26877 25835 26911
rect 25777 26871 25835 26877
rect 10376 26812 12296 26840
rect 10376 26800 10382 26812
rect 14826 26800 14832 26852
rect 14884 26840 14890 26852
rect 14921 26843 14979 26849
rect 14921 26840 14933 26843
rect 14884 26812 14933 26840
rect 14884 26800 14890 26812
rect 14921 26809 14933 26812
rect 14967 26809 14979 26843
rect 19610 26840 19616 26852
rect 14921 26803 14979 26809
rect 16960 26812 19616 26840
rect 7837 26775 7895 26781
rect 7837 26741 7849 26775
rect 7883 26741 7895 26775
rect 8294 26772 8300 26784
rect 8255 26744 8300 26772
rect 7837 26735 7895 26741
rect 8294 26732 8300 26744
rect 8352 26732 8358 26784
rect 10870 26772 10876 26784
rect 10831 26744 10876 26772
rect 10870 26732 10876 26744
rect 10928 26732 10934 26784
rect 12802 26732 12808 26784
rect 12860 26772 12866 26784
rect 13173 26775 13231 26781
rect 13173 26772 13185 26775
rect 12860 26744 13185 26772
rect 12860 26732 12866 26744
rect 13173 26741 13185 26744
rect 13219 26741 13231 26775
rect 14090 26772 14096 26784
rect 14051 26744 14096 26772
rect 13173 26735 13231 26741
rect 14090 26732 14096 26744
rect 14148 26732 14154 26784
rect 15286 26732 15292 26784
rect 15344 26772 15350 26784
rect 16960 26772 16988 26812
rect 19610 26800 19616 26812
rect 19668 26840 19674 26852
rect 19668 26812 22094 26840
rect 19668 26800 19674 26812
rect 17126 26772 17132 26784
rect 15344 26744 16988 26772
rect 17087 26744 17132 26772
rect 15344 26732 15350 26744
rect 17126 26732 17132 26744
rect 17184 26732 17190 26784
rect 18138 26732 18144 26784
rect 18196 26772 18202 26784
rect 18325 26775 18383 26781
rect 18325 26772 18337 26775
rect 18196 26744 18337 26772
rect 18196 26732 18202 26744
rect 18325 26741 18337 26744
rect 18371 26772 18383 26775
rect 18414 26772 18420 26784
rect 18371 26744 18420 26772
rect 18371 26741 18383 26744
rect 18325 26735 18383 26741
rect 18414 26732 18420 26744
rect 18472 26732 18478 26784
rect 19058 26732 19064 26784
rect 19116 26772 19122 26784
rect 21542 26772 21548 26784
rect 19116 26744 21548 26772
rect 19116 26732 19122 26744
rect 21542 26732 21548 26744
rect 21600 26732 21606 26784
rect 22066 26772 22094 26812
rect 22186 26800 22192 26852
rect 22244 26840 22250 26852
rect 25792 26840 25820 26871
rect 22244 26812 25820 26840
rect 22244 26800 22250 26812
rect 22370 26772 22376 26784
rect 22066 26744 22376 26772
rect 22370 26732 22376 26744
rect 22428 26732 22434 26784
rect 22554 26772 22560 26784
rect 22515 26744 22560 26772
rect 22554 26732 22560 26744
rect 22612 26732 22618 26784
rect 23290 26772 23296 26784
rect 23251 26744 23296 26772
rect 23290 26732 23296 26744
rect 23348 26732 23354 26784
rect 23477 26775 23535 26781
rect 23477 26741 23489 26775
rect 23523 26772 23535 26775
rect 24302 26772 24308 26784
rect 23523 26744 24308 26772
rect 23523 26741 23535 26744
rect 23477 26735 23535 26741
rect 24302 26732 24308 26744
rect 24360 26772 24366 26784
rect 25130 26772 25136 26784
rect 24360 26744 25136 26772
rect 24360 26732 24366 26744
rect 25130 26732 25136 26744
rect 25188 26732 25194 26784
rect 28626 26772 28632 26784
rect 28587 26744 28632 26772
rect 28626 26732 28632 26744
rect 28684 26732 28690 26784
rect 1104 26682 29440 26704
rect 1104 26630 4492 26682
rect 4544 26630 4556 26682
rect 4608 26630 4620 26682
rect 4672 26630 4684 26682
rect 4736 26630 4748 26682
rect 4800 26630 11576 26682
rect 11628 26630 11640 26682
rect 11692 26630 11704 26682
rect 11756 26630 11768 26682
rect 11820 26630 11832 26682
rect 11884 26630 18660 26682
rect 18712 26630 18724 26682
rect 18776 26630 18788 26682
rect 18840 26630 18852 26682
rect 18904 26630 18916 26682
rect 18968 26630 25744 26682
rect 25796 26630 25808 26682
rect 25860 26630 25872 26682
rect 25924 26630 25936 26682
rect 25988 26630 26000 26682
rect 26052 26630 29440 26682
rect 1104 26608 29440 26630
rect 1578 26568 1584 26580
rect 1539 26540 1584 26568
rect 1578 26528 1584 26540
rect 1636 26528 1642 26580
rect 5534 26568 5540 26580
rect 5495 26540 5540 26568
rect 5534 26528 5540 26540
rect 5592 26528 5598 26580
rect 7098 26568 7104 26580
rect 7059 26540 7104 26568
rect 7098 26528 7104 26540
rect 7156 26528 7162 26580
rect 7742 26528 7748 26580
rect 7800 26568 7806 26580
rect 10965 26571 11023 26577
rect 10965 26568 10977 26571
rect 7800 26540 10977 26568
rect 7800 26528 7806 26540
rect 10965 26537 10977 26540
rect 11011 26537 11023 26571
rect 11974 26568 11980 26580
rect 11935 26540 11980 26568
rect 10965 26531 11023 26537
rect 11974 26528 11980 26540
rect 12032 26528 12038 26580
rect 12342 26528 12348 26580
rect 12400 26568 12406 26580
rect 14366 26568 14372 26580
rect 12400 26540 14372 26568
rect 12400 26528 12406 26540
rect 14366 26528 14372 26540
rect 14424 26568 14430 26580
rect 14461 26571 14519 26577
rect 14461 26568 14473 26571
rect 14424 26540 14473 26568
rect 14424 26528 14430 26540
rect 14461 26537 14473 26540
rect 14507 26537 14519 26571
rect 15194 26568 15200 26580
rect 15155 26540 15200 26568
rect 14461 26531 14519 26537
rect 15194 26528 15200 26540
rect 15252 26528 15258 26580
rect 16298 26528 16304 26580
rect 16356 26568 16362 26580
rect 16485 26571 16543 26577
rect 16485 26568 16497 26571
rect 16356 26540 16497 26568
rect 16356 26528 16362 26540
rect 16485 26537 16497 26540
rect 16531 26537 16543 26571
rect 18049 26571 18107 26577
rect 18049 26568 18061 26571
rect 16485 26531 16543 26537
rect 16592 26540 18061 26568
rect 5718 26460 5724 26512
rect 5776 26500 5782 26512
rect 6273 26503 6331 26509
rect 6273 26500 6285 26503
rect 5776 26472 6285 26500
rect 5776 26460 5782 26472
rect 6273 26469 6285 26472
rect 6319 26500 6331 26503
rect 10042 26500 10048 26512
rect 6319 26472 10048 26500
rect 6319 26469 6331 26472
rect 6273 26463 6331 26469
rect 10042 26460 10048 26472
rect 10100 26460 10106 26512
rect 10505 26503 10563 26509
rect 10505 26469 10517 26503
rect 10551 26500 10563 26503
rect 10551 26472 12480 26500
rect 10551 26469 10563 26472
rect 10505 26463 10563 26469
rect 4985 26435 5043 26441
rect 4985 26401 4997 26435
rect 5031 26432 5043 26435
rect 8294 26432 8300 26444
rect 5031 26404 7236 26432
rect 5031 26401 5043 26404
rect 4985 26395 5043 26401
rect 4893 26367 4951 26373
rect 4893 26333 4905 26367
rect 4939 26333 4951 26367
rect 5074 26364 5080 26376
rect 5035 26336 5080 26364
rect 4893 26327 4951 26333
rect 4908 26296 4936 26327
rect 5074 26324 5080 26336
rect 5132 26324 5138 26376
rect 5534 26364 5540 26376
rect 5495 26336 5540 26364
rect 5534 26324 5540 26336
rect 5592 26324 5598 26376
rect 5718 26364 5724 26376
rect 5679 26336 5724 26364
rect 5718 26324 5724 26336
rect 5776 26324 5782 26376
rect 7006 26364 7012 26376
rect 6967 26336 7012 26364
rect 7006 26324 7012 26336
rect 7064 26324 7070 26376
rect 7208 26373 7236 26404
rect 7576 26404 8300 26432
rect 7576 26373 7604 26404
rect 8294 26392 8300 26404
rect 8352 26432 8358 26444
rect 8478 26432 8484 26444
rect 8352 26404 8484 26432
rect 8352 26392 8358 26404
rect 8478 26392 8484 26404
rect 8536 26392 8542 26444
rect 10870 26432 10876 26444
rect 9968 26404 10876 26432
rect 7193 26367 7251 26373
rect 7193 26333 7205 26367
rect 7239 26333 7251 26367
rect 7193 26327 7251 26333
rect 7561 26367 7619 26373
rect 7561 26333 7573 26367
rect 7607 26333 7619 26367
rect 7561 26327 7619 26333
rect 7837 26367 7895 26373
rect 7837 26333 7849 26367
rect 7883 26364 7895 26367
rect 8386 26364 8392 26376
rect 7883 26336 8392 26364
rect 7883 26333 7895 26336
rect 7837 26327 7895 26333
rect 8386 26324 8392 26336
rect 8444 26324 8450 26376
rect 9968 26373 9996 26404
rect 10870 26392 10876 26404
rect 10928 26392 10934 26444
rect 11238 26432 11244 26444
rect 11199 26404 11244 26432
rect 11238 26392 11244 26404
rect 11296 26392 11302 26444
rect 11333 26435 11391 26441
rect 11333 26401 11345 26435
rect 11379 26432 11391 26435
rect 12342 26432 12348 26444
rect 11379 26404 12348 26432
rect 11379 26401 11391 26404
rect 11333 26395 11391 26401
rect 12342 26392 12348 26404
rect 12400 26392 12406 26444
rect 9953 26367 10011 26373
rect 9953 26333 9965 26367
rect 9999 26333 10011 26367
rect 9953 26327 10011 26333
rect 10091 26367 10149 26373
rect 10091 26333 10103 26367
rect 10137 26333 10149 26367
rect 10091 26327 10149 26333
rect 10321 26367 10379 26373
rect 10321 26333 10333 26367
rect 10367 26364 10379 26367
rect 10502 26364 10508 26376
rect 10367 26336 10508 26364
rect 10367 26333 10379 26336
rect 10321 26327 10379 26333
rect 5350 26296 5356 26308
rect 4908 26268 5356 26296
rect 5350 26256 5356 26268
rect 5408 26256 5414 26308
rect 9493 26299 9551 26305
rect 9493 26265 9505 26299
rect 9539 26296 9551 26299
rect 9858 26296 9864 26308
rect 9539 26268 9864 26296
rect 9539 26265 9551 26268
rect 9493 26259 9551 26265
rect 9858 26256 9864 26268
rect 9916 26256 9922 26308
rect 7834 26188 7840 26240
rect 7892 26228 7898 26240
rect 8294 26228 8300 26240
rect 7892 26200 8300 26228
rect 7892 26188 7898 26200
rect 8294 26188 8300 26200
rect 8352 26188 8358 26240
rect 10106 26228 10134 26327
rect 10502 26324 10508 26336
rect 10560 26324 10566 26376
rect 11149 26367 11207 26373
rect 11149 26333 11161 26367
rect 11195 26333 11207 26367
rect 11149 26327 11207 26333
rect 11425 26367 11483 26373
rect 11425 26333 11437 26367
rect 11471 26364 11483 26367
rect 11514 26364 11520 26376
rect 11471 26336 11520 26364
rect 11471 26333 11483 26336
rect 11425 26327 11483 26333
rect 10226 26305 10232 26308
rect 10225 26259 10232 26305
rect 10284 26296 10290 26308
rect 11164 26296 11192 26327
rect 11514 26324 11520 26336
rect 11572 26364 11578 26376
rect 12161 26367 12219 26373
rect 12161 26364 12173 26367
rect 11572 26336 12173 26364
rect 11572 26324 11578 26336
rect 12161 26333 12173 26336
rect 12207 26333 12219 26367
rect 12161 26327 12219 26333
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12452 26373 12480 26472
rect 12710 26460 12716 26512
rect 12768 26500 12774 26512
rect 16592 26500 16620 26540
rect 18049 26537 18061 26540
rect 18095 26537 18107 26571
rect 18049 26531 18107 26537
rect 19794 26528 19800 26580
rect 19852 26568 19858 26580
rect 19981 26571 20039 26577
rect 19981 26568 19993 26571
rect 19852 26540 19993 26568
rect 19852 26528 19858 26540
rect 19981 26537 19993 26540
rect 20027 26537 20039 26571
rect 20990 26568 20996 26580
rect 20951 26540 20996 26568
rect 19981 26531 20039 26537
rect 20990 26528 20996 26540
rect 21048 26528 21054 26580
rect 22370 26528 22376 26580
rect 22428 26568 22434 26580
rect 22557 26571 22615 26577
rect 22557 26568 22569 26571
rect 22428 26540 22569 26568
rect 22428 26528 22434 26540
rect 22557 26537 22569 26540
rect 22603 26568 22615 26571
rect 23566 26568 23572 26580
rect 22603 26540 23572 26568
rect 22603 26537 22615 26540
rect 22557 26531 22615 26537
rect 23566 26528 23572 26540
rect 23624 26528 23630 26580
rect 23658 26528 23664 26580
rect 23716 26568 23722 26580
rect 24489 26571 24547 26577
rect 24489 26568 24501 26571
rect 23716 26540 24501 26568
rect 23716 26528 23722 26540
rect 24489 26537 24501 26540
rect 24535 26537 24547 26571
rect 24489 26531 24547 26537
rect 12768 26472 16620 26500
rect 16761 26503 16819 26509
rect 12768 26460 12774 26472
rect 16761 26469 16773 26503
rect 16807 26500 16819 26503
rect 17402 26500 17408 26512
rect 16807 26472 17408 26500
rect 16807 26469 16819 26472
rect 16761 26463 16819 26469
rect 17402 26460 17408 26472
rect 17460 26460 17466 26512
rect 18322 26460 18328 26512
rect 18380 26500 18386 26512
rect 18966 26500 18972 26512
rect 18380 26472 18972 26500
rect 18380 26460 18386 26472
rect 18966 26460 18972 26472
rect 19024 26460 19030 26512
rect 19426 26500 19432 26512
rect 19260 26472 19432 26500
rect 15562 26392 15568 26444
rect 15620 26432 15626 26444
rect 19260 26432 19288 26472
rect 19426 26460 19432 26472
rect 19484 26500 19490 26512
rect 20346 26500 20352 26512
rect 19484 26472 20352 26500
rect 19484 26460 19490 26472
rect 20346 26460 20352 26472
rect 20404 26460 20410 26512
rect 21542 26460 21548 26512
rect 21600 26500 21606 26512
rect 23106 26500 23112 26512
rect 21600 26472 22140 26500
rect 23067 26472 23112 26500
rect 21600 26460 21606 26472
rect 19886 26432 19892 26444
rect 15620 26404 18644 26432
rect 15620 26392 15626 26404
rect 12437 26367 12495 26373
rect 12308 26336 12353 26364
rect 12308 26324 12314 26336
rect 12437 26333 12449 26367
rect 12483 26333 12495 26367
rect 12437 26327 12495 26333
rect 12529 26367 12587 26373
rect 12529 26333 12541 26367
rect 12575 26364 12587 26367
rect 12802 26364 12808 26376
rect 12575 26336 12808 26364
rect 12575 26333 12587 26336
rect 12529 26327 12587 26333
rect 12802 26324 12808 26336
rect 12860 26324 12866 26376
rect 15286 26364 15292 26376
rect 13372 26336 15292 26364
rect 12710 26296 12716 26308
rect 10284 26268 10325 26296
rect 11164 26268 12716 26296
rect 10226 26256 10232 26259
rect 10284 26256 10290 26268
rect 12710 26256 12716 26268
rect 12768 26256 12774 26308
rect 10410 26228 10416 26240
rect 10106 26200 10416 26228
rect 10410 26188 10416 26200
rect 10468 26188 10474 26240
rect 12250 26188 12256 26240
rect 12308 26228 12314 26240
rect 13372 26228 13400 26336
rect 15286 26324 15292 26336
rect 15344 26324 15350 26376
rect 15381 26367 15439 26373
rect 15381 26333 15393 26367
rect 15427 26364 15439 26367
rect 15654 26364 15660 26376
rect 15427 26336 15660 26364
rect 15427 26333 15439 26336
rect 15381 26327 15439 26333
rect 15654 26324 15660 26336
rect 15712 26324 15718 26376
rect 15749 26367 15807 26373
rect 15749 26333 15761 26367
rect 15795 26364 15807 26367
rect 15838 26364 15844 26376
rect 15795 26336 15844 26364
rect 15795 26333 15807 26336
rect 15749 26327 15807 26333
rect 15838 26324 15844 26336
rect 15896 26324 15902 26376
rect 16666 26364 16672 26376
rect 16627 26336 16672 26364
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 16853 26367 16911 26373
rect 16853 26333 16865 26367
rect 16899 26333 16911 26367
rect 16853 26327 16911 26333
rect 14090 26296 14096 26308
rect 14003 26268 14096 26296
rect 14090 26256 14096 26268
rect 14148 26256 14154 26308
rect 14274 26296 14280 26308
rect 14235 26268 14280 26296
rect 14274 26256 14280 26268
rect 14332 26256 14338 26308
rect 15473 26299 15531 26305
rect 15473 26265 15485 26299
rect 15519 26265 15531 26299
rect 15473 26259 15531 26265
rect 15565 26299 15623 26305
rect 15565 26265 15577 26299
rect 15611 26296 15623 26299
rect 16574 26296 16580 26308
rect 15611 26268 16580 26296
rect 15611 26265 15623 26268
rect 15565 26259 15623 26265
rect 12308 26200 13400 26228
rect 13541 26231 13599 26237
rect 12308 26188 12314 26200
rect 13541 26197 13553 26231
rect 13587 26228 13599 26231
rect 13906 26228 13912 26240
rect 13587 26200 13912 26228
rect 13587 26197 13599 26200
rect 13541 26191 13599 26197
rect 13906 26188 13912 26200
rect 13964 26188 13970 26240
rect 14108 26228 14136 26256
rect 15488 26228 15516 26259
rect 16574 26256 16580 26268
rect 16632 26256 16638 26308
rect 16868 26296 16896 26327
rect 16942 26324 16948 26376
rect 17000 26364 17006 26376
rect 17126 26364 17132 26376
rect 17000 26336 17045 26364
rect 17087 26336 17132 26364
rect 17000 26324 17006 26336
rect 17126 26324 17132 26336
rect 17184 26324 17190 26376
rect 18233 26367 18291 26373
rect 18233 26333 18245 26367
rect 18279 26333 18291 26367
rect 18233 26327 18291 26333
rect 18138 26296 18144 26308
rect 16868 26268 18144 26296
rect 18138 26256 18144 26268
rect 18196 26256 18202 26308
rect 15654 26228 15660 26240
rect 14108 26200 15660 26228
rect 15654 26188 15660 26200
rect 15712 26228 15718 26240
rect 16206 26228 16212 26240
rect 15712 26200 16212 26228
rect 15712 26188 15718 26200
rect 16206 26188 16212 26200
rect 16264 26188 16270 26240
rect 18248 26228 18276 26327
rect 18322 26324 18328 26376
rect 18380 26364 18386 26376
rect 18616 26373 18644 26404
rect 18800 26404 19473 26432
rect 18574 26367 18644 26373
rect 18380 26336 18425 26364
rect 18380 26324 18386 26336
rect 18574 26333 18586 26367
rect 18620 26336 18644 26367
rect 18693 26367 18751 26373
rect 18620 26333 18632 26336
rect 18574 26327 18632 26333
rect 18693 26333 18705 26367
rect 18739 26358 18751 26367
rect 18800 26358 18828 26404
rect 18739 26333 18828 26358
rect 18693 26330 18828 26333
rect 18693 26327 18751 26330
rect 19058 26324 19064 26376
rect 19116 26364 19122 26376
rect 19445 26373 19473 26404
rect 19536 26404 19892 26432
rect 19337 26367 19395 26373
rect 19337 26364 19349 26367
rect 19116 26336 19349 26364
rect 19116 26324 19122 26336
rect 19337 26333 19349 26336
rect 19383 26333 19395 26367
rect 19337 26327 19395 26333
rect 19430 26367 19488 26373
rect 19430 26333 19442 26367
rect 19476 26333 19488 26367
rect 19430 26327 19488 26333
rect 18417 26299 18475 26305
rect 18417 26265 18429 26299
rect 18463 26296 18475 26299
rect 18874 26296 18880 26308
rect 18463 26268 18880 26296
rect 18463 26265 18475 26268
rect 18417 26259 18475 26265
rect 18874 26256 18880 26268
rect 18932 26256 18938 26308
rect 18966 26256 18972 26308
rect 19024 26296 19030 26308
rect 19536 26296 19564 26404
rect 19886 26392 19892 26404
rect 19944 26432 19950 26444
rect 22112 26441 22140 26472
rect 23106 26460 23112 26472
rect 23164 26460 23170 26512
rect 22097 26435 22155 26441
rect 19944 26404 20944 26432
rect 19944 26392 19950 26404
rect 19610 26324 19616 26376
rect 19668 26364 19674 26376
rect 19668 26336 19713 26364
rect 19668 26324 19674 26336
rect 19794 26324 19800 26376
rect 19852 26373 19858 26376
rect 19852 26364 19860 26373
rect 20438 26364 20444 26376
rect 19852 26336 19897 26364
rect 20399 26336 20444 26364
rect 19852 26327 19860 26336
rect 19852 26324 19858 26327
rect 20438 26324 20444 26336
rect 20496 26324 20502 26376
rect 20806 26364 20812 26376
rect 20767 26336 20812 26364
rect 20806 26324 20812 26336
rect 20864 26324 20870 26376
rect 19702 26296 19708 26308
rect 19024 26268 19564 26296
rect 19663 26268 19708 26296
rect 19024 26256 19030 26268
rect 19702 26256 19708 26268
rect 19760 26256 19766 26308
rect 20625 26299 20683 26305
rect 20625 26265 20637 26299
rect 20671 26265 20683 26299
rect 20625 26259 20683 26265
rect 20717 26299 20775 26305
rect 20717 26265 20729 26299
rect 20763 26296 20775 26299
rect 20916 26296 20944 26404
rect 22097 26401 22109 26435
rect 22143 26432 22155 26435
rect 22186 26432 22192 26444
rect 22143 26404 22192 26432
rect 22143 26401 22155 26404
rect 22097 26395 22155 26401
rect 22186 26392 22192 26404
rect 22244 26392 22250 26444
rect 24854 26392 24860 26444
rect 24912 26432 24918 26444
rect 26142 26432 26148 26444
rect 24912 26404 26148 26432
rect 24912 26392 24918 26404
rect 24397 26367 24455 26373
rect 24397 26333 24409 26367
rect 24443 26364 24455 26367
rect 24486 26364 24492 26376
rect 24443 26336 24492 26364
rect 24443 26333 24455 26336
rect 24397 26327 24455 26333
rect 24486 26324 24492 26336
rect 24544 26324 24550 26376
rect 25792 26373 25820 26404
rect 26142 26392 26148 26404
rect 26200 26392 26206 26444
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26364 24639 26367
rect 25777 26367 25835 26373
rect 24627 26336 25636 26364
rect 24627 26333 24639 26336
rect 24581 26327 24639 26333
rect 20763 26268 20944 26296
rect 20763 26265 20775 26268
rect 20717 26259 20775 26265
rect 19242 26228 19248 26240
rect 18248 26200 19248 26228
rect 19242 26188 19248 26200
rect 19300 26228 19306 26240
rect 20640 26228 20668 26259
rect 25608 26240 25636 26336
rect 25777 26333 25789 26367
rect 25823 26333 25835 26367
rect 25958 26364 25964 26376
rect 25919 26336 25964 26364
rect 25777 26327 25835 26333
rect 25958 26324 25964 26336
rect 26016 26324 26022 26376
rect 28261 26299 28319 26305
rect 28261 26265 28273 26299
rect 28307 26296 28319 26299
rect 28350 26296 28356 26308
rect 28307 26268 28356 26296
rect 28307 26265 28319 26268
rect 28261 26259 28319 26265
rect 28350 26256 28356 26268
rect 28408 26256 28414 26308
rect 28626 26296 28632 26308
rect 28587 26268 28632 26296
rect 28626 26256 28632 26268
rect 28684 26256 28690 26308
rect 19300 26200 20668 26228
rect 19300 26188 19306 26200
rect 21358 26188 21364 26240
rect 21416 26228 21422 26240
rect 21453 26231 21511 26237
rect 21453 26228 21465 26231
rect 21416 26200 21465 26228
rect 21416 26188 21422 26200
rect 21453 26197 21465 26200
rect 21499 26197 21511 26231
rect 21453 26191 21511 26197
rect 25590 26188 25596 26240
rect 25648 26228 25654 26240
rect 25777 26231 25835 26237
rect 25777 26228 25789 26231
rect 25648 26200 25789 26228
rect 25648 26188 25654 26200
rect 25777 26197 25789 26200
rect 25823 26197 25835 26231
rect 25777 26191 25835 26197
rect 1104 26138 29600 26160
rect 1104 26086 8034 26138
rect 8086 26086 8098 26138
rect 8150 26086 8162 26138
rect 8214 26086 8226 26138
rect 8278 26086 8290 26138
rect 8342 26086 15118 26138
rect 15170 26086 15182 26138
rect 15234 26086 15246 26138
rect 15298 26086 15310 26138
rect 15362 26086 15374 26138
rect 15426 26086 22202 26138
rect 22254 26086 22266 26138
rect 22318 26086 22330 26138
rect 22382 26086 22394 26138
rect 22446 26086 22458 26138
rect 22510 26086 29286 26138
rect 29338 26086 29350 26138
rect 29402 26086 29414 26138
rect 29466 26086 29478 26138
rect 29530 26086 29542 26138
rect 29594 26086 29600 26138
rect 1104 26064 29600 26086
rect 5074 25984 5080 26036
rect 5132 26024 5138 26036
rect 5169 26027 5227 26033
rect 5169 26024 5181 26027
rect 5132 25996 5181 26024
rect 5132 25984 5138 25996
rect 5169 25993 5181 25996
rect 5215 25993 5227 26027
rect 5169 25987 5227 25993
rect 7006 25984 7012 26036
rect 7064 25984 7070 26036
rect 7190 26024 7196 26036
rect 7151 25996 7196 26024
rect 7190 25984 7196 25996
rect 7248 25984 7254 26036
rect 8754 26024 8760 26036
rect 8715 25996 8760 26024
rect 8754 25984 8760 25996
rect 8812 25984 8818 26036
rect 9858 25984 9864 26036
rect 9916 26024 9922 26036
rect 10502 26024 10508 26036
rect 9916 25996 10508 26024
rect 9916 25984 9922 25996
rect 10502 25984 10508 25996
rect 10560 25984 10566 26036
rect 11514 26024 11520 26036
rect 11475 25996 11520 26024
rect 11514 25984 11520 25996
rect 11572 25984 11578 26036
rect 13354 26024 13360 26036
rect 13315 25996 13360 26024
rect 13354 25984 13360 25996
rect 13412 25984 13418 26036
rect 13906 25984 13912 26036
rect 13964 26024 13970 26036
rect 14274 26024 14280 26036
rect 13964 25996 14280 26024
rect 13964 25984 13970 25996
rect 14274 25984 14280 25996
rect 14332 25984 14338 26036
rect 15010 26024 15016 26036
rect 14971 25996 15016 26024
rect 15010 25984 15016 25996
rect 15068 25984 15074 26036
rect 19242 25984 19248 26036
rect 19300 26024 19306 26036
rect 19429 26027 19487 26033
rect 19429 26024 19441 26027
rect 19300 25996 19441 26024
rect 19300 25984 19306 25996
rect 19429 25993 19441 25996
rect 19475 25993 19487 26027
rect 19429 25987 19487 25993
rect 19521 26027 19579 26033
rect 19521 25993 19533 26027
rect 19567 26024 19579 26027
rect 20254 26024 20260 26036
rect 19567 25996 20260 26024
rect 19567 25993 19579 25996
rect 19521 25987 19579 25993
rect 20254 25984 20260 25996
rect 20312 26024 20318 26036
rect 20717 26027 20775 26033
rect 20717 26024 20729 26027
rect 20312 25996 20729 26024
rect 20312 25984 20318 25996
rect 20717 25993 20729 25996
rect 20763 26024 20775 26027
rect 20806 26024 20812 26036
rect 20763 25996 20812 26024
rect 20763 25993 20775 25996
rect 20717 25987 20775 25993
rect 20806 25984 20812 25996
rect 20864 25984 20870 26036
rect 23566 25984 23572 26036
rect 23624 26024 23630 26036
rect 23661 26027 23719 26033
rect 23661 26024 23673 26027
rect 23624 25996 23673 26024
rect 23624 25984 23630 25996
rect 23661 25993 23673 25996
rect 23707 25993 23719 26027
rect 23661 25987 23719 25993
rect 25860 26027 25918 26033
rect 25860 25993 25872 26027
rect 25906 26024 25918 26027
rect 26142 26024 26148 26036
rect 25906 25996 26148 26024
rect 25906 25993 25918 25996
rect 25860 25987 25918 25993
rect 5537 25959 5595 25965
rect 5537 25956 5549 25959
rect 5092 25928 5549 25956
rect 5092 25900 5120 25928
rect 5537 25925 5549 25928
rect 5583 25956 5595 25959
rect 7024 25956 7052 25984
rect 7653 25959 7711 25965
rect 7653 25956 7665 25959
rect 5583 25928 6914 25956
rect 7024 25928 7665 25956
rect 5583 25925 5595 25928
rect 5537 25919 5595 25925
rect 4338 25888 4344 25900
rect 4299 25860 4344 25888
rect 4338 25848 4344 25860
rect 4396 25848 4402 25900
rect 5074 25848 5080 25900
rect 5132 25848 5138 25900
rect 5258 25848 5264 25900
rect 5316 25888 5322 25900
rect 5353 25891 5411 25897
rect 5353 25888 5365 25891
rect 5316 25860 5365 25888
rect 5316 25848 5322 25860
rect 5353 25857 5365 25860
rect 5399 25857 5411 25891
rect 5353 25851 5411 25857
rect 5626 25848 5632 25900
rect 5684 25888 5690 25900
rect 5684 25860 5729 25888
rect 5684 25848 5690 25860
rect 4246 25820 4252 25832
rect 4207 25792 4252 25820
rect 4246 25780 4252 25792
rect 4304 25780 4310 25832
rect 6730 25820 6736 25832
rect 6691 25792 6736 25820
rect 6730 25780 6736 25792
rect 6788 25780 6794 25832
rect 6886 25820 6914 25928
rect 7653 25925 7665 25928
rect 7699 25925 7711 25959
rect 10962 25956 10968 25968
rect 7653 25919 7711 25925
rect 8128 25928 10968 25956
rect 7006 25888 7012 25900
rect 6967 25860 7012 25888
rect 7006 25848 7012 25860
rect 7064 25848 7070 25900
rect 7190 25848 7196 25900
rect 7248 25888 7254 25900
rect 7834 25888 7840 25900
rect 7248 25860 7840 25888
rect 7248 25848 7254 25860
rect 7834 25848 7840 25860
rect 7892 25848 7898 25900
rect 7926 25848 7932 25900
rect 7984 25888 7990 25900
rect 8128 25897 8156 25928
rect 10962 25916 10968 25928
rect 11020 25916 11026 25968
rect 12066 25956 12072 25968
rect 11716 25928 12072 25956
rect 8021 25891 8079 25897
rect 8021 25888 8033 25891
rect 7984 25860 8033 25888
rect 7984 25848 7990 25860
rect 8021 25857 8033 25860
rect 8067 25857 8079 25891
rect 8021 25851 8079 25857
rect 8113 25891 8171 25897
rect 8113 25857 8125 25891
rect 8159 25857 8171 25891
rect 8113 25851 8171 25857
rect 8386 25848 8392 25900
rect 8444 25888 8450 25900
rect 8662 25888 8668 25900
rect 8444 25860 8668 25888
rect 8444 25848 8450 25860
rect 8662 25848 8668 25860
rect 8720 25848 8726 25900
rect 8849 25891 8907 25897
rect 8849 25857 8861 25891
rect 8895 25888 8907 25891
rect 9214 25888 9220 25900
rect 8895 25860 9220 25888
rect 8895 25857 8907 25860
rect 8849 25851 8907 25857
rect 9214 25848 9220 25860
rect 9272 25888 9278 25900
rect 9309 25891 9367 25897
rect 9309 25888 9321 25891
rect 9272 25860 9321 25888
rect 9272 25848 9278 25860
rect 9309 25857 9321 25860
rect 9355 25857 9367 25891
rect 10410 25888 10416 25900
rect 10371 25860 10416 25888
rect 9309 25851 9367 25857
rect 10410 25848 10416 25860
rect 10468 25848 10474 25900
rect 11716 25897 11744 25928
rect 12066 25916 12072 25928
rect 12124 25956 12130 25968
rect 12618 25956 12624 25968
rect 12124 25928 12624 25956
rect 12124 25916 12130 25928
rect 12618 25916 12624 25928
rect 12676 25916 12682 25968
rect 13541 25959 13599 25965
rect 13541 25925 13553 25959
rect 13587 25956 13599 25959
rect 13998 25956 14004 25968
rect 13587 25928 14004 25956
rect 13587 25925 13599 25928
rect 13541 25919 13599 25925
rect 13998 25916 14004 25928
rect 14056 25916 14062 25968
rect 16758 25956 16764 25968
rect 15166 25928 16764 25956
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 12526 25888 12532 25900
rect 11701 25851 11759 25857
rect 11808 25860 12532 25888
rect 11808 25820 11836 25860
rect 12526 25848 12532 25860
rect 12584 25848 12590 25900
rect 13725 25891 13783 25897
rect 13725 25857 13737 25891
rect 13771 25888 13783 25891
rect 14090 25888 14096 25900
rect 13771 25860 14096 25888
rect 13771 25857 13783 25860
rect 13725 25851 13783 25857
rect 14090 25848 14096 25860
rect 14148 25848 14154 25900
rect 14366 25888 14372 25900
rect 14327 25860 14372 25888
rect 14366 25848 14372 25860
rect 14424 25848 14430 25900
rect 14458 25848 14464 25900
rect 14516 25888 14522 25900
rect 15166 25897 15194 25928
rect 16758 25916 16764 25928
rect 16816 25916 16822 25968
rect 18322 25916 18328 25968
rect 18380 25956 18386 25968
rect 18874 25956 18880 25968
rect 18380 25928 18880 25956
rect 18380 25916 18386 25928
rect 18874 25916 18880 25928
rect 18932 25956 18938 25968
rect 19797 25959 19855 25965
rect 19797 25956 19809 25959
rect 18932 25928 19809 25956
rect 18932 25916 18938 25928
rect 19797 25925 19809 25928
rect 19843 25956 19855 25959
rect 20438 25956 20444 25968
rect 19843 25928 20444 25956
rect 19843 25925 19855 25928
rect 19797 25919 19855 25925
rect 20438 25916 20444 25928
rect 20496 25916 20502 25968
rect 21358 25956 21364 25968
rect 20732 25928 21364 25956
rect 15153 25891 15211 25897
rect 15153 25888 15165 25891
rect 14516 25860 15165 25888
rect 14516 25848 14522 25860
rect 15153 25857 15165 25860
rect 15199 25857 15211 25891
rect 15286 25888 15292 25900
rect 15247 25860 15292 25888
rect 15153 25851 15211 25857
rect 15286 25848 15292 25860
rect 15344 25848 15350 25900
rect 15381 25891 15439 25897
rect 15381 25857 15393 25891
rect 15427 25857 15439 25891
rect 15562 25888 15568 25900
rect 15523 25860 15568 25888
rect 15381 25851 15439 25857
rect 6886 25792 11836 25820
rect 11885 25823 11943 25829
rect 11885 25789 11897 25823
rect 11931 25820 11943 25823
rect 12158 25820 12164 25832
rect 11931 25792 12164 25820
rect 11931 25789 11943 25792
rect 11885 25783 11943 25789
rect 4709 25755 4767 25761
rect 4709 25721 4721 25755
rect 4755 25752 4767 25755
rect 5534 25752 5540 25764
rect 4755 25724 5540 25752
rect 4755 25721 4767 25724
rect 4709 25715 4767 25721
rect 5534 25712 5540 25724
rect 5592 25712 5598 25764
rect 7929 25755 7987 25761
rect 7929 25721 7941 25755
rect 7975 25752 7987 25755
rect 8202 25752 8208 25764
rect 7975 25724 8208 25752
rect 7975 25721 7987 25724
rect 7929 25715 7987 25721
rect 8202 25712 8208 25724
rect 8260 25712 8266 25764
rect 10226 25712 10232 25764
rect 10284 25752 10290 25764
rect 10965 25755 11023 25761
rect 10965 25752 10977 25755
rect 10284 25724 10977 25752
rect 10284 25712 10290 25724
rect 10965 25721 10977 25724
rect 11011 25752 11023 25755
rect 11900 25752 11928 25783
rect 12158 25780 12164 25792
rect 12216 25780 12222 25832
rect 14826 25780 14832 25832
rect 14884 25820 14890 25832
rect 15396 25820 15424 25851
rect 15562 25848 15568 25860
rect 15620 25848 15626 25900
rect 15657 25891 15715 25897
rect 15657 25857 15669 25891
rect 15703 25857 15715 25891
rect 15657 25851 15715 25857
rect 15672 25820 15700 25851
rect 19150 25848 19156 25900
rect 19208 25888 19214 25900
rect 19245 25891 19303 25897
rect 19245 25888 19257 25891
rect 19208 25860 19257 25888
rect 19208 25848 19214 25860
rect 19245 25857 19257 25860
rect 19291 25857 19303 25891
rect 19245 25851 19303 25857
rect 19613 25891 19671 25897
rect 19613 25857 19625 25891
rect 19659 25857 19671 25891
rect 19613 25851 19671 25857
rect 17218 25820 17224 25832
rect 14884 25792 15424 25820
rect 15626 25792 17224 25820
rect 14884 25780 14890 25792
rect 11011 25724 11928 25752
rect 14461 25755 14519 25761
rect 11011 25721 11023 25724
rect 10965 25715 11023 25721
rect 14461 25721 14473 25755
rect 14507 25752 14519 25755
rect 15378 25752 15384 25764
rect 14507 25724 15384 25752
rect 14507 25721 14519 25724
rect 14461 25715 14519 25721
rect 15378 25712 15384 25724
rect 15436 25712 15442 25764
rect 6822 25684 6828 25696
rect 6783 25656 6828 25684
rect 6822 25644 6828 25656
rect 6880 25644 6886 25696
rect 12250 25644 12256 25696
rect 12308 25684 12314 25696
rect 12805 25687 12863 25693
rect 12805 25684 12817 25687
rect 12308 25656 12817 25684
rect 12308 25644 12314 25656
rect 12805 25653 12817 25656
rect 12851 25653 12863 25687
rect 12805 25647 12863 25653
rect 12894 25644 12900 25696
rect 12952 25684 12958 25696
rect 15626 25684 15654 25792
rect 17218 25780 17224 25792
rect 17276 25780 17282 25832
rect 18046 25780 18052 25832
rect 18104 25820 18110 25832
rect 18325 25823 18383 25829
rect 18325 25820 18337 25823
rect 18104 25792 18337 25820
rect 18104 25780 18110 25792
rect 18325 25789 18337 25792
rect 18371 25789 18383 25823
rect 19628 25820 19656 25851
rect 19702 25848 19708 25900
rect 19760 25888 19766 25900
rect 20732 25897 20760 25928
rect 21358 25916 21364 25928
rect 21416 25956 21422 25968
rect 22373 25959 22431 25965
rect 22373 25956 22385 25959
rect 21416 25928 22385 25956
rect 21416 25916 21422 25928
rect 22373 25925 22385 25928
rect 22419 25925 22431 25959
rect 22373 25919 22431 25925
rect 20717 25891 20775 25897
rect 20717 25888 20729 25891
rect 19760 25860 20729 25888
rect 19760 25848 19766 25860
rect 20717 25857 20729 25860
rect 20763 25857 20775 25891
rect 20898 25888 20904 25900
rect 20859 25860 20904 25888
rect 20717 25851 20775 25857
rect 20898 25848 20904 25860
rect 20956 25848 20962 25900
rect 23676 25888 23704 25987
rect 26142 25984 26148 25996
rect 26200 25984 26206 26036
rect 24946 25916 24952 25968
rect 25004 25956 25010 25968
rect 25958 25956 25964 25968
rect 25004 25928 25964 25956
rect 25004 25916 25010 25928
rect 25958 25916 25964 25928
rect 26016 25956 26022 25968
rect 26237 25959 26295 25965
rect 26237 25956 26249 25959
rect 26016 25928 26249 25956
rect 26016 25916 26022 25928
rect 26237 25925 26249 25928
rect 26283 25956 26295 25959
rect 26878 25956 26884 25968
rect 26283 25928 26884 25956
rect 26283 25925 26295 25928
rect 26237 25919 26295 25925
rect 26878 25916 26884 25928
rect 26936 25916 26942 25968
rect 25593 25891 25651 25897
rect 25593 25888 25605 25891
rect 23676 25860 25605 25888
rect 25593 25857 25605 25860
rect 25639 25857 25651 25891
rect 25593 25851 25651 25857
rect 19886 25820 19892 25832
rect 19628 25792 19892 25820
rect 18325 25783 18383 25789
rect 19886 25780 19892 25792
rect 19944 25780 19950 25832
rect 16758 25752 16764 25764
rect 16671 25724 16764 25752
rect 16758 25712 16764 25724
rect 16816 25752 16822 25764
rect 19794 25752 19800 25764
rect 16816 25724 19800 25752
rect 16816 25712 16822 25724
rect 19794 25712 19800 25724
rect 19852 25752 19858 25764
rect 21821 25755 21879 25761
rect 21821 25752 21833 25755
rect 19852 25724 21833 25752
rect 19852 25712 19858 25724
rect 21821 25721 21833 25724
rect 21867 25752 21879 25755
rect 22738 25752 22744 25764
rect 21867 25724 22744 25752
rect 21867 25721 21879 25724
rect 21821 25715 21879 25721
rect 22738 25712 22744 25724
rect 22796 25752 22802 25764
rect 23290 25752 23296 25764
rect 22796 25724 23296 25752
rect 22796 25712 22802 25724
rect 23290 25712 23296 25724
rect 23348 25712 23354 25764
rect 27706 25712 27712 25764
rect 27764 25752 27770 25764
rect 28629 25755 28687 25761
rect 28629 25752 28641 25755
rect 27764 25724 28641 25752
rect 27764 25712 27770 25724
rect 28629 25721 28641 25724
rect 28675 25721 28687 25755
rect 28629 25715 28687 25721
rect 12952 25656 15654 25684
rect 17865 25687 17923 25693
rect 12952 25644 12958 25656
rect 17865 25653 17877 25687
rect 17911 25684 17923 25687
rect 18230 25684 18236 25696
rect 17911 25656 18236 25684
rect 17911 25653 17923 25656
rect 17865 25647 17923 25653
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 25869 25687 25927 25693
rect 25869 25653 25881 25687
rect 25915 25684 25927 25687
rect 26142 25684 26148 25696
rect 25915 25656 26148 25684
rect 25915 25653 25927 25656
rect 25869 25647 25927 25653
rect 26142 25644 26148 25656
rect 26200 25644 26206 25696
rect 27614 25684 27620 25696
rect 27575 25656 27620 25684
rect 27614 25644 27620 25656
rect 27672 25644 27678 25696
rect 28169 25687 28227 25693
rect 28169 25653 28181 25687
rect 28215 25684 28227 25687
rect 28534 25684 28540 25696
rect 28215 25656 28540 25684
rect 28215 25653 28227 25656
rect 28169 25647 28227 25653
rect 28534 25644 28540 25656
rect 28592 25644 28598 25696
rect 1104 25594 29440 25616
rect 1104 25542 4492 25594
rect 4544 25542 4556 25594
rect 4608 25542 4620 25594
rect 4672 25542 4684 25594
rect 4736 25542 4748 25594
rect 4800 25542 11576 25594
rect 11628 25542 11640 25594
rect 11692 25542 11704 25594
rect 11756 25542 11768 25594
rect 11820 25542 11832 25594
rect 11884 25542 18660 25594
rect 18712 25542 18724 25594
rect 18776 25542 18788 25594
rect 18840 25542 18852 25594
rect 18904 25542 18916 25594
rect 18968 25542 25744 25594
rect 25796 25542 25808 25594
rect 25860 25542 25872 25594
rect 25924 25542 25936 25594
rect 25988 25542 26000 25594
rect 26052 25542 29440 25594
rect 1104 25520 29440 25542
rect 4246 25440 4252 25492
rect 4304 25480 4310 25492
rect 4341 25483 4399 25489
rect 4341 25480 4353 25483
rect 4304 25452 4353 25480
rect 4304 25440 4310 25452
rect 4341 25449 4353 25452
rect 4387 25449 4399 25483
rect 5258 25480 5264 25492
rect 5219 25452 5264 25480
rect 4341 25443 4399 25449
rect 5258 25440 5264 25452
rect 5316 25440 5322 25492
rect 7006 25440 7012 25492
rect 7064 25480 7070 25492
rect 7101 25483 7159 25489
rect 7101 25480 7113 25483
rect 7064 25452 7113 25480
rect 7064 25440 7070 25452
rect 7101 25449 7113 25452
rect 7147 25449 7159 25483
rect 8202 25480 8208 25492
rect 8163 25452 8208 25480
rect 7101 25443 7159 25449
rect 8202 25440 8208 25452
rect 8260 25440 8266 25492
rect 13541 25483 13599 25489
rect 13541 25449 13553 25483
rect 13587 25480 13599 25483
rect 14090 25480 14096 25492
rect 13587 25452 14096 25480
rect 13587 25449 13599 25452
rect 13541 25443 13599 25449
rect 14090 25440 14096 25452
rect 14148 25440 14154 25492
rect 15562 25440 15568 25492
rect 15620 25480 15626 25492
rect 15749 25483 15807 25489
rect 15749 25480 15761 25483
rect 15620 25452 15761 25480
rect 15620 25440 15626 25452
rect 15749 25449 15761 25452
rect 15795 25449 15807 25483
rect 15749 25443 15807 25449
rect 16114 25440 16120 25492
rect 16172 25480 16178 25492
rect 17037 25483 17095 25489
rect 17037 25480 17049 25483
rect 16172 25452 17049 25480
rect 16172 25440 16178 25452
rect 17037 25449 17049 25452
rect 17083 25449 17095 25483
rect 17402 25480 17408 25492
rect 17315 25452 17408 25480
rect 17037 25443 17095 25449
rect 17402 25440 17408 25452
rect 17460 25480 17466 25492
rect 18230 25480 18236 25492
rect 17460 25452 18236 25480
rect 17460 25440 17466 25452
rect 18230 25440 18236 25452
rect 18288 25440 18294 25492
rect 19242 25480 19248 25492
rect 19203 25452 19248 25480
rect 19242 25440 19248 25452
rect 19300 25440 19306 25492
rect 20809 25483 20867 25489
rect 20809 25449 20821 25483
rect 20855 25480 20867 25483
rect 20898 25480 20904 25492
rect 20855 25452 20904 25480
rect 20855 25449 20867 25452
rect 20809 25443 20867 25449
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 21358 25440 21364 25492
rect 21416 25480 21422 25492
rect 21453 25483 21511 25489
rect 21453 25480 21465 25483
rect 21416 25452 21465 25480
rect 21416 25440 21422 25452
rect 21453 25449 21465 25452
rect 21499 25449 21511 25483
rect 21453 25443 21511 25449
rect 22373 25483 22431 25489
rect 22373 25449 22385 25483
rect 22419 25480 22431 25483
rect 23106 25480 23112 25492
rect 22419 25452 23112 25480
rect 22419 25449 22431 25452
rect 22373 25443 22431 25449
rect 23106 25440 23112 25452
rect 23164 25440 23170 25492
rect 23290 25440 23296 25492
rect 23348 25480 23354 25492
rect 23477 25483 23535 25489
rect 23477 25480 23489 25483
rect 23348 25452 23489 25480
rect 23348 25440 23354 25452
rect 23477 25449 23489 25452
rect 23523 25449 23535 25483
rect 26878 25480 26884 25492
rect 26839 25452 26884 25480
rect 23477 25443 23535 25449
rect 26878 25440 26884 25452
rect 26936 25440 26942 25492
rect 27614 25440 27620 25492
rect 27672 25480 27678 25492
rect 28442 25480 28448 25492
rect 27672 25452 28448 25480
rect 27672 25440 27678 25452
rect 28442 25440 28448 25452
rect 28500 25480 28506 25492
rect 28537 25483 28595 25489
rect 28537 25480 28549 25483
rect 28500 25452 28549 25480
rect 28500 25440 28506 25452
rect 28537 25449 28549 25452
rect 28583 25449 28595 25483
rect 28537 25443 28595 25449
rect 7742 25304 7748 25356
rect 7800 25344 7806 25356
rect 7800 25316 8064 25344
rect 7800 25304 7806 25316
rect 4614 25276 4620 25288
rect 4575 25248 4620 25276
rect 4614 25236 4620 25248
rect 4672 25236 4678 25288
rect 5074 25276 5080 25288
rect 5035 25248 5080 25276
rect 5074 25236 5080 25248
rect 5132 25236 5138 25288
rect 5258 25276 5264 25288
rect 5219 25248 5264 25276
rect 5258 25236 5264 25248
rect 5316 25236 5322 25288
rect 6822 25236 6828 25288
rect 6880 25276 6886 25288
rect 7377 25279 7435 25285
rect 7377 25276 7389 25279
rect 6880 25248 7389 25276
rect 6880 25236 6886 25248
rect 7377 25245 7389 25248
rect 7423 25245 7435 25279
rect 7834 25276 7840 25288
rect 7795 25248 7840 25276
rect 7377 25239 7435 25245
rect 4341 25211 4399 25217
rect 4341 25177 4353 25211
rect 4387 25208 4399 25211
rect 5276 25208 5304 25236
rect 4387 25180 5304 25208
rect 7101 25211 7159 25217
rect 4387 25177 4399 25180
rect 4341 25171 4399 25177
rect 7101 25177 7113 25211
rect 7147 25208 7159 25211
rect 7190 25208 7196 25220
rect 7147 25180 7196 25208
rect 7147 25177 7159 25180
rect 7101 25171 7159 25177
rect 7190 25168 7196 25180
rect 7248 25168 7254 25220
rect 7392 25208 7420 25239
rect 7834 25236 7840 25248
rect 7892 25236 7898 25288
rect 8036 25285 8064 25316
rect 8021 25279 8079 25285
rect 8021 25245 8033 25279
rect 8067 25245 8079 25279
rect 8220 25276 8248 25440
rect 25038 25412 25044 25424
rect 17420 25384 25044 25412
rect 8662 25304 8668 25356
rect 8720 25344 8726 25356
rect 9677 25347 9735 25353
rect 9677 25344 9689 25347
rect 8720 25316 9689 25344
rect 8720 25304 8726 25316
rect 9677 25313 9689 25316
rect 9723 25344 9735 25347
rect 16666 25344 16672 25356
rect 9723 25316 16672 25344
rect 9723 25313 9735 25316
rect 9677 25307 9735 25313
rect 16666 25304 16672 25316
rect 16724 25344 16730 25356
rect 17313 25347 17371 25353
rect 17313 25344 17325 25347
rect 16724 25316 17325 25344
rect 16724 25304 16730 25316
rect 17313 25313 17325 25316
rect 17359 25313 17371 25347
rect 17313 25307 17371 25313
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8220 25248 8953 25276
rect 8021 25239 8079 25245
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25276 9183 25279
rect 9306 25276 9312 25288
rect 9171 25248 9312 25276
rect 9171 25245 9183 25248
rect 9125 25239 9183 25245
rect 9306 25236 9312 25248
rect 9364 25236 9370 25288
rect 12158 25276 12164 25288
rect 12071 25248 12164 25276
rect 12158 25236 12164 25248
rect 12216 25276 12222 25288
rect 13538 25276 13544 25288
rect 12216 25248 13544 25276
rect 12216 25236 12222 25248
rect 13538 25236 13544 25248
rect 13596 25236 13602 25288
rect 15381 25279 15439 25285
rect 15381 25276 15393 25279
rect 14844 25248 15393 25276
rect 9033 25211 9091 25217
rect 9033 25208 9045 25211
rect 7392 25180 9045 25208
rect 9033 25177 9045 25180
rect 9079 25177 9091 25211
rect 10410 25208 10416 25220
rect 10371 25180 10416 25208
rect 9033 25171 9091 25177
rect 10410 25168 10416 25180
rect 10468 25208 10474 25220
rect 11241 25211 11299 25217
rect 11241 25208 11253 25211
rect 10468 25180 11253 25208
rect 10468 25168 10474 25180
rect 11241 25177 11253 25180
rect 11287 25208 11299 25211
rect 12250 25208 12256 25220
rect 11287 25180 12256 25208
rect 11287 25177 11299 25180
rect 11241 25171 11299 25177
rect 12250 25168 12256 25180
rect 12308 25168 12314 25220
rect 4525 25143 4583 25149
rect 4525 25109 4537 25143
rect 4571 25140 4583 25143
rect 5074 25140 5080 25152
rect 4571 25112 5080 25140
rect 4571 25109 4583 25112
rect 4525 25103 4583 25109
rect 5074 25100 5080 25112
rect 5132 25100 5138 25152
rect 6454 25100 6460 25152
rect 6512 25140 6518 25152
rect 6730 25140 6736 25152
rect 6512 25112 6736 25140
rect 6512 25100 6518 25112
rect 6730 25100 6736 25112
rect 6788 25140 6794 25152
rect 7285 25143 7343 25149
rect 7285 25140 7297 25143
rect 6788 25112 7297 25140
rect 6788 25100 6794 25112
rect 7285 25109 7297 25112
rect 7331 25109 7343 25143
rect 7285 25103 7343 25109
rect 10689 25143 10747 25149
rect 10689 25109 10701 25143
rect 10735 25140 10747 25143
rect 10870 25140 10876 25152
rect 10735 25112 10876 25140
rect 10735 25109 10747 25112
rect 10689 25103 10747 25109
rect 10870 25100 10876 25112
rect 10928 25100 10934 25152
rect 12526 25100 12532 25152
rect 12584 25140 12590 25152
rect 12713 25143 12771 25149
rect 12713 25140 12725 25143
rect 12584 25112 12725 25140
rect 12584 25100 12590 25112
rect 12713 25109 12725 25112
rect 12759 25109 12771 25143
rect 12713 25103 12771 25109
rect 13906 25100 13912 25152
rect 13964 25140 13970 25152
rect 14844 25149 14872 25248
rect 15381 25245 15393 25248
rect 15427 25245 15439 25279
rect 15381 25239 15439 25245
rect 15565 25279 15623 25285
rect 15565 25245 15577 25279
rect 15611 25276 15623 25279
rect 15654 25276 15660 25288
rect 15611 25248 15660 25276
rect 15611 25245 15623 25248
rect 15565 25239 15623 25245
rect 15654 25236 15660 25248
rect 15712 25276 15718 25288
rect 15712 25248 16344 25276
rect 15712 25236 15718 25248
rect 16316 25149 16344 25248
rect 17328 25208 17356 25307
rect 17420 25285 17448 25384
rect 25038 25372 25044 25384
rect 25096 25372 25102 25424
rect 22002 25344 22008 25356
rect 19628 25316 22008 25344
rect 17405 25279 17463 25285
rect 17405 25245 17417 25279
rect 17451 25245 17463 25279
rect 17405 25239 17463 25245
rect 19429 25279 19487 25285
rect 19429 25245 19441 25279
rect 19475 25276 19487 25279
rect 19518 25276 19524 25288
rect 19475 25248 19524 25276
rect 19475 25245 19487 25248
rect 19429 25239 19487 25245
rect 19518 25236 19524 25248
rect 19576 25236 19582 25288
rect 19628 25285 19656 25316
rect 22002 25304 22008 25316
rect 22060 25304 22066 25356
rect 22830 25344 22836 25356
rect 22388 25316 22836 25344
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 19705 25279 19763 25285
rect 19705 25245 19717 25279
rect 19751 25276 19763 25279
rect 19794 25276 19800 25288
rect 19751 25248 19800 25276
rect 19751 25245 19763 25248
rect 19705 25239 19763 25245
rect 19794 25236 19800 25248
rect 19852 25236 19858 25288
rect 22388 25276 22416 25316
rect 22830 25304 22836 25316
rect 22888 25304 22894 25356
rect 24673 25347 24731 25353
rect 24673 25313 24685 25347
rect 24719 25344 24731 25347
rect 26142 25344 26148 25356
rect 24719 25316 26148 25344
rect 24719 25313 24731 25316
rect 24673 25307 24731 25313
rect 22554 25276 22560 25288
rect 20180 25248 22416 25276
rect 22515 25248 22560 25276
rect 17678 25208 17684 25220
rect 17328 25180 17684 25208
rect 17678 25168 17684 25180
rect 17736 25208 17742 25220
rect 17865 25211 17923 25217
rect 17865 25208 17877 25211
rect 17736 25180 17877 25208
rect 17736 25168 17742 25180
rect 17865 25177 17877 25180
rect 17911 25177 17923 25211
rect 19536 25208 19564 25236
rect 20180 25217 20208 25248
rect 22554 25236 22560 25248
rect 22612 25236 22618 25288
rect 24578 25276 24584 25288
rect 24539 25248 24584 25276
rect 24578 25236 24584 25248
rect 24636 25236 24642 25288
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25276 24823 25279
rect 25130 25276 25136 25288
rect 24811 25248 25136 25276
rect 24811 25245 24823 25248
rect 24765 25239 24823 25245
rect 25130 25236 25136 25248
rect 25188 25236 25194 25288
rect 25682 25276 25688 25288
rect 25643 25248 25688 25276
rect 25682 25236 25688 25248
rect 25740 25236 25746 25288
rect 26068 25285 26096 25316
rect 26142 25304 26148 25316
rect 26200 25304 26206 25356
rect 25869 25279 25927 25285
rect 25869 25245 25881 25279
rect 25915 25245 25927 25279
rect 25869 25239 25927 25245
rect 26053 25279 26111 25285
rect 26053 25245 26065 25279
rect 26099 25245 26111 25279
rect 26053 25239 26111 25245
rect 20165 25211 20223 25217
rect 20165 25208 20177 25211
rect 19536 25180 20177 25208
rect 17865 25171 17923 25177
rect 20165 25177 20177 25180
rect 20211 25177 20223 25211
rect 20165 25171 20223 25177
rect 20990 25168 20996 25220
rect 21048 25208 21054 25220
rect 21266 25208 21272 25220
rect 21048 25180 21272 25208
rect 21048 25168 21054 25180
rect 21266 25168 21272 25180
rect 21324 25208 21330 25220
rect 21361 25211 21419 25217
rect 21361 25208 21373 25211
rect 21324 25180 21373 25208
rect 21324 25168 21330 25180
rect 21361 25177 21373 25180
rect 21407 25177 21419 25211
rect 21361 25171 21419 25177
rect 23382 25168 23388 25220
rect 23440 25208 23446 25220
rect 25225 25211 25283 25217
rect 25225 25208 25237 25211
rect 23440 25180 25237 25208
rect 23440 25168 23446 25180
rect 25225 25177 25237 25180
rect 25271 25177 25283 25211
rect 25225 25171 25283 25177
rect 25590 25168 25596 25220
rect 25648 25208 25654 25220
rect 25884 25208 25912 25239
rect 25648 25180 25912 25208
rect 26068 25208 26096 25239
rect 26234 25236 26240 25288
rect 26292 25276 26298 25288
rect 26292 25248 27108 25276
rect 26292 25236 26298 25248
rect 27080 25217 27108 25248
rect 26849 25211 26907 25217
rect 26849 25208 26861 25211
rect 26068 25180 26861 25208
rect 25648 25168 25654 25180
rect 26849 25177 26861 25180
rect 26895 25177 26907 25211
rect 26849 25171 26907 25177
rect 27065 25211 27123 25217
rect 27065 25177 27077 25211
rect 27111 25177 27123 25211
rect 27065 25171 27123 25177
rect 14093 25143 14151 25149
rect 14093 25140 14105 25143
rect 13964 25112 14105 25140
rect 13964 25100 13970 25112
rect 14093 25109 14105 25112
rect 14139 25140 14151 25143
rect 14829 25143 14887 25149
rect 14829 25140 14841 25143
rect 14139 25112 14841 25140
rect 14139 25109 14151 25112
rect 14093 25103 14151 25109
rect 14829 25109 14841 25112
rect 14875 25109 14887 25143
rect 14829 25103 14887 25109
rect 16301 25143 16359 25149
rect 16301 25109 16313 25143
rect 16347 25140 16359 25143
rect 16390 25140 16396 25152
rect 16347 25112 16396 25140
rect 16347 25109 16359 25112
rect 16301 25103 16359 25109
rect 16390 25100 16396 25112
rect 16448 25100 16454 25152
rect 18230 25100 18236 25152
rect 18288 25140 18294 25152
rect 18417 25143 18475 25149
rect 18417 25140 18429 25143
rect 18288 25112 18429 25140
rect 18288 25100 18294 25112
rect 18417 25109 18429 25112
rect 18463 25109 18475 25143
rect 18417 25103 18475 25109
rect 22922 25100 22928 25152
rect 22980 25140 22986 25152
rect 26697 25143 26755 25149
rect 26697 25140 26709 25143
rect 22980 25112 26709 25140
rect 22980 25100 22986 25112
rect 26697 25109 26709 25112
rect 26743 25109 26755 25143
rect 26697 25103 26755 25109
rect 28077 25143 28135 25149
rect 28077 25109 28089 25143
rect 28123 25140 28135 25143
rect 28258 25140 28264 25152
rect 28123 25112 28264 25140
rect 28123 25109 28135 25112
rect 28077 25103 28135 25109
rect 28258 25100 28264 25112
rect 28316 25100 28322 25152
rect 1104 25050 29600 25072
rect 1104 24998 8034 25050
rect 8086 24998 8098 25050
rect 8150 24998 8162 25050
rect 8214 24998 8226 25050
rect 8278 24998 8290 25050
rect 8342 24998 15118 25050
rect 15170 24998 15182 25050
rect 15234 24998 15246 25050
rect 15298 24998 15310 25050
rect 15362 24998 15374 25050
rect 15426 24998 22202 25050
rect 22254 24998 22266 25050
rect 22318 24998 22330 25050
rect 22382 24998 22394 25050
rect 22446 24998 22458 25050
rect 22510 24998 29286 25050
rect 29338 24998 29350 25050
rect 29402 24998 29414 25050
rect 29466 24998 29478 25050
rect 29530 24998 29542 25050
rect 29594 24998 29600 25050
rect 1104 24976 29600 24998
rect 4982 24896 4988 24948
rect 5040 24936 5046 24948
rect 5166 24936 5172 24948
rect 5040 24908 5172 24936
rect 5040 24896 5046 24908
rect 5166 24896 5172 24908
rect 5224 24896 5230 24948
rect 7926 24896 7932 24948
rect 7984 24936 7990 24948
rect 8113 24939 8171 24945
rect 8113 24936 8125 24939
rect 7984 24908 8125 24936
rect 7984 24896 7990 24908
rect 8113 24905 8125 24908
rect 8159 24905 8171 24939
rect 8113 24899 8171 24905
rect 10870 24896 10876 24948
rect 10928 24936 10934 24948
rect 14826 24936 14832 24948
rect 10928 24908 14832 24936
rect 10928 24896 10934 24908
rect 14826 24896 14832 24908
rect 14884 24896 14890 24948
rect 22465 24939 22523 24945
rect 22465 24905 22477 24939
rect 22511 24936 22523 24939
rect 22554 24936 22560 24948
rect 22511 24908 22560 24936
rect 22511 24905 22523 24908
rect 22465 24899 22523 24905
rect 22554 24896 22560 24908
rect 22612 24896 22618 24948
rect 25682 24896 25688 24948
rect 25740 24936 25746 24948
rect 25869 24939 25927 24945
rect 25869 24936 25881 24939
rect 25740 24908 25881 24936
rect 25740 24896 25746 24908
rect 25869 24905 25881 24908
rect 25915 24905 25927 24939
rect 25869 24899 25927 24905
rect 7834 24868 7840 24880
rect 6886 24840 7840 24868
rect 1394 24800 1400 24812
rect 1355 24772 1400 24800
rect 1394 24760 1400 24772
rect 1452 24760 1458 24812
rect 4525 24803 4583 24809
rect 4525 24769 4537 24803
rect 4571 24769 4583 24803
rect 4525 24763 4583 24769
rect 4709 24803 4767 24809
rect 4709 24769 4721 24803
rect 4755 24800 4767 24803
rect 4890 24800 4896 24812
rect 4755 24772 4896 24800
rect 4755 24769 4767 24772
rect 4709 24763 4767 24769
rect 4540 24732 4568 24763
rect 4890 24760 4896 24772
rect 4948 24800 4954 24812
rect 5258 24800 5264 24812
rect 4948 24772 5264 24800
rect 4948 24760 4954 24772
rect 5258 24760 5264 24772
rect 5316 24800 5322 24812
rect 6886 24800 6914 24840
rect 7834 24828 7840 24840
rect 7892 24868 7898 24880
rect 15470 24868 15476 24880
rect 7892 24840 8248 24868
rect 7892 24828 7898 24840
rect 8220 24812 8248 24840
rect 13832 24840 15476 24868
rect 5316 24772 6914 24800
rect 5316 24760 5322 24772
rect 7742 24760 7748 24812
rect 7800 24800 7806 24812
rect 8021 24803 8079 24809
rect 8021 24800 8033 24803
rect 7800 24772 8033 24800
rect 7800 24760 7806 24772
rect 8021 24769 8033 24772
rect 8067 24769 8079 24803
rect 8202 24800 8208 24812
rect 8163 24772 8208 24800
rect 8021 24763 8079 24769
rect 8202 24760 8208 24772
rect 8260 24760 8266 24812
rect 12802 24800 12808 24812
rect 12268 24772 12808 24800
rect 4614 24732 4620 24744
rect 4527 24704 4620 24732
rect 4614 24692 4620 24704
rect 4672 24732 4678 24744
rect 5074 24732 5080 24744
rect 4672 24704 5080 24732
rect 4672 24692 4678 24704
rect 5074 24692 5080 24704
rect 5132 24732 5138 24744
rect 11422 24732 11428 24744
rect 5132 24704 11428 24732
rect 5132 24692 5138 24704
rect 11422 24692 11428 24704
rect 11480 24692 11486 24744
rect 9490 24624 9496 24676
rect 9548 24664 9554 24676
rect 10321 24667 10379 24673
rect 10321 24664 10333 24667
rect 9548 24636 10333 24664
rect 9548 24624 9554 24636
rect 10321 24633 10333 24636
rect 10367 24664 10379 24667
rect 12268 24664 12296 24772
rect 12802 24760 12808 24772
rect 12860 24760 12866 24812
rect 13081 24803 13139 24809
rect 13081 24769 13093 24803
rect 13127 24769 13139 24803
rect 13081 24763 13139 24769
rect 12529 24735 12587 24741
rect 12529 24701 12541 24735
rect 12575 24732 12587 24735
rect 13096 24732 13124 24763
rect 13262 24760 13268 24812
rect 13320 24800 13326 24812
rect 13449 24803 13507 24809
rect 13449 24800 13461 24803
rect 13320 24772 13461 24800
rect 13320 24760 13326 24772
rect 13449 24769 13461 24772
rect 13495 24800 13507 24803
rect 13832 24800 13860 24840
rect 15470 24828 15476 24840
rect 15528 24828 15534 24880
rect 22649 24871 22707 24877
rect 22649 24837 22661 24871
rect 22695 24868 22707 24871
rect 22922 24868 22928 24880
rect 22695 24840 22928 24868
rect 22695 24837 22707 24840
rect 22649 24831 22707 24837
rect 22922 24828 22928 24840
rect 22980 24828 22986 24880
rect 13495 24772 13860 24800
rect 13495 24769 13507 24772
rect 13449 24763 13507 24769
rect 13906 24760 13912 24812
rect 13964 24800 13970 24812
rect 21818 24800 21824 24812
rect 13964 24772 14057 24800
rect 21779 24772 21824 24800
rect 13964 24760 13970 24772
rect 21818 24760 21824 24772
rect 21876 24760 21882 24812
rect 22833 24803 22891 24809
rect 22833 24769 22845 24803
rect 22879 24800 22891 24803
rect 23382 24800 23388 24812
rect 22879 24772 23388 24800
rect 22879 24769 22891 24772
rect 22833 24763 22891 24769
rect 23382 24760 23388 24772
rect 23440 24760 23446 24812
rect 24946 24760 24952 24812
rect 25004 24800 25010 24812
rect 25504 24809 25562 24815
rect 25682 24809 25688 24812
rect 25225 24803 25283 24809
rect 25225 24800 25237 24803
rect 25004 24772 25237 24800
rect 25004 24760 25010 24772
rect 25225 24769 25237 24772
rect 25271 24769 25283 24803
rect 25225 24763 25283 24769
rect 25409 24803 25467 24809
rect 25409 24769 25421 24803
rect 25455 24769 25467 24803
rect 25504 24775 25516 24809
rect 25550 24775 25562 24809
rect 25504 24769 25562 24775
rect 25639 24803 25688 24809
rect 25639 24769 25651 24803
rect 25685 24769 25688 24803
rect 25409 24763 25467 24769
rect 13354 24732 13360 24744
rect 12575 24704 13360 24732
rect 12575 24701 12587 24704
rect 12529 24695 12587 24701
rect 13354 24692 13360 24704
rect 13412 24732 13418 24744
rect 13924 24732 13952 24760
rect 13412 24704 13952 24732
rect 13412 24692 13418 24704
rect 13998 24692 14004 24744
rect 14056 24732 14062 24744
rect 14056 24704 14101 24732
rect 14056 24692 14062 24704
rect 25314 24692 25320 24744
rect 25372 24732 25378 24744
rect 25424 24732 25452 24763
rect 25372 24704 25452 24732
rect 25372 24692 25378 24704
rect 14734 24664 14740 24676
rect 10367 24636 12296 24664
rect 12406 24636 14740 24664
rect 10367 24633 10379 24636
rect 10321 24627 10379 24633
rect 1578 24596 1584 24608
rect 1539 24568 1584 24596
rect 1578 24556 1584 24568
rect 1636 24556 1642 24608
rect 4893 24599 4951 24605
rect 4893 24565 4905 24599
rect 4939 24596 4951 24599
rect 5534 24596 5540 24608
rect 4939 24568 5540 24596
rect 4939 24565 4951 24568
rect 4893 24559 4951 24565
rect 5534 24556 5540 24568
rect 5592 24556 5598 24608
rect 7190 24556 7196 24608
rect 7248 24596 7254 24608
rect 7469 24599 7527 24605
rect 7469 24596 7481 24599
rect 7248 24568 7481 24596
rect 7248 24556 7254 24568
rect 7469 24565 7481 24568
rect 7515 24565 7527 24599
rect 7469 24559 7527 24565
rect 8846 24556 8852 24608
rect 8904 24596 8910 24608
rect 9217 24599 9275 24605
rect 9217 24596 9229 24599
rect 8904 24568 9229 24596
rect 8904 24556 8910 24568
rect 9217 24565 9229 24568
rect 9263 24565 9275 24599
rect 9217 24559 9275 24565
rect 10042 24556 10048 24608
rect 10100 24596 10106 24608
rect 12406 24596 12434 24636
rect 14734 24624 14740 24636
rect 14792 24624 14798 24676
rect 10100 24568 12434 24596
rect 10100 24556 10106 24568
rect 17218 24556 17224 24608
rect 17276 24596 17282 24608
rect 18785 24599 18843 24605
rect 18785 24596 18797 24599
rect 17276 24568 18797 24596
rect 17276 24556 17282 24568
rect 18785 24565 18797 24568
rect 18831 24596 18843 24599
rect 19058 24596 19064 24608
rect 18831 24568 19064 24596
rect 18831 24565 18843 24568
rect 18785 24559 18843 24565
rect 19058 24556 19064 24568
rect 19116 24556 19122 24608
rect 19521 24599 19579 24605
rect 19521 24565 19533 24599
rect 19567 24596 19579 24599
rect 19794 24596 19800 24608
rect 19567 24568 19800 24596
rect 19567 24565 19579 24568
rect 19521 24559 19579 24565
rect 19794 24556 19800 24568
rect 19852 24596 19858 24608
rect 19981 24599 20039 24605
rect 19981 24596 19993 24599
rect 19852 24568 19993 24596
rect 19852 24556 19858 24568
rect 19981 24565 19993 24568
rect 20027 24565 20039 24599
rect 19981 24559 20039 24565
rect 24210 24556 24216 24608
rect 24268 24596 24274 24608
rect 24305 24599 24363 24605
rect 24305 24596 24317 24599
rect 24268 24568 24317 24596
rect 24268 24556 24274 24568
rect 24305 24565 24317 24568
rect 24351 24596 24363 24599
rect 25519 24596 25547 24769
rect 25639 24763 25688 24769
rect 25682 24760 25688 24763
rect 25740 24760 25746 24812
rect 26329 24667 26387 24673
rect 26329 24633 26341 24667
rect 26375 24664 26387 24667
rect 27525 24667 27583 24673
rect 27525 24664 27537 24667
rect 26375 24636 27537 24664
rect 26375 24633 26387 24636
rect 26329 24627 26387 24633
rect 27525 24633 27537 24636
rect 27571 24633 27583 24667
rect 27525 24627 27583 24633
rect 25590 24596 25596 24608
rect 24351 24568 25596 24596
rect 24351 24565 24363 24568
rect 24305 24559 24363 24565
rect 25590 24556 25596 24568
rect 25648 24596 25654 24608
rect 26344 24596 26372 24627
rect 26970 24596 26976 24608
rect 25648 24568 26372 24596
rect 26931 24568 26976 24596
rect 25648 24556 25654 24568
rect 26970 24556 26976 24568
rect 27028 24556 27034 24608
rect 28445 24599 28503 24605
rect 28445 24565 28457 24599
rect 28491 24596 28503 24599
rect 28534 24596 28540 24608
rect 28491 24568 28540 24596
rect 28491 24565 28503 24568
rect 28445 24559 28503 24565
rect 28534 24556 28540 24568
rect 28592 24556 28598 24608
rect 1104 24506 29440 24528
rect 1104 24454 4492 24506
rect 4544 24454 4556 24506
rect 4608 24454 4620 24506
rect 4672 24454 4684 24506
rect 4736 24454 4748 24506
rect 4800 24454 11576 24506
rect 11628 24454 11640 24506
rect 11692 24454 11704 24506
rect 11756 24454 11768 24506
rect 11820 24454 11832 24506
rect 11884 24454 18660 24506
rect 18712 24454 18724 24506
rect 18776 24454 18788 24506
rect 18840 24454 18852 24506
rect 18904 24454 18916 24506
rect 18968 24454 25744 24506
rect 25796 24454 25808 24506
rect 25860 24454 25872 24506
rect 25924 24454 25936 24506
rect 25988 24454 26000 24506
rect 26052 24454 29440 24506
rect 1104 24432 29440 24454
rect 1394 24392 1400 24404
rect 1355 24364 1400 24392
rect 1394 24352 1400 24364
rect 1452 24352 1458 24404
rect 1578 24352 1584 24404
rect 1636 24392 1642 24404
rect 10042 24392 10048 24404
rect 1636 24364 10048 24392
rect 1636 24352 1642 24364
rect 10042 24352 10048 24364
rect 10100 24352 10106 24404
rect 10413 24395 10471 24401
rect 10413 24361 10425 24395
rect 10459 24361 10471 24395
rect 10413 24355 10471 24361
rect 5626 24324 5632 24336
rect 5587 24296 5632 24324
rect 5626 24284 5632 24296
rect 5684 24284 5690 24336
rect 5644 24256 5672 24284
rect 10428 24256 10456 24355
rect 11422 24352 11428 24404
rect 11480 24392 11486 24404
rect 11609 24395 11667 24401
rect 11609 24392 11621 24395
rect 11480 24364 11621 24392
rect 11480 24352 11486 24364
rect 11609 24361 11621 24364
rect 11655 24361 11667 24395
rect 12526 24392 12532 24404
rect 12439 24364 12532 24392
rect 11609 24355 11667 24361
rect 12526 24352 12532 24364
rect 12584 24392 12590 24404
rect 19242 24392 19248 24404
rect 12584 24364 19248 24392
rect 12584 24352 12590 24364
rect 19242 24352 19248 24364
rect 19300 24352 19306 24404
rect 23750 24392 23756 24404
rect 23663 24364 23756 24392
rect 23750 24352 23756 24364
rect 23808 24392 23814 24404
rect 27890 24392 27896 24404
rect 23808 24364 27896 24392
rect 23808 24352 23814 24364
rect 27890 24352 27896 24364
rect 27948 24352 27954 24404
rect 18601 24327 18659 24333
rect 18601 24293 18613 24327
rect 18647 24324 18659 24327
rect 22557 24327 22615 24333
rect 22557 24324 22569 24327
rect 18647 24296 22569 24324
rect 18647 24293 18659 24296
rect 18601 24287 18659 24293
rect 22557 24293 22569 24296
rect 22603 24293 22615 24327
rect 23768 24324 23796 24352
rect 22557 24287 22615 24293
rect 22848 24296 23796 24324
rect 24857 24327 24915 24333
rect 4264 24228 5672 24256
rect 9232 24228 10456 24256
rect 4154 24148 4160 24200
rect 4212 24188 4218 24200
rect 4264 24197 4292 24228
rect 4249 24191 4307 24197
rect 4249 24188 4261 24191
rect 4212 24160 4261 24188
rect 4212 24148 4218 24160
rect 4249 24157 4261 24160
rect 4295 24157 4307 24191
rect 4249 24151 4307 24157
rect 4338 24148 4344 24200
rect 4396 24188 4402 24200
rect 4433 24191 4491 24197
rect 4433 24188 4445 24191
rect 4396 24160 4445 24188
rect 4396 24148 4402 24160
rect 4433 24157 4445 24160
rect 4479 24157 4491 24191
rect 4890 24188 4896 24200
rect 4851 24160 4896 24188
rect 4433 24151 4491 24157
rect 4890 24148 4896 24160
rect 4948 24148 4954 24200
rect 5074 24188 5080 24200
rect 5035 24160 5080 24188
rect 5074 24148 5080 24160
rect 5132 24148 5138 24200
rect 5534 24188 5540 24200
rect 5495 24160 5540 24188
rect 5534 24148 5540 24160
rect 5592 24148 5598 24200
rect 5721 24191 5779 24197
rect 5721 24157 5733 24191
rect 5767 24157 5779 24191
rect 5721 24151 5779 24157
rect 7653 24191 7711 24197
rect 7653 24157 7665 24191
rect 7699 24188 7711 24191
rect 8846 24188 8852 24200
rect 7699 24160 8852 24188
rect 7699 24157 7711 24160
rect 7653 24151 7711 24157
rect 4614 24080 4620 24132
rect 4672 24120 4678 24132
rect 4985 24123 5043 24129
rect 4985 24120 4997 24123
rect 4672 24092 4997 24120
rect 4672 24080 4678 24092
rect 4985 24089 4997 24092
rect 5031 24120 5043 24123
rect 5736 24120 5764 24151
rect 8846 24148 8852 24160
rect 8904 24148 8910 24200
rect 9030 24148 9036 24200
rect 9088 24188 9094 24200
rect 9232 24197 9260 24228
rect 12710 24216 12716 24268
rect 12768 24256 12774 24268
rect 12768 24228 18276 24256
rect 12768 24216 12774 24228
rect 9217 24191 9275 24197
rect 9217 24188 9229 24191
rect 9088 24160 9229 24188
rect 9088 24148 9094 24160
rect 9217 24157 9229 24160
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 9306 24148 9312 24200
rect 9364 24188 9370 24200
rect 10137 24191 10195 24197
rect 9364 24160 9409 24188
rect 9364 24148 9370 24160
rect 10137 24157 10149 24191
rect 10183 24188 10195 24191
rect 10226 24188 10232 24200
rect 10183 24160 10232 24188
rect 10183 24157 10195 24160
rect 10137 24151 10195 24157
rect 10226 24148 10232 24160
rect 10284 24148 10290 24200
rect 11793 24191 11851 24197
rect 11793 24157 11805 24191
rect 11839 24188 11851 24191
rect 12986 24188 12992 24200
rect 11839 24160 12992 24188
rect 11839 24157 11851 24160
rect 11793 24151 11851 24157
rect 12986 24148 12992 24160
rect 13044 24148 13050 24200
rect 13998 24148 14004 24200
rect 14056 24188 14062 24200
rect 14553 24191 14611 24197
rect 14553 24188 14565 24191
rect 14056 24160 14565 24188
rect 14056 24148 14062 24160
rect 14553 24157 14565 24160
rect 14599 24157 14611 24191
rect 14553 24151 14611 24157
rect 5031 24092 5764 24120
rect 7009 24123 7067 24129
rect 5031 24089 5043 24092
rect 4985 24083 5043 24089
rect 7009 24089 7021 24123
rect 7055 24120 7067 24123
rect 8113 24123 8171 24129
rect 8113 24120 8125 24123
rect 7055 24092 8125 24120
rect 7055 24089 7067 24092
rect 7009 24083 7067 24089
rect 8113 24089 8125 24092
rect 8159 24089 8171 24123
rect 8113 24083 8171 24089
rect 4246 24012 4252 24064
rect 4304 24052 4310 24064
rect 4341 24055 4399 24061
rect 4341 24052 4353 24055
rect 4304 24024 4353 24052
rect 4304 24012 4310 24024
rect 4341 24021 4353 24024
rect 4387 24021 4399 24055
rect 4341 24015 4399 24021
rect 6822 24012 6828 24064
rect 6880 24052 6886 24064
rect 7024 24052 7052 24083
rect 9950 24080 9956 24132
rect 10008 24120 10014 24132
rect 10410 24120 10416 24132
rect 10008 24092 10416 24120
rect 10008 24080 10014 24092
rect 10410 24080 10416 24092
rect 10468 24120 10474 24132
rect 11057 24123 11115 24129
rect 11057 24120 11069 24123
rect 10468 24092 11069 24120
rect 10468 24080 10474 24092
rect 11057 24089 11069 24092
rect 11103 24089 11115 24123
rect 11057 24083 11115 24089
rect 11977 24123 12035 24129
rect 11977 24089 11989 24123
rect 12023 24120 12035 24123
rect 12526 24120 12532 24132
rect 12023 24092 12532 24120
rect 12023 24089 12035 24092
rect 11977 24083 12035 24089
rect 12526 24080 12532 24092
rect 12584 24080 12590 24132
rect 13906 24080 13912 24132
rect 13964 24120 13970 24132
rect 18248 24120 18276 24228
rect 18322 24216 18328 24268
rect 18380 24256 18386 24268
rect 18417 24259 18475 24265
rect 18417 24256 18429 24259
rect 18380 24228 18429 24256
rect 18380 24216 18386 24228
rect 18417 24225 18429 24228
rect 18463 24225 18475 24259
rect 18417 24219 18475 24225
rect 21729 24259 21787 24265
rect 21729 24225 21741 24259
rect 21775 24256 21787 24259
rect 22002 24256 22008 24268
rect 21775 24228 22008 24256
rect 21775 24225 21787 24228
rect 21729 24219 21787 24225
rect 22002 24216 22008 24228
rect 22060 24216 22066 24268
rect 18693 24191 18751 24197
rect 18693 24157 18705 24191
rect 18739 24188 18751 24191
rect 19058 24188 19064 24200
rect 18739 24160 19064 24188
rect 18739 24157 18751 24160
rect 18693 24151 18751 24157
rect 19058 24148 19064 24160
rect 19116 24148 19122 24200
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24188 19763 24191
rect 19794 24188 19800 24200
rect 19751 24160 19800 24188
rect 19751 24157 19763 24160
rect 19705 24151 19763 24157
rect 19794 24148 19800 24160
rect 19852 24148 19858 24200
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24188 20131 24191
rect 21818 24188 21824 24200
rect 20119 24160 21824 24188
rect 20119 24157 20131 24160
rect 20073 24151 20131 24157
rect 21818 24148 21824 24160
rect 21876 24188 21882 24200
rect 22738 24197 22744 24200
rect 21913 24191 21971 24197
rect 21913 24188 21925 24191
rect 21876 24160 21925 24188
rect 21876 24148 21882 24160
rect 21913 24157 21925 24160
rect 21959 24157 21971 24191
rect 22736 24188 22744 24197
rect 22699 24160 22744 24188
rect 21913 24151 21971 24157
rect 22736 24151 22744 24160
rect 22738 24148 22744 24151
rect 22796 24148 22802 24200
rect 22848 24197 22876 24296
rect 24857 24293 24869 24327
rect 24903 24324 24915 24327
rect 25406 24324 25412 24336
rect 24903 24296 25412 24324
rect 24903 24293 24915 24296
rect 24857 24287 24915 24293
rect 25406 24284 25412 24296
rect 25464 24284 25470 24336
rect 23566 24256 23572 24268
rect 23124 24228 23572 24256
rect 23124 24197 23152 24228
rect 23566 24216 23572 24228
rect 23624 24216 23630 24268
rect 24946 24216 24952 24268
rect 25004 24216 25010 24268
rect 25222 24256 25228 24268
rect 25135 24228 25228 24256
rect 25222 24216 25228 24228
rect 25280 24256 25286 24268
rect 26234 24256 26240 24268
rect 25280 24228 26240 24256
rect 25280 24216 25286 24228
rect 26234 24216 26240 24228
rect 26292 24216 26298 24268
rect 22833 24191 22891 24197
rect 22833 24157 22845 24191
rect 22879 24157 22891 24191
rect 22833 24151 22891 24157
rect 23108 24191 23166 24197
rect 23108 24157 23120 24191
rect 23154 24157 23166 24191
rect 23108 24151 23166 24157
rect 23198 24148 23204 24200
rect 23256 24188 23262 24200
rect 24964 24188 24992 24216
rect 25314 24188 25320 24200
rect 23256 24160 23301 24188
rect 24964 24160 25320 24188
rect 23256 24148 23262 24160
rect 25314 24148 25320 24160
rect 25372 24188 25378 24200
rect 25501 24191 25559 24197
rect 25501 24188 25513 24191
rect 25372 24160 25513 24188
rect 25372 24148 25378 24160
rect 25501 24157 25513 24160
rect 25547 24157 25559 24191
rect 25501 24151 25559 24157
rect 25590 24148 25596 24200
rect 25648 24188 25654 24200
rect 25961 24191 26019 24197
rect 25961 24188 25973 24191
rect 25648 24160 25973 24188
rect 25648 24148 25654 24160
rect 25961 24157 25973 24160
rect 26007 24157 26019 24191
rect 25961 24151 26019 24157
rect 26142 24148 26148 24200
rect 26200 24188 26206 24200
rect 26697 24191 26755 24197
rect 26697 24188 26709 24191
rect 26200 24160 26709 24188
rect 26200 24148 26206 24160
rect 26697 24157 26709 24160
rect 26743 24157 26755 24191
rect 26697 24151 26755 24157
rect 20898 24120 20904 24132
rect 13964 24092 14688 24120
rect 18248 24092 20904 24120
rect 13964 24080 13970 24092
rect 6880 24024 7052 24052
rect 6880 24012 6886 24024
rect 8202 24012 8208 24064
rect 8260 24052 8266 24064
rect 9401 24055 9459 24061
rect 9401 24052 9413 24055
rect 8260 24024 9413 24052
rect 8260 24012 8266 24024
rect 9401 24021 9413 24024
rect 9447 24052 9459 24055
rect 9582 24052 9588 24064
rect 9447 24024 9588 24052
rect 9447 24021 9459 24024
rect 9401 24015 9459 24021
rect 9582 24012 9588 24024
rect 9640 24012 9646 24064
rect 10597 24055 10655 24061
rect 10597 24021 10609 24055
rect 10643 24052 10655 24055
rect 10686 24052 10692 24064
rect 10643 24024 10692 24052
rect 10643 24021 10655 24024
rect 10597 24015 10655 24021
rect 10686 24012 10692 24024
rect 10744 24012 10750 24064
rect 14660 24061 14688 24092
rect 20898 24080 20904 24092
rect 20956 24120 20962 24132
rect 21085 24123 21143 24129
rect 21085 24120 21097 24123
rect 20956 24092 21097 24120
rect 20956 24080 20962 24092
rect 21085 24089 21097 24092
rect 21131 24089 21143 24123
rect 21085 24083 21143 24089
rect 22925 24123 22983 24129
rect 22925 24089 22937 24123
rect 22971 24089 22983 24123
rect 22925 24083 22983 24089
rect 14645 24055 14703 24061
rect 14645 24021 14657 24055
rect 14691 24052 14703 24055
rect 15010 24052 15016 24064
rect 14691 24024 15016 24052
rect 14691 24021 14703 24024
rect 14645 24015 14703 24021
rect 15010 24012 15016 24024
rect 15068 24012 15074 24064
rect 17218 24012 17224 24064
rect 17276 24052 17282 24064
rect 18417 24055 18475 24061
rect 18417 24052 18429 24055
rect 17276 24024 18429 24052
rect 17276 24012 17282 24024
rect 18417 24021 18429 24024
rect 18463 24021 18475 24055
rect 18417 24015 18475 24021
rect 19978 24012 19984 24064
rect 20036 24052 20042 24064
rect 20533 24055 20591 24061
rect 20533 24052 20545 24055
rect 20036 24024 20545 24052
rect 20036 24012 20042 24024
rect 20533 24021 20545 24024
rect 20579 24021 20591 24055
rect 20533 24015 20591 24021
rect 22094 24012 22100 24064
rect 22152 24052 22158 24064
rect 22940 24052 22968 24083
rect 24578 24080 24584 24132
rect 24636 24120 24642 24132
rect 24854 24120 24860 24132
rect 24636 24092 24860 24120
rect 24636 24080 24642 24092
rect 24854 24080 24860 24092
rect 24912 24120 24918 24132
rect 25016 24123 25074 24129
rect 25016 24120 25028 24123
rect 24912 24092 25028 24120
rect 24912 24080 24918 24092
rect 25016 24089 25028 24092
rect 25062 24089 25074 24123
rect 25016 24083 25074 24089
rect 25130 24080 25136 24132
rect 25188 24120 25194 24132
rect 25188 24092 26188 24120
rect 25188 24080 25194 24092
rect 26160 24061 26188 24092
rect 22152 24024 22968 24052
rect 26145 24055 26203 24061
rect 22152 24012 22158 24024
rect 26145 24021 26157 24055
rect 26191 24021 26203 24055
rect 26145 24015 26203 24021
rect 27341 24055 27399 24061
rect 27341 24021 27353 24055
rect 27387 24052 27399 24055
rect 27798 24052 27804 24064
rect 27387 24024 27804 24052
rect 27387 24021 27399 24024
rect 27341 24015 27399 24021
rect 27798 24012 27804 24024
rect 27856 24012 27862 24064
rect 28077 24055 28135 24061
rect 28077 24021 28089 24055
rect 28123 24052 28135 24055
rect 28534 24052 28540 24064
rect 28123 24024 28540 24052
rect 28123 24021 28135 24024
rect 28077 24015 28135 24021
rect 28534 24012 28540 24024
rect 28592 24012 28598 24064
rect 28718 24052 28724 24064
rect 28679 24024 28724 24052
rect 28718 24012 28724 24024
rect 28776 24012 28782 24064
rect 1104 23962 29600 23984
rect 1104 23910 8034 23962
rect 8086 23910 8098 23962
rect 8150 23910 8162 23962
rect 8214 23910 8226 23962
rect 8278 23910 8290 23962
rect 8342 23910 15118 23962
rect 15170 23910 15182 23962
rect 15234 23910 15246 23962
rect 15298 23910 15310 23962
rect 15362 23910 15374 23962
rect 15426 23910 22202 23962
rect 22254 23910 22266 23962
rect 22318 23910 22330 23962
rect 22382 23910 22394 23962
rect 22446 23910 22458 23962
rect 22510 23910 29286 23962
rect 29338 23910 29350 23962
rect 29402 23910 29414 23962
rect 29466 23910 29478 23962
rect 29530 23910 29542 23962
rect 29594 23910 29600 23962
rect 1104 23888 29600 23910
rect 4614 23848 4620 23860
rect 4575 23820 4620 23848
rect 4614 23808 4620 23820
rect 4672 23808 4678 23860
rect 6546 23808 6552 23860
rect 6604 23848 6610 23860
rect 6733 23851 6791 23857
rect 6733 23848 6745 23851
rect 6604 23820 6745 23848
rect 6604 23808 6610 23820
rect 6733 23817 6745 23820
rect 6779 23817 6791 23851
rect 9030 23848 9036 23860
rect 8991 23820 9036 23848
rect 6733 23811 6791 23817
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 10226 23848 10232 23860
rect 10187 23820 10232 23848
rect 10226 23808 10232 23820
rect 10284 23808 10290 23860
rect 10502 23808 10508 23860
rect 10560 23848 10566 23860
rect 12161 23851 12219 23857
rect 12161 23848 12173 23851
rect 10560 23820 12173 23848
rect 10560 23808 10566 23820
rect 12161 23817 12173 23820
rect 12207 23848 12219 23851
rect 14458 23848 14464 23860
rect 12207 23820 14464 23848
rect 12207 23817 12219 23820
rect 12161 23811 12219 23817
rect 14458 23808 14464 23820
rect 14516 23808 14522 23860
rect 14642 23848 14648 23860
rect 14603 23820 14648 23848
rect 14642 23808 14648 23820
rect 14700 23808 14706 23860
rect 18322 23808 18328 23860
rect 18380 23848 18386 23860
rect 18969 23851 19027 23857
rect 18969 23848 18981 23851
rect 18380 23820 18981 23848
rect 18380 23808 18386 23820
rect 18969 23817 18981 23820
rect 19015 23848 19027 23851
rect 19150 23848 19156 23860
rect 19015 23820 19156 23848
rect 19015 23817 19027 23820
rect 18969 23811 19027 23817
rect 19150 23808 19156 23820
rect 19208 23808 19214 23860
rect 19610 23808 19616 23860
rect 19668 23848 19674 23860
rect 19889 23851 19947 23857
rect 19889 23848 19901 23851
rect 19668 23820 19901 23848
rect 19668 23808 19674 23820
rect 19889 23817 19901 23820
rect 19935 23848 19947 23851
rect 20806 23848 20812 23860
rect 19935 23820 20812 23848
rect 19935 23817 19947 23820
rect 19889 23811 19947 23817
rect 20806 23808 20812 23820
rect 20864 23808 20870 23860
rect 21818 23848 21824 23860
rect 21779 23820 21824 23848
rect 21818 23808 21824 23820
rect 21876 23808 21882 23860
rect 22925 23851 22983 23857
rect 22925 23817 22937 23851
rect 22971 23848 22983 23851
rect 23198 23848 23204 23860
rect 22971 23820 23204 23848
rect 22971 23817 22983 23820
rect 22925 23811 22983 23817
rect 23198 23808 23204 23820
rect 23256 23808 23262 23860
rect 25222 23808 25228 23860
rect 25280 23808 25286 23860
rect 6365 23783 6423 23789
rect 6365 23780 6377 23783
rect 5184 23752 6377 23780
rect 5184 23721 5212 23752
rect 6365 23749 6377 23752
rect 6411 23749 6423 23783
rect 6365 23743 6423 23749
rect 7837 23783 7895 23789
rect 7837 23749 7849 23783
rect 7883 23780 7895 23783
rect 8110 23780 8116 23792
rect 7883 23752 8116 23780
rect 7883 23749 7895 23752
rect 7837 23743 7895 23749
rect 8110 23740 8116 23752
rect 8168 23780 8174 23792
rect 9306 23780 9312 23792
rect 8168 23752 9312 23780
rect 8168 23740 8174 23752
rect 9306 23740 9312 23752
rect 9364 23780 9370 23792
rect 9364 23752 9704 23780
rect 9364 23740 9370 23752
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23712 4767 23715
rect 5169 23715 5227 23721
rect 5169 23712 5181 23715
rect 4755 23684 5181 23712
rect 4755 23681 4767 23684
rect 4709 23675 4767 23681
rect 5169 23681 5181 23684
rect 5215 23681 5227 23715
rect 5169 23675 5227 23681
rect 5353 23715 5411 23721
rect 5353 23681 5365 23715
rect 5399 23712 5411 23715
rect 6178 23712 6184 23724
rect 5399 23684 6184 23712
rect 5399 23681 5411 23684
rect 5353 23675 5411 23681
rect 4249 23647 4307 23653
rect 4249 23613 4261 23647
rect 4295 23644 4307 23647
rect 5368 23644 5396 23675
rect 6178 23672 6184 23684
rect 6236 23672 6242 23724
rect 6454 23672 6460 23724
rect 6512 23712 6518 23724
rect 6549 23715 6607 23721
rect 6549 23712 6561 23715
rect 6512 23684 6561 23712
rect 6512 23672 6518 23684
rect 6549 23681 6561 23684
rect 6595 23681 6607 23715
rect 6822 23712 6828 23724
rect 6735 23684 6828 23712
rect 6549 23675 6607 23681
rect 6822 23672 6828 23684
rect 6880 23712 6886 23724
rect 7653 23715 7711 23721
rect 7653 23712 7665 23715
rect 6880 23684 7665 23712
rect 6880 23672 6886 23684
rect 7653 23681 7665 23684
rect 7699 23681 7711 23715
rect 7653 23675 7711 23681
rect 4295 23616 5396 23644
rect 4295 23613 4307 23616
rect 4249 23607 4307 23613
rect 6270 23604 6276 23656
rect 6328 23644 6334 23656
rect 6840 23644 6868 23672
rect 6328 23616 6868 23644
rect 7469 23647 7527 23653
rect 6328 23604 6334 23616
rect 7469 23613 7481 23647
rect 7515 23644 7527 23647
rect 7515 23616 7604 23644
rect 7515 23613 7527 23616
rect 7469 23607 7527 23613
rect 4338 23536 4344 23588
rect 4396 23576 4402 23588
rect 5261 23579 5319 23585
rect 5261 23576 5273 23579
rect 4396 23548 5273 23576
rect 4396 23536 4402 23548
rect 5261 23545 5273 23548
rect 5307 23545 5319 23579
rect 5261 23539 5319 23545
rect 3970 23468 3976 23520
rect 4028 23508 4034 23520
rect 4433 23511 4491 23517
rect 4433 23508 4445 23511
rect 4028 23480 4445 23508
rect 4028 23468 4034 23480
rect 4433 23477 4445 23480
rect 4479 23477 4491 23511
rect 7576 23508 7604 23616
rect 7668 23576 7696 23675
rect 8846 23672 8852 23724
rect 8904 23712 8910 23724
rect 8941 23715 8999 23721
rect 8941 23712 8953 23715
rect 8904 23684 8953 23712
rect 8904 23672 8910 23684
rect 8941 23681 8953 23684
rect 8987 23681 8999 23715
rect 8941 23675 8999 23681
rect 9125 23715 9183 23721
rect 9125 23681 9137 23715
rect 9171 23681 9183 23715
rect 9125 23675 9183 23681
rect 9140 23644 9168 23675
rect 9490 23672 9496 23724
rect 9548 23712 9554 23724
rect 9676 23721 9704 23752
rect 9585 23715 9643 23721
rect 9585 23712 9597 23715
rect 9548 23684 9597 23712
rect 9548 23672 9554 23684
rect 9585 23681 9597 23684
rect 9631 23681 9643 23715
rect 9676 23715 9736 23721
rect 9676 23684 9690 23715
rect 9585 23675 9643 23681
rect 9678 23681 9690 23684
rect 9724 23681 9736 23715
rect 9858 23712 9864 23724
rect 9819 23684 9864 23712
rect 9678 23675 9736 23681
rect 9858 23672 9864 23684
rect 9916 23672 9922 23724
rect 9953 23715 10011 23721
rect 9953 23681 9965 23715
rect 9999 23681 10011 23715
rect 9953 23675 10011 23681
rect 10091 23715 10149 23721
rect 10091 23681 10103 23715
rect 10137 23712 10149 23715
rect 10520 23712 10548 23808
rect 14829 23783 14887 23789
rect 14829 23749 14841 23783
rect 14875 23780 14887 23783
rect 15838 23780 15844 23792
rect 14875 23752 15844 23780
rect 14875 23749 14887 23752
rect 14829 23743 14887 23749
rect 15838 23740 15844 23752
rect 15896 23740 15902 23792
rect 21726 23780 21732 23792
rect 19168 23752 21732 23780
rect 10137 23684 10548 23712
rect 12989 23715 13047 23721
rect 10137 23681 10149 23684
rect 10091 23675 10149 23681
rect 12989 23681 13001 23715
rect 13035 23712 13047 23715
rect 13449 23715 13507 23721
rect 13449 23712 13461 23715
rect 13035 23684 13461 23712
rect 13035 23681 13047 23684
rect 12989 23675 13047 23681
rect 13449 23681 13461 23684
rect 13495 23681 13507 23715
rect 13449 23675 13507 23681
rect 9968 23644 9996 23675
rect 13538 23672 13544 23724
rect 13596 23712 13602 23724
rect 13633 23715 13691 23721
rect 13633 23712 13645 23715
rect 13596 23684 13645 23712
rect 13596 23672 13602 23684
rect 13633 23681 13645 23684
rect 13679 23681 13691 23715
rect 13633 23675 13691 23681
rect 13817 23715 13875 23721
rect 13817 23681 13829 23715
rect 13863 23712 13875 23715
rect 14366 23712 14372 23724
rect 13863 23684 14372 23712
rect 13863 23681 13875 23684
rect 13817 23675 13875 23681
rect 14366 23672 14372 23684
rect 14424 23672 14430 23724
rect 16945 23715 17003 23721
rect 16945 23681 16957 23715
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23681 17095 23715
rect 17037 23675 17095 23681
rect 17129 23715 17187 23721
rect 17129 23681 17141 23715
rect 17175 23712 17187 23715
rect 17218 23712 17224 23724
rect 17175 23684 17224 23712
rect 17175 23681 17187 23684
rect 17129 23675 17187 23681
rect 11609 23647 11667 23653
rect 11609 23644 11621 23647
rect 9048 23616 11621 23644
rect 8389 23579 8447 23585
rect 8389 23576 8401 23579
rect 7668 23548 8401 23576
rect 8389 23545 8401 23548
rect 8435 23576 8447 23579
rect 9048 23576 9076 23616
rect 11609 23613 11621 23616
rect 11655 23644 11667 23647
rect 12710 23644 12716 23656
rect 11655 23616 12716 23644
rect 11655 23613 11667 23616
rect 11609 23607 11667 23613
rect 12710 23604 12716 23616
rect 12768 23604 12774 23656
rect 16960 23644 16988 23675
rect 12820 23616 16988 23644
rect 12820 23585 12848 23616
rect 13464 23588 13492 23616
rect 17052 23588 17080 23675
rect 17218 23672 17224 23684
rect 17276 23672 17282 23724
rect 19168 23721 19196 23752
rect 21726 23740 21732 23752
rect 21784 23780 21790 23792
rect 22002 23780 22008 23792
rect 21784 23752 22008 23780
rect 21784 23740 21790 23752
rect 22002 23740 22008 23752
rect 22060 23740 22066 23792
rect 22094 23740 22100 23792
rect 22152 23780 22158 23792
rect 22465 23783 22523 23789
rect 22465 23780 22477 23783
rect 22152 23752 22477 23780
rect 22152 23740 22158 23752
rect 22465 23749 22477 23752
rect 22511 23780 22523 23783
rect 22554 23780 22560 23792
rect 22511 23752 22560 23780
rect 22511 23749 22523 23752
rect 22465 23743 22523 23749
rect 22554 23740 22560 23752
rect 22612 23740 22618 23792
rect 25240 23780 25268 23808
rect 24964 23752 25268 23780
rect 17313 23715 17371 23721
rect 17313 23681 17325 23715
rect 17359 23681 17371 23715
rect 17313 23675 17371 23681
rect 19153 23715 19211 23721
rect 19153 23681 19165 23715
rect 19199 23681 19211 23715
rect 19153 23675 19211 23681
rect 19337 23715 19395 23721
rect 19337 23681 19349 23715
rect 19383 23681 19395 23715
rect 19337 23675 19395 23681
rect 8435 23548 9076 23576
rect 12805 23579 12863 23585
rect 8435 23545 8447 23548
rect 8389 23539 8447 23545
rect 12805 23545 12817 23579
rect 12851 23545 12863 23579
rect 12805 23539 12863 23545
rect 13446 23536 13452 23588
rect 13504 23536 13510 23588
rect 14182 23536 14188 23588
rect 14240 23576 14246 23588
rect 15197 23579 15255 23585
rect 15197 23576 15209 23579
rect 14240 23548 15209 23576
rect 14240 23536 14246 23548
rect 15197 23545 15209 23548
rect 15243 23545 15255 23579
rect 15746 23576 15752 23588
rect 15659 23548 15752 23576
rect 15197 23539 15255 23545
rect 15746 23536 15752 23548
rect 15804 23576 15810 23588
rect 15804 23548 16896 23576
rect 15804 23536 15810 23548
rect 8846 23508 8852 23520
rect 7576 23480 8852 23508
rect 4433 23471 4491 23477
rect 8846 23468 8852 23480
rect 8904 23468 8910 23520
rect 10778 23508 10784 23520
rect 10739 23480 10784 23508
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 14826 23508 14832 23520
rect 14787 23480 14832 23508
rect 14826 23468 14832 23480
rect 14884 23468 14890 23520
rect 16669 23511 16727 23517
rect 16669 23477 16681 23511
rect 16715 23508 16727 23511
rect 16758 23508 16764 23520
rect 16715 23480 16764 23508
rect 16715 23477 16727 23480
rect 16669 23471 16727 23477
rect 16758 23468 16764 23480
rect 16816 23468 16822 23520
rect 16868 23508 16896 23548
rect 17034 23536 17040 23588
rect 17092 23536 17098 23588
rect 17328 23576 17356 23675
rect 19352 23644 19380 23675
rect 19426 23672 19432 23724
rect 19484 23712 19490 23724
rect 20993 23715 21051 23721
rect 20993 23712 21005 23715
rect 19484 23684 21005 23712
rect 19484 23672 19490 23684
rect 20993 23681 21005 23684
rect 21039 23712 21051 23715
rect 22922 23712 22928 23724
rect 21039 23684 22928 23712
rect 21039 23681 21051 23684
rect 20993 23675 21051 23681
rect 22922 23672 22928 23684
rect 22980 23672 22986 23724
rect 24964 23721 24992 23752
rect 24765 23715 24823 23721
rect 24765 23681 24777 23715
rect 24811 23681 24823 23715
rect 24765 23675 24823 23681
rect 24949 23715 25007 23721
rect 24949 23681 24961 23715
rect 24995 23681 25007 23715
rect 24949 23675 25007 23681
rect 25225 23715 25283 23721
rect 25225 23681 25237 23715
rect 25271 23712 25283 23715
rect 25314 23712 25320 23724
rect 25271 23684 25320 23712
rect 25271 23681 25283 23684
rect 25225 23675 25283 23681
rect 19794 23644 19800 23656
rect 19352 23616 19800 23644
rect 19794 23604 19800 23616
rect 19852 23644 19858 23656
rect 20349 23647 20407 23653
rect 20349 23644 20361 23647
rect 19852 23616 20361 23644
rect 19852 23604 19858 23616
rect 20349 23613 20361 23616
rect 20395 23613 20407 23647
rect 23934 23644 23940 23656
rect 20349 23607 20407 23613
rect 22756 23616 23940 23644
rect 20714 23576 20720 23588
rect 17328 23548 20720 23576
rect 20714 23536 20720 23548
rect 20772 23536 20778 23588
rect 22756 23585 22784 23616
rect 23934 23604 23940 23616
rect 23992 23604 23998 23656
rect 24780 23644 24808 23675
rect 25314 23672 25320 23684
rect 25372 23672 25378 23724
rect 25961 23715 26019 23721
rect 25961 23681 25973 23715
rect 26007 23712 26019 23715
rect 26142 23712 26148 23724
rect 26007 23684 26148 23712
rect 26007 23681 26019 23684
rect 25961 23675 26019 23681
rect 26142 23672 26148 23684
rect 26200 23672 26206 23724
rect 28258 23672 28264 23724
rect 28316 23712 28322 23724
rect 28445 23715 28503 23721
rect 28445 23712 28457 23715
rect 28316 23684 28457 23712
rect 28316 23672 28322 23684
rect 28445 23681 28457 23684
rect 28491 23681 28503 23715
rect 28445 23675 28503 23681
rect 24854 23644 24860 23656
rect 24767 23616 24860 23644
rect 24854 23604 24860 23616
rect 24912 23644 24918 23656
rect 25498 23644 25504 23656
rect 24912 23616 25504 23644
rect 24912 23604 24918 23616
rect 25498 23604 25504 23616
rect 25556 23644 25562 23656
rect 25556 23616 25820 23644
rect 25556 23604 25562 23616
rect 25792 23585 25820 23616
rect 22741 23579 22799 23585
rect 22741 23545 22753 23579
rect 22787 23545 22799 23579
rect 24581 23579 24639 23585
rect 24581 23576 24593 23579
rect 22741 23539 22799 23545
rect 22848 23548 24593 23576
rect 17494 23508 17500 23520
rect 16868 23480 17500 23508
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 19886 23508 19892 23520
rect 19392 23480 19892 23508
rect 19392 23468 19398 23480
rect 19886 23468 19892 23480
rect 19944 23468 19950 23520
rect 21174 23468 21180 23520
rect 21232 23508 21238 23520
rect 22848 23508 22876 23548
rect 24581 23545 24593 23548
rect 24627 23545 24639 23579
rect 24581 23539 24639 23545
rect 25777 23579 25835 23585
rect 25777 23545 25789 23579
rect 25823 23545 25835 23579
rect 25777 23539 25835 23545
rect 26878 23536 26884 23588
rect 26936 23576 26942 23588
rect 27801 23579 27859 23585
rect 27801 23576 27813 23579
rect 26936 23548 27813 23576
rect 26936 23536 26942 23548
rect 27801 23545 27813 23548
rect 27847 23545 27859 23579
rect 27801 23539 27859 23545
rect 21232 23480 22876 23508
rect 21232 23468 21238 23480
rect 22922 23468 22928 23520
rect 22980 23508 22986 23520
rect 23385 23511 23443 23517
rect 23385 23508 23397 23511
rect 22980 23480 23397 23508
rect 22980 23468 22986 23480
rect 23385 23477 23397 23480
rect 23431 23477 23443 23511
rect 25130 23508 25136 23520
rect 25091 23480 25136 23508
rect 23385 23471 23443 23477
rect 25130 23468 25136 23480
rect 25188 23468 25194 23520
rect 27065 23511 27123 23517
rect 27065 23477 27077 23511
rect 27111 23508 27123 23511
rect 27522 23508 27528 23520
rect 27111 23480 27528 23508
rect 27111 23477 27123 23480
rect 27065 23471 27123 23477
rect 27522 23468 27528 23480
rect 27580 23468 27586 23520
rect 28626 23508 28632 23520
rect 28587 23480 28632 23508
rect 28626 23468 28632 23480
rect 28684 23468 28690 23520
rect 1104 23418 29440 23440
rect 1104 23366 4492 23418
rect 4544 23366 4556 23418
rect 4608 23366 4620 23418
rect 4672 23366 4684 23418
rect 4736 23366 4748 23418
rect 4800 23366 11576 23418
rect 11628 23366 11640 23418
rect 11692 23366 11704 23418
rect 11756 23366 11768 23418
rect 11820 23366 11832 23418
rect 11884 23366 18660 23418
rect 18712 23366 18724 23418
rect 18776 23366 18788 23418
rect 18840 23366 18852 23418
rect 18904 23366 18916 23418
rect 18968 23366 25744 23418
rect 25796 23366 25808 23418
rect 25860 23366 25872 23418
rect 25924 23366 25936 23418
rect 25988 23366 26000 23418
rect 26052 23366 29440 23418
rect 1104 23344 29440 23366
rect 4338 23304 4344 23316
rect 4299 23276 4344 23304
rect 4338 23264 4344 23276
rect 4396 23264 4402 23316
rect 6178 23304 6184 23316
rect 6139 23276 6184 23304
rect 6178 23264 6184 23276
rect 6236 23264 6242 23316
rect 10962 23264 10968 23316
rect 11020 23304 11026 23316
rect 11333 23307 11391 23313
rect 11333 23304 11345 23307
rect 11020 23276 11345 23304
rect 11020 23264 11026 23276
rect 11333 23273 11345 23276
rect 11379 23273 11391 23307
rect 14182 23304 14188 23316
rect 11333 23267 11391 23273
rect 12268 23276 14188 23304
rect 7742 23128 7748 23180
rect 7800 23128 7806 23180
rect 10045 23171 10103 23177
rect 10045 23137 10057 23171
rect 10091 23168 10103 23171
rect 11057 23171 11115 23177
rect 10091 23140 10916 23168
rect 10091 23137 10103 23140
rect 10045 23131 10103 23137
rect 4154 23060 4160 23112
rect 4212 23100 4218 23112
rect 4249 23103 4307 23109
rect 4249 23100 4261 23103
rect 4212 23072 4261 23100
rect 4212 23060 4218 23072
rect 4249 23069 4261 23072
rect 4295 23069 4307 23103
rect 4249 23063 4307 23069
rect 4338 23060 4344 23112
rect 4396 23100 4402 23112
rect 4709 23103 4767 23109
rect 4396 23072 4441 23100
rect 4396 23060 4402 23072
rect 4709 23069 4721 23103
rect 4755 23100 4767 23103
rect 4982 23100 4988 23112
rect 4755 23072 4988 23100
rect 4755 23069 4767 23072
rect 4709 23063 4767 23069
rect 4982 23060 4988 23072
rect 5040 23060 5046 23112
rect 6181 23103 6239 23109
rect 6181 23069 6193 23103
rect 6227 23100 6239 23103
rect 6546 23100 6552 23112
rect 6227 23072 6552 23100
rect 6227 23069 6239 23072
rect 6181 23063 6239 23069
rect 6546 23060 6552 23072
rect 6604 23060 6610 23112
rect 7374 23060 7380 23112
rect 7432 23100 7438 23112
rect 7607 23103 7665 23109
rect 7607 23100 7619 23103
rect 7432 23072 7619 23100
rect 7432 23060 7438 23072
rect 7607 23069 7619 23072
rect 7653 23069 7665 23103
rect 7760 23100 7788 23128
rect 7965 23103 8023 23109
rect 7965 23100 7977 23103
rect 7760 23072 7977 23100
rect 7607 23063 7665 23069
rect 7965 23069 7977 23072
rect 8011 23069 8023 23103
rect 8110 23100 8116 23112
rect 8071 23072 8116 23100
rect 7965 23063 8023 23069
rect 8110 23060 8116 23072
rect 8168 23060 8174 23112
rect 9582 23060 9588 23112
rect 9640 23100 9646 23112
rect 9953 23103 10011 23109
rect 9953 23100 9965 23103
rect 9640 23072 9965 23100
rect 9640 23060 9646 23072
rect 9953 23069 9965 23072
rect 9999 23069 10011 23103
rect 9953 23063 10011 23069
rect 10173 23103 10231 23109
rect 10173 23069 10185 23103
rect 10219 23100 10231 23103
rect 10318 23100 10324 23112
rect 10219 23072 10324 23100
rect 10219 23069 10231 23072
rect 10173 23063 10231 23069
rect 10318 23060 10324 23072
rect 10376 23060 10382 23112
rect 10686 23100 10692 23112
rect 10647 23072 10692 23100
rect 10686 23060 10692 23072
rect 10744 23060 10750 23112
rect 10888 23109 10916 23140
rect 11057 23137 11069 23171
rect 11103 23168 11115 23171
rect 12161 23171 12219 23177
rect 12161 23168 12173 23171
rect 11103 23140 12173 23168
rect 11103 23137 11115 23140
rect 11057 23131 11115 23137
rect 12161 23137 12173 23140
rect 12207 23137 12219 23171
rect 12161 23131 12219 23137
rect 10873 23103 10931 23109
rect 10873 23069 10885 23103
rect 10919 23069 10931 23103
rect 10873 23063 10931 23069
rect 10965 23103 11023 23109
rect 10965 23069 10977 23103
rect 11011 23069 11023 23103
rect 10965 23063 11023 23069
rect 11149 23103 11207 23109
rect 11149 23069 11161 23103
rect 11195 23100 11207 23103
rect 12268 23100 12296 23276
rect 14182 23264 14188 23276
rect 14240 23264 14246 23316
rect 14366 23264 14372 23316
rect 14424 23304 14430 23316
rect 15838 23304 15844 23316
rect 14424 23276 15148 23304
rect 15799 23276 15844 23304
rect 14424 23264 14430 23276
rect 13170 23236 13176 23248
rect 12406 23208 13176 23236
rect 12406 23168 12434 23208
rect 13170 23196 13176 23208
rect 13228 23236 13234 23248
rect 15120 23236 15148 23276
rect 15838 23264 15844 23276
rect 15896 23264 15902 23316
rect 17034 23304 17040 23316
rect 16995 23276 17040 23304
rect 17034 23264 17040 23276
rect 17092 23264 17098 23316
rect 19150 23264 19156 23316
rect 19208 23304 19214 23316
rect 19208 23276 19840 23304
rect 19208 23264 19214 23276
rect 19334 23236 19340 23248
rect 13228 23208 15056 23236
rect 15120 23208 19340 23236
rect 13228 23196 13234 23208
rect 12360 23140 12434 23168
rect 12621 23171 12679 23177
rect 12360 23109 12388 23140
rect 12621 23137 12633 23171
rect 12667 23168 12679 23171
rect 13262 23168 13268 23180
rect 12667 23140 13268 23168
rect 12667 23137 12679 23140
rect 12621 23131 12679 23137
rect 13262 23128 13268 23140
rect 13320 23128 13326 23180
rect 15028 23112 15056 23208
rect 19334 23196 19340 23208
rect 19392 23196 19398 23248
rect 15102 23128 15108 23180
rect 15160 23168 15166 23180
rect 16393 23171 16451 23177
rect 16393 23168 16405 23171
rect 15160 23140 16405 23168
rect 15160 23128 15166 23140
rect 16393 23137 16405 23140
rect 16439 23168 16451 23171
rect 16942 23168 16948 23180
rect 16439 23140 16948 23168
rect 16439 23137 16451 23140
rect 16393 23131 16451 23137
rect 16942 23128 16948 23140
rect 17000 23128 17006 23180
rect 19245 23171 19303 23177
rect 19245 23168 19257 23171
rect 18432 23140 19257 23168
rect 11195 23072 12296 23100
rect 12345 23103 12403 23109
rect 11195 23069 11207 23072
rect 11149 23063 11207 23069
rect 12345 23069 12357 23103
rect 12391 23069 12403 23103
rect 12526 23100 12532 23112
rect 12487 23072 12532 23100
rect 12345 23063 12403 23069
rect 5721 23035 5779 23041
rect 5721 23001 5733 23035
rect 5767 23032 5779 23035
rect 6270 23032 6276 23044
rect 5767 23004 6276 23032
rect 5767 23001 5779 23004
rect 5721 22995 5779 23001
rect 6270 22992 6276 23004
rect 6328 22992 6334 23044
rect 6454 23032 6460 23044
rect 6415 23004 6460 23032
rect 6454 22992 6460 23004
rect 6512 22992 6518 23044
rect 7745 23035 7803 23041
rect 7745 23032 7757 23035
rect 7024 23004 7757 23032
rect 7024 22976 7052 23004
rect 7745 23001 7757 23004
rect 7791 23001 7803 23035
rect 7745 22995 7803 23001
rect 7837 23035 7895 23041
rect 7837 23001 7849 23035
rect 7883 23032 7895 23035
rect 9600 23032 9628 23060
rect 7883 23004 9628 23032
rect 9769 23035 9827 23041
rect 7883 23001 7895 23004
rect 7837 22995 7895 23001
rect 9769 23001 9781 23035
rect 9815 23001 9827 23035
rect 10042 23032 10048 23044
rect 9955 23004 10048 23032
rect 9769 22995 9827 23001
rect 1489 22967 1547 22973
rect 1489 22933 1501 22967
rect 1535 22964 1547 22967
rect 1578 22964 1584 22976
rect 1535 22936 1584 22964
rect 1535 22933 1547 22936
rect 1489 22927 1547 22933
rect 1578 22924 1584 22936
rect 1636 22924 1642 22976
rect 3786 22924 3792 22976
rect 3844 22964 3850 22976
rect 4065 22967 4123 22973
rect 4065 22964 4077 22967
rect 3844 22936 4077 22964
rect 3844 22924 3850 22936
rect 4065 22933 4077 22936
rect 4111 22933 4123 22967
rect 7006 22964 7012 22976
rect 6967 22936 7012 22964
rect 4065 22927 4123 22933
rect 7006 22924 7012 22936
rect 7064 22924 7070 22976
rect 7466 22964 7472 22976
rect 7427 22936 7472 22964
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 9309 22967 9367 22973
rect 9309 22933 9321 22967
rect 9355 22964 9367 22967
rect 9784 22964 9812 22995
rect 10042 22992 10048 23004
rect 10100 23032 10106 23044
rect 10778 23032 10784 23044
rect 10100 23004 10784 23032
rect 10100 22992 10106 23004
rect 10778 22992 10784 23004
rect 10836 22992 10842 23044
rect 10980 23032 11008 23063
rect 12526 23060 12532 23072
rect 12584 23060 12590 23112
rect 13357 23103 13415 23109
rect 13357 23069 13369 23103
rect 13403 23100 13415 23103
rect 13538 23100 13544 23112
rect 13403 23072 13544 23100
rect 13403 23069 13415 23072
rect 13357 23063 13415 23069
rect 13538 23060 13544 23072
rect 13596 23060 13602 23112
rect 14366 23100 14372 23112
rect 14327 23072 14372 23100
rect 14366 23060 14372 23072
rect 14424 23060 14430 23112
rect 15010 23060 15016 23112
rect 15068 23100 15074 23112
rect 15378 23109 15384 23112
rect 15197 23103 15255 23109
rect 15197 23100 15209 23103
rect 15068 23072 15209 23100
rect 15068 23060 15074 23072
rect 15197 23069 15209 23072
rect 15243 23069 15255 23103
rect 15197 23063 15255 23069
rect 15345 23103 15384 23109
rect 15345 23069 15357 23103
rect 15345 23063 15384 23069
rect 15378 23060 15384 23063
rect 15436 23060 15442 23112
rect 15703 23103 15761 23109
rect 15703 23069 15715 23103
rect 15749 23100 15761 23103
rect 16298 23100 16304 23112
rect 15749 23072 16304 23100
rect 15749 23069 15761 23072
rect 15703 23063 15761 23069
rect 16298 23060 16304 23072
rect 16356 23060 16362 23112
rect 16482 23060 16488 23112
rect 16540 23100 16546 23112
rect 18432 23109 18460 23140
rect 19245 23137 19257 23140
rect 19291 23137 19303 23171
rect 19245 23131 19303 23137
rect 16856 23103 16914 23109
rect 16856 23100 16868 23103
rect 16540 23072 16585 23100
rect 16684 23072 16868 23100
rect 16540 23060 16546 23072
rect 16684 23044 16712 23072
rect 16856 23069 16868 23072
rect 16902 23069 16914 23103
rect 16856 23063 16914 23069
rect 18417 23103 18475 23109
rect 18417 23069 18429 23103
rect 18463 23069 18475 23103
rect 18417 23063 18475 23069
rect 18693 23103 18751 23109
rect 18693 23069 18705 23103
rect 18739 23100 18751 23103
rect 18966 23100 18972 23112
rect 18739 23072 18972 23100
rect 18739 23069 18751 23072
rect 18693 23063 18751 23069
rect 18966 23060 18972 23072
rect 19024 23060 19030 23112
rect 19426 23060 19432 23112
rect 19484 23109 19490 23112
rect 19484 23103 19533 23109
rect 19484 23069 19487 23103
rect 19521 23069 19533 23103
rect 19484 23063 19533 23069
rect 19484 23060 19490 23063
rect 19591 23060 19597 23112
rect 19649 23109 19655 23112
rect 19649 23103 19668 23109
rect 19656 23069 19668 23103
rect 19649 23063 19668 23069
rect 19710 23103 19768 23109
rect 19710 23069 19722 23103
rect 19756 23100 19768 23103
rect 19812 23100 19840 23276
rect 19886 23264 19892 23316
rect 19944 23304 19950 23316
rect 20717 23307 20775 23313
rect 20717 23304 20729 23307
rect 19944 23276 20729 23304
rect 19944 23264 19950 23276
rect 20717 23273 20729 23276
rect 20763 23273 20775 23307
rect 20717 23267 20775 23273
rect 20806 23264 20812 23316
rect 20864 23304 20870 23316
rect 22738 23304 22744 23316
rect 20864 23276 22744 23304
rect 20864 23264 20870 23276
rect 22738 23264 22744 23276
rect 22796 23264 22802 23316
rect 21082 23128 21088 23180
rect 21140 23168 21146 23180
rect 24673 23171 24731 23177
rect 24673 23168 24685 23171
rect 21140 23140 24685 23168
rect 21140 23128 21146 23140
rect 24673 23137 24685 23140
rect 24719 23137 24731 23171
rect 24673 23131 24731 23137
rect 25222 23128 25228 23180
rect 25280 23168 25286 23180
rect 25501 23171 25559 23177
rect 25501 23168 25513 23171
rect 25280 23140 25513 23168
rect 25280 23128 25286 23140
rect 25501 23137 25513 23140
rect 25547 23137 25559 23171
rect 25501 23131 25559 23137
rect 26234 23128 26240 23180
rect 26292 23168 26298 23180
rect 26881 23171 26939 23177
rect 26881 23168 26893 23171
rect 26292 23140 26893 23168
rect 26292 23128 26298 23140
rect 26881 23137 26893 23140
rect 26927 23137 26939 23171
rect 26881 23131 26939 23137
rect 26970 23128 26976 23180
rect 27028 23168 27034 23180
rect 27525 23171 27583 23177
rect 27525 23168 27537 23171
rect 27028 23140 27537 23168
rect 27028 23128 27034 23140
rect 27525 23137 27537 23140
rect 27571 23137 27583 23171
rect 27798 23168 27804 23180
rect 27759 23140 27804 23168
rect 27525 23131 27583 23137
rect 27798 23128 27804 23140
rect 27856 23128 27862 23180
rect 28074 23168 28080 23180
rect 28035 23140 28080 23168
rect 28074 23128 28080 23140
rect 28132 23128 28138 23180
rect 28442 23128 28448 23180
rect 28500 23168 28506 23180
rect 28721 23171 28779 23177
rect 28721 23168 28733 23171
rect 28500 23140 28733 23168
rect 28500 23128 28506 23140
rect 28721 23137 28733 23140
rect 28767 23137 28779 23171
rect 28721 23131 28779 23137
rect 19756 23072 19840 23100
rect 19889 23103 19947 23109
rect 19756 23069 19768 23072
rect 19710 23063 19768 23069
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 19978 23100 19984 23112
rect 19935 23072 19984 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 19649 23060 19655 23063
rect 19978 23060 19984 23072
rect 20036 23060 20042 23112
rect 20898 23100 20904 23112
rect 20859 23072 20904 23100
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 21174 23100 21180 23112
rect 21135 23072 21180 23100
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 21818 23060 21824 23112
rect 21876 23100 21882 23112
rect 21913 23103 21971 23109
rect 21913 23100 21925 23103
rect 21876 23072 21925 23100
rect 21876 23060 21882 23072
rect 21913 23069 21925 23072
rect 21959 23069 21971 23103
rect 21913 23063 21971 23069
rect 14090 23032 14096 23044
rect 10980 23004 14096 23032
rect 14090 22992 14096 23004
rect 14148 22992 14154 23044
rect 15473 23035 15531 23041
rect 15473 23001 15485 23035
rect 15519 23001 15531 23035
rect 15473 22995 15531 23001
rect 15565 23035 15623 23041
rect 15565 23001 15577 23035
rect 15611 23032 15623 23035
rect 16666 23032 16672 23044
rect 15611 23004 16672 23032
rect 15611 23001 15623 23004
rect 15565 22995 15623 23001
rect 10410 22964 10416 22976
rect 9355 22936 10416 22964
rect 9355 22933 9367 22936
rect 9309 22927 9367 22933
rect 10410 22924 10416 22936
rect 10468 22924 10474 22976
rect 15488 22964 15516 22995
rect 16666 22992 16672 23004
rect 16724 22992 16730 23044
rect 20916 23032 20944 23060
rect 21266 23032 21272 23044
rect 20916 23004 21272 23032
rect 21266 22992 21272 23004
rect 21324 22992 21330 23044
rect 21928 23032 21956 23063
rect 24210 23060 24216 23112
rect 24268 23100 24274 23112
rect 24489 23103 24547 23109
rect 24489 23100 24501 23103
rect 24268 23072 24501 23100
rect 24268 23060 24274 23072
rect 24489 23069 24501 23072
rect 24535 23069 24547 23103
rect 24762 23100 24768 23112
rect 24723 23072 24768 23100
rect 24489 23063 24547 23069
rect 24762 23060 24768 23072
rect 24820 23060 24826 23112
rect 25133 23103 25191 23109
rect 25133 23069 25145 23103
rect 25179 23100 25191 23103
rect 25314 23100 25320 23112
rect 25179 23072 25320 23100
rect 25179 23069 25191 23072
rect 25133 23063 25191 23069
rect 25314 23060 25320 23072
rect 25372 23060 25378 23112
rect 27706 23109 27712 23112
rect 27684 23103 27712 23109
rect 27684 23069 27696 23103
rect 27684 23063 27712 23069
rect 27706 23060 27712 23063
rect 27764 23060 27770 23112
rect 28534 23100 28540 23112
rect 28495 23072 28540 23100
rect 28534 23060 28540 23072
rect 28592 23060 28598 23112
rect 23293 23035 23351 23041
rect 23293 23032 23305 23035
rect 21928 23004 23305 23032
rect 23293 23001 23305 23004
rect 23339 23001 23351 23035
rect 23293 22995 23351 23001
rect 15654 22964 15660 22976
rect 15488 22936 15660 22964
rect 15654 22924 15660 22936
rect 15712 22924 15718 22976
rect 16853 22967 16911 22973
rect 16853 22933 16865 22967
rect 16899 22964 16911 22967
rect 18233 22967 18291 22973
rect 18233 22964 18245 22967
rect 16899 22936 18245 22964
rect 16899 22933 16911 22936
rect 16853 22927 16911 22933
rect 18233 22933 18245 22936
rect 18279 22933 18291 22967
rect 18233 22927 18291 22933
rect 18601 22967 18659 22973
rect 18601 22933 18613 22967
rect 18647 22964 18659 22967
rect 19334 22964 19340 22976
rect 18647 22936 19340 22964
rect 18647 22933 18659 22936
rect 18601 22927 18659 22933
rect 19334 22924 19340 22936
rect 19392 22964 19398 22976
rect 19702 22964 19708 22976
rect 19392 22936 19708 22964
rect 19392 22924 19398 22936
rect 19702 22924 19708 22936
rect 19760 22924 19766 22976
rect 21082 22964 21088 22976
rect 21043 22936 21088 22964
rect 21082 22924 21088 22936
rect 21140 22924 21146 22976
rect 22002 22924 22008 22976
rect 22060 22964 22066 22976
rect 22189 22967 22247 22973
rect 22189 22964 22201 22967
rect 22060 22936 22201 22964
rect 22060 22924 22066 22936
rect 22189 22933 22201 22936
rect 22235 22933 22247 22967
rect 25958 22964 25964 22976
rect 25919 22936 25964 22964
rect 22189 22927 22247 22933
rect 25958 22924 25964 22936
rect 26016 22924 26022 22976
rect 1104 22874 29600 22896
rect 1104 22822 8034 22874
rect 8086 22822 8098 22874
rect 8150 22822 8162 22874
rect 8214 22822 8226 22874
rect 8278 22822 8290 22874
rect 8342 22822 15118 22874
rect 15170 22822 15182 22874
rect 15234 22822 15246 22874
rect 15298 22822 15310 22874
rect 15362 22822 15374 22874
rect 15426 22822 22202 22874
rect 22254 22822 22266 22874
rect 22318 22822 22330 22874
rect 22382 22822 22394 22874
rect 22446 22822 22458 22874
rect 22510 22822 29286 22874
rect 29338 22822 29350 22874
rect 29402 22822 29414 22874
rect 29466 22822 29478 22874
rect 29530 22822 29542 22874
rect 29594 22822 29600 22874
rect 1104 22800 29600 22822
rect 4157 22763 4215 22769
rect 4157 22729 4169 22763
rect 4203 22760 4215 22763
rect 4982 22760 4988 22772
rect 4203 22732 4988 22760
rect 4203 22729 4215 22732
rect 4157 22723 4215 22729
rect 4982 22720 4988 22732
rect 5040 22720 5046 22772
rect 6546 22720 6552 22772
rect 6604 22760 6610 22772
rect 6825 22763 6883 22769
rect 6825 22760 6837 22763
rect 6604 22732 6837 22760
rect 6604 22720 6610 22732
rect 6825 22729 6837 22732
rect 6871 22729 6883 22763
rect 9674 22760 9680 22772
rect 9587 22732 9680 22760
rect 6825 22723 6883 22729
rect 9674 22720 9680 22732
rect 9732 22760 9738 22772
rect 10229 22763 10287 22769
rect 10229 22760 10241 22763
rect 9732 22732 10241 22760
rect 9732 22720 9738 22732
rect 10229 22729 10241 22732
rect 10275 22760 10287 22763
rect 10318 22760 10324 22772
rect 10275 22732 10324 22760
rect 10275 22729 10287 22732
rect 10229 22723 10287 22729
rect 10318 22720 10324 22732
rect 10376 22720 10382 22772
rect 10410 22720 10416 22772
rect 10468 22760 10474 22772
rect 12069 22763 12127 22769
rect 12069 22760 12081 22763
rect 10468 22732 12081 22760
rect 10468 22720 10474 22732
rect 12069 22729 12081 22732
rect 12115 22729 12127 22763
rect 12986 22760 12992 22772
rect 12947 22732 12992 22760
rect 12069 22723 12127 22729
rect 12986 22720 12992 22732
rect 13044 22720 13050 22772
rect 14826 22720 14832 22772
rect 14884 22760 14890 22772
rect 15013 22763 15071 22769
rect 15013 22760 15025 22763
rect 14884 22732 15025 22760
rect 14884 22720 14890 22732
rect 15013 22729 15025 22732
rect 15059 22729 15071 22763
rect 16666 22760 16672 22772
rect 16627 22732 16672 22760
rect 15013 22723 15071 22729
rect 16666 22720 16672 22732
rect 16724 22720 16730 22772
rect 18138 22720 18144 22772
rect 18196 22760 18202 22772
rect 18322 22760 18328 22772
rect 18196 22732 18328 22760
rect 18196 22720 18202 22732
rect 18322 22720 18328 22732
rect 18380 22760 18386 22772
rect 18693 22763 18751 22769
rect 18693 22760 18705 22763
rect 18380 22732 18705 22760
rect 18380 22720 18386 22732
rect 18693 22729 18705 22732
rect 18739 22729 18751 22763
rect 18693 22723 18751 22729
rect 19334 22720 19340 22772
rect 19392 22760 19398 22772
rect 19392 22732 19437 22760
rect 19392 22720 19398 22732
rect 20806 22720 20812 22772
rect 20864 22760 20870 22772
rect 21177 22763 21235 22769
rect 21177 22760 21189 22763
rect 20864 22732 21189 22760
rect 20864 22720 20870 22732
rect 21177 22729 21189 22732
rect 21223 22729 21235 22763
rect 21177 22723 21235 22729
rect 24762 22720 24768 22772
rect 24820 22760 24826 22772
rect 25317 22763 25375 22769
rect 25317 22760 25329 22763
rect 24820 22732 25329 22760
rect 24820 22720 24826 22732
rect 25317 22729 25329 22732
rect 25363 22760 25375 22763
rect 25958 22760 25964 22772
rect 25363 22732 25964 22760
rect 25363 22729 25375 22732
rect 25317 22723 25375 22729
rect 25958 22720 25964 22732
rect 26016 22760 26022 22772
rect 26053 22763 26111 22769
rect 26053 22760 26065 22763
rect 26016 22732 26065 22760
rect 26016 22720 26022 22732
rect 26053 22729 26065 22732
rect 26099 22729 26111 22763
rect 26053 22723 26111 22729
rect 3326 22692 3332 22704
rect 3287 22664 3332 22692
rect 3326 22652 3332 22664
rect 3384 22652 3390 22704
rect 6454 22652 6460 22704
rect 6512 22692 6518 22704
rect 7469 22695 7527 22701
rect 7469 22692 7481 22695
rect 6512 22664 7481 22692
rect 6512 22652 6518 22664
rect 7469 22661 7481 22664
rect 7515 22661 7527 22695
rect 8846 22692 8852 22704
rect 8759 22664 8852 22692
rect 7469 22655 7527 22661
rect 8846 22652 8852 22664
rect 8904 22692 8910 22704
rect 10042 22692 10048 22704
rect 8904 22664 10048 22692
rect 8904 22652 8910 22664
rect 10042 22652 10048 22664
rect 10100 22652 10106 22704
rect 11974 22692 11980 22704
rect 11935 22664 11980 22692
rect 11974 22652 11980 22664
rect 12032 22652 12038 22704
rect 13538 22692 13544 22704
rect 13004 22664 13544 22692
rect 1578 22624 1584 22636
rect 1539 22596 1584 22624
rect 1578 22584 1584 22596
rect 1636 22584 1642 22636
rect 2222 22584 2228 22636
rect 2280 22624 2286 22636
rect 2501 22627 2559 22633
rect 2501 22624 2513 22627
rect 2280 22596 2513 22624
rect 2280 22584 2286 22596
rect 2501 22593 2513 22596
rect 2547 22593 2559 22627
rect 2501 22587 2559 22593
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 3050 22624 3056 22636
rect 3007 22596 3056 22624
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 3050 22584 3056 22596
rect 3108 22584 3114 22636
rect 3970 22624 3976 22636
rect 3931 22596 3976 22624
rect 3970 22584 3976 22596
rect 4028 22584 4034 22636
rect 4246 22584 4252 22636
rect 4304 22624 4310 22636
rect 6917 22627 6975 22633
rect 4304 22596 4349 22624
rect 4304 22584 4310 22596
rect 6917 22593 6929 22627
rect 6963 22593 6975 22627
rect 6917 22587 6975 22593
rect 1762 22488 1768 22500
rect 1723 22460 1768 22488
rect 1762 22448 1768 22460
rect 1820 22448 1826 22500
rect 6932 22488 6960 22587
rect 7282 22584 7288 22636
rect 7340 22624 7346 22636
rect 7377 22627 7435 22633
rect 7377 22624 7389 22627
rect 7340 22596 7389 22624
rect 7340 22584 7346 22596
rect 7377 22593 7389 22596
rect 7423 22593 7435 22627
rect 7558 22624 7564 22636
rect 7519 22596 7564 22624
rect 7377 22587 7435 22593
rect 7558 22584 7564 22596
rect 7616 22584 7622 22636
rect 13004 22633 13032 22664
rect 13538 22652 13544 22664
rect 13596 22692 13602 22704
rect 13633 22695 13691 22701
rect 13633 22692 13645 22695
rect 13596 22664 13645 22692
rect 13596 22652 13602 22664
rect 13633 22661 13645 22664
rect 13679 22692 13691 22695
rect 14185 22695 14243 22701
rect 14185 22692 14197 22695
rect 13679 22664 14197 22692
rect 13679 22661 13691 22664
rect 13633 22655 13691 22661
rect 14185 22661 14197 22664
rect 14231 22692 14243 22695
rect 15746 22692 15752 22704
rect 14231 22664 15752 22692
rect 14231 22661 14243 22664
rect 14185 22655 14243 22661
rect 15746 22652 15752 22664
rect 15804 22652 15810 22704
rect 19352 22692 19380 22720
rect 21082 22692 21088 22704
rect 19352 22664 21088 22692
rect 21082 22652 21088 22664
rect 21140 22652 21146 22704
rect 23106 22692 23112 22704
rect 22664 22664 23112 22692
rect 12989 22627 13047 22633
rect 12989 22593 13001 22627
rect 13035 22593 13047 22627
rect 15010 22624 15016 22636
rect 14971 22596 15016 22624
rect 12989 22587 13047 22593
rect 15010 22584 15016 22596
rect 15068 22584 15074 22636
rect 15197 22627 15255 22633
rect 15197 22593 15209 22627
rect 15243 22593 15255 22627
rect 16850 22624 16856 22636
rect 16811 22596 16856 22624
rect 15197 22587 15255 22593
rect 8846 22488 8852 22500
rect 6932 22460 8852 22488
rect 8846 22448 8852 22460
rect 8904 22448 8910 22500
rect 15212 22488 15240 22587
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 16942 22584 16948 22636
rect 17000 22624 17006 22636
rect 17865 22627 17923 22633
rect 17000 22596 17045 22624
rect 17000 22584 17006 22596
rect 17865 22593 17877 22627
rect 17911 22624 17923 22627
rect 19242 22624 19248 22636
rect 17911 22596 19248 22624
rect 17911 22593 17923 22596
rect 17865 22587 17923 22593
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 21542 22584 21548 22636
rect 21600 22624 21606 22636
rect 21818 22624 21824 22636
rect 21600 22596 21824 22624
rect 21600 22584 21606 22596
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 22554 22624 22560 22636
rect 22515 22596 22560 22624
rect 22554 22584 22560 22596
rect 22612 22584 22618 22636
rect 22664 22633 22692 22664
rect 23106 22652 23112 22664
rect 23164 22652 23170 22704
rect 24210 22652 24216 22704
rect 24268 22692 24274 22704
rect 25434 22695 25492 22701
rect 25434 22692 25446 22695
rect 24268 22664 25446 22692
rect 24268 22652 24274 22664
rect 25434 22661 25446 22664
rect 25480 22692 25492 22695
rect 26973 22695 27031 22701
rect 26973 22692 26985 22695
rect 25480 22664 26985 22692
rect 25480 22661 25492 22664
rect 25434 22655 25492 22661
rect 26973 22661 26985 22664
rect 27019 22661 27031 22695
rect 26973 22655 27031 22661
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22593 22707 22627
rect 22830 22624 22836 22636
rect 22791 22596 22836 22624
rect 22649 22587 22707 22593
rect 22830 22584 22836 22596
rect 22888 22584 22894 22636
rect 22925 22627 22983 22633
rect 22925 22593 22937 22627
rect 22971 22624 22983 22627
rect 23569 22627 23627 22633
rect 23569 22624 23581 22627
rect 22971 22596 23581 22624
rect 22971 22593 22983 22596
rect 22925 22587 22983 22593
rect 23569 22593 23581 22596
rect 23615 22593 23627 22627
rect 23569 22587 23627 22593
rect 24949 22627 25007 22633
rect 24949 22593 24961 22627
rect 24995 22624 25007 22627
rect 25130 22624 25136 22636
rect 24995 22596 25136 22624
rect 24995 22593 25007 22596
rect 24949 22587 25007 22593
rect 16390 22516 16396 22568
rect 16448 22556 16454 22568
rect 22097 22559 22155 22565
rect 16448 22528 19656 22556
rect 16448 22516 16454 22528
rect 19628 22500 19656 22528
rect 22097 22525 22109 22559
rect 22143 22556 22155 22559
rect 22848 22556 22876 22584
rect 22143 22528 22876 22556
rect 22143 22525 22155 22528
rect 22097 22519 22155 22525
rect 17862 22488 17868 22500
rect 15212 22460 17868 22488
rect 17862 22448 17868 22460
rect 17920 22448 17926 22500
rect 19610 22448 19616 22500
rect 19668 22488 19674 22500
rect 20717 22491 20775 22497
rect 20717 22488 20729 22491
rect 19668 22460 20729 22488
rect 19668 22448 19674 22460
rect 20717 22457 20729 22460
rect 20763 22488 20775 22491
rect 21910 22488 21916 22500
rect 20763 22460 21916 22488
rect 20763 22457 20775 22460
rect 20717 22451 20775 22457
rect 21910 22448 21916 22460
rect 21968 22448 21974 22500
rect 22738 22448 22744 22500
rect 22796 22488 22802 22500
rect 22940 22488 22968 22587
rect 25130 22584 25136 22596
rect 25188 22584 25194 22636
rect 27985 22627 28043 22633
rect 27985 22593 27997 22627
rect 28031 22624 28043 22627
rect 28074 22624 28080 22636
rect 28031 22596 28080 22624
rect 28031 22593 28043 22596
rect 27985 22587 28043 22593
rect 28074 22584 28080 22596
rect 28132 22584 28138 22636
rect 25225 22559 25283 22565
rect 25225 22525 25237 22559
rect 25271 22556 25283 22559
rect 25314 22556 25320 22568
rect 25271 22528 25320 22556
rect 25271 22525 25283 22528
rect 25225 22519 25283 22525
rect 25314 22516 25320 22528
rect 25372 22516 25378 22568
rect 22796 22460 22968 22488
rect 22796 22448 22802 22460
rect 24026 22448 24032 22500
rect 24084 22488 24090 22500
rect 24121 22491 24179 22497
rect 24121 22488 24133 22491
rect 24084 22460 24133 22488
rect 24084 22448 24090 22460
rect 24121 22457 24133 22460
rect 24167 22457 24179 22491
rect 24121 22451 24179 22457
rect 3510 22380 3516 22432
rect 3568 22420 3574 22432
rect 3789 22423 3847 22429
rect 3789 22420 3801 22423
rect 3568 22392 3801 22420
rect 3568 22380 3574 22392
rect 3789 22389 3801 22392
rect 3835 22389 3847 22423
rect 8202 22420 8208 22432
rect 8163 22392 8208 22420
rect 3789 22383 3847 22389
rect 8202 22380 8208 22392
rect 8260 22380 8266 22432
rect 9950 22380 9956 22432
rect 10008 22420 10014 22432
rect 10689 22423 10747 22429
rect 10689 22420 10701 22423
rect 10008 22392 10701 22420
rect 10008 22380 10014 22392
rect 10689 22389 10701 22392
rect 10735 22389 10747 22423
rect 10689 22383 10747 22389
rect 19886 22380 19892 22432
rect 19944 22420 19950 22432
rect 20073 22423 20131 22429
rect 20073 22420 20085 22423
rect 19944 22392 20085 22420
rect 19944 22380 19950 22392
rect 20073 22389 20085 22392
rect 20119 22389 20131 22423
rect 20073 22383 20131 22389
rect 23109 22423 23167 22429
rect 23109 22389 23121 22423
rect 23155 22420 23167 22423
rect 23382 22420 23388 22432
rect 23155 22392 23388 22420
rect 23155 22389 23167 22392
rect 23109 22383 23167 22389
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 25590 22420 25596 22432
rect 25551 22392 25596 22420
rect 25590 22380 25596 22392
rect 25648 22380 25654 22432
rect 27890 22380 27896 22432
rect 27948 22420 27954 22432
rect 28077 22423 28135 22429
rect 28077 22420 28089 22423
rect 27948 22392 28089 22420
rect 27948 22380 27954 22392
rect 28077 22389 28089 22392
rect 28123 22389 28135 22423
rect 28077 22383 28135 22389
rect 1104 22330 29440 22352
rect 1104 22278 4492 22330
rect 4544 22278 4556 22330
rect 4608 22278 4620 22330
rect 4672 22278 4684 22330
rect 4736 22278 4748 22330
rect 4800 22278 11576 22330
rect 11628 22278 11640 22330
rect 11692 22278 11704 22330
rect 11756 22278 11768 22330
rect 11820 22278 11832 22330
rect 11884 22278 18660 22330
rect 18712 22278 18724 22330
rect 18776 22278 18788 22330
rect 18840 22278 18852 22330
rect 18904 22278 18916 22330
rect 18968 22278 25744 22330
rect 25796 22278 25808 22330
rect 25860 22278 25872 22330
rect 25924 22278 25936 22330
rect 25988 22278 26000 22330
rect 26052 22278 29440 22330
rect 1104 22256 29440 22278
rect 2222 22216 2228 22228
rect 2183 22188 2228 22216
rect 2222 22176 2228 22188
rect 2280 22176 2286 22228
rect 11241 22219 11299 22225
rect 11241 22185 11253 22219
rect 11287 22216 11299 22219
rect 11974 22216 11980 22228
rect 11287 22188 11980 22216
rect 11287 22185 11299 22188
rect 11241 22179 11299 22185
rect 7377 22151 7435 22157
rect 7377 22117 7389 22151
rect 7423 22148 7435 22151
rect 7558 22148 7564 22160
rect 7423 22120 7564 22148
rect 7423 22117 7435 22120
rect 7377 22111 7435 22117
rect 7558 22108 7564 22120
rect 7616 22148 7622 22160
rect 7616 22120 9536 22148
rect 7616 22108 7622 22120
rect 9508 22094 9536 22120
rect 2041 22083 2099 22089
rect 2041 22049 2053 22083
rect 2087 22080 2099 22083
rect 2958 22080 2964 22092
rect 2087 22052 2964 22080
rect 2087 22049 2099 22052
rect 2041 22043 2099 22049
rect 2958 22040 2964 22052
rect 3016 22040 3022 22092
rect 6825 22083 6883 22089
rect 6825 22049 6837 22083
rect 6871 22080 6883 22083
rect 7006 22080 7012 22092
rect 6871 22052 7012 22080
rect 6871 22049 6883 22052
rect 6825 22043 6883 22049
rect 7006 22040 7012 22052
rect 7064 22080 7070 22092
rect 9508 22089 9573 22094
rect 9493 22083 9573 22089
rect 7064 22052 7512 22080
rect 7064 22040 7070 22052
rect 1670 21972 1676 22024
rect 1728 22012 1734 22024
rect 1949 22015 2007 22021
rect 1949 22012 1961 22015
rect 1728 21984 1961 22012
rect 1728 21972 1734 21984
rect 1949 21981 1961 21984
rect 1995 22012 2007 22015
rect 2777 22015 2835 22021
rect 2777 22012 2789 22015
rect 1995 21984 2789 22012
rect 1995 21981 2007 21984
rect 1949 21975 2007 21981
rect 2777 21981 2789 21984
rect 2823 21981 2835 22015
rect 3970 22012 3976 22024
rect 3931 21984 3976 22012
rect 2777 21975 2835 21981
rect 3970 21972 3976 21984
rect 4028 21972 4034 22024
rect 6546 21972 6552 22024
rect 6604 22012 6610 22024
rect 7484 22021 7512 22052
rect 9493 22049 9505 22083
rect 9539 22066 9573 22083
rect 9677 22083 9735 22089
rect 9539 22049 9551 22066
rect 9493 22043 9551 22049
rect 9677 22049 9689 22083
rect 9723 22080 9735 22083
rect 11256 22080 11284 22179
rect 11974 22176 11980 22188
rect 12032 22216 12038 22228
rect 12437 22219 12495 22225
rect 12437 22216 12449 22219
rect 12032 22188 12449 22216
rect 12032 22176 12038 22188
rect 12437 22185 12449 22188
rect 12483 22185 12495 22219
rect 19058 22216 19064 22228
rect 12437 22179 12495 22185
rect 18064 22188 19064 22216
rect 9723 22052 11284 22080
rect 9723 22049 9735 22052
rect 9677 22043 9735 22049
rect 9876 22024 9904 22052
rect 13170 22040 13176 22092
rect 13228 22080 13234 22092
rect 14918 22080 14924 22092
rect 13228 22052 14688 22080
rect 14879 22052 14924 22080
rect 13228 22040 13234 22052
rect 7285 22015 7343 22021
rect 7285 22012 7297 22015
rect 6604 21984 7297 22012
rect 6604 21972 6610 21984
rect 7285 21981 7297 21984
rect 7331 21981 7343 22015
rect 7285 21975 7343 21981
rect 7469 22015 7527 22021
rect 7469 21981 7481 22015
rect 7515 22012 7527 22015
rect 7834 22012 7840 22024
rect 7515 21984 7840 22012
rect 7515 21981 7527 21984
rect 7469 21975 7527 21981
rect 7300 21944 7328 21975
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 9858 21972 9864 22024
rect 9916 21972 9922 22024
rect 14182 21972 14188 22024
rect 14240 22012 14246 22024
rect 14369 22015 14427 22021
rect 14369 22012 14381 22015
rect 14240 21984 14381 22012
rect 14240 21972 14246 21984
rect 14369 21981 14381 21984
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 7374 21944 7380 21956
rect 7287 21916 7380 21944
rect 7374 21904 7380 21916
rect 7432 21944 7438 21956
rect 7929 21947 7987 21953
rect 7929 21944 7941 21947
rect 7432 21916 7941 21944
rect 7432 21904 7438 21916
rect 7929 21913 7941 21916
rect 7975 21944 7987 21947
rect 8202 21944 8208 21956
rect 7975 21916 8208 21944
rect 7975 21913 7987 21916
rect 7929 21907 7987 21913
rect 8202 21904 8208 21916
rect 8260 21944 8266 21956
rect 8662 21944 8668 21956
rect 8260 21916 8668 21944
rect 8260 21904 8266 21916
rect 8662 21904 8668 21916
rect 8720 21904 8726 21956
rect 9398 21904 9404 21956
rect 9456 21944 9462 21956
rect 10594 21944 10600 21956
rect 9456 21916 10600 21944
rect 9456 21904 9462 21916
rect 10594 21904 10600 21916
rect 10652 21904 10658 21956
rect 14384 21944 14412 21975
rect 14458 21972 14464 22024
rect 14516 22012 14522 22024
rect 14660 22021 14688 22052
rect 14918 22040 14924 22052
rect 14976 22040 14982 22092
rect 14645 22015 14703 22021
rect 14516 21984 14561 22012
rect 14516 21972 14522 21984
rect 14645 21981 14657 22015
rect 14691 21981 14703 22015
rect 14645 21975 14703 21981
rect 14734 21972 14740 22024
rect 14792 22012 14798 22024
rect 18064 22012 18092 22188
rect 19058 22176 19064 22188
rect 19116 22216 19122 22228
rect 19245 22219 19303 22225
rect 19245 22216 19257 22219
rect 19116 22188 19257 22216
rect 19116 22176 19122 22188
rect 19245 22185 19257 22188
rect 19291 22185 19303 22219
rect 19245 22179 19303 22185
rect 22002 22176 22008 22228
rect 22060 22216 22066 22228
rect 22060 22188 22140 22216
rect 22060 22176 22066 22188
rect 21818 22148 21824 22160
rect 21744 22120 21824 22148
rect 19242 22080 19248 22092
rect 18524 22052 19248 22080
rect 18125 22015 18183 22021
rect 18125 22012 18137 22015
rect 14792 21984 14837 22012
rect 18064 21984 18137 22012
rect 14792 21972 14798 21984
rect 18125 21981 18137 21984
rect 18171 21981 18183 22015
rect 18322 22012 18328 22024
rect 18283 21984 18328 22012
rect 18125 21975 18183 21981
rect 18322 21972 18328 21984
rect 18380 21972 18386 22024
rect 18524 22021 18552 22052
rect 19242 22040 19248 22052
rect 19300 22040 19306 22092
rect 19886 22080 19892 22092
rect 19847 22052 19892 22080
rect 19886 22040 19892 22052
rect 19944 22040 19950 22092
rect 21358 22089 21364 22092
rect 21336 22083 21364 22089
rect 21336 22049 21348 22083
rect 21336 22043 21364 22049
rect 21358 22040 21364 22043
rect 21416 22040 21422 22092
rect 21453 22083 21511 22089
rect 21453 22049 21465 22083
rect 21499 22080 21511 22083
rect 21634 22080 21640 22092
rect 21499 22052 21640 22080
rect 21499 22049 21511 22052
rect 21453 22043 21511 22049
rect 21634 22040 21640 22052
rect 21692 22040 21698 22092
rect 21744 22089 21772 22120
rect 21818 22108 21824 22120
rect 21876 22148 21882 22160
rect 22112 22148 22140 22188
rect 23032 22188 28120 22216
rect 23032 22148 23060 22188
rect 21876 22120 23060 22148
rect 21876 22108 21882 22120
rect 21729 22083 21787 22089
rect 21729 22049 21741 22083
rect 21775 22080 21787 22083
rect 21775 22052 21809 22080
rect 21775 22049 21787 22052
rect 21729 22043 21787 22049
rect 22002 22040 22008 22092
rect 22060 22080 22066 22092
rect 23032 22089 23060 22120
rect 28092 22092 28120 22188
rect 23017 22083 23075 22089
rect 22060 22052 22416 22080
rect 22060 22040 22066 22052
rect 18509 22015 18567 22021
rect 18509 21981 18521 22015
rect 18555 21981 18567 22015
rect 18509 21975 18567 21981
rect 18601 22015 18659 22021
rect 18601 21981 18613 22015
rect 18647 22012 18659 22015
rect 18966 22012 18972 22024
rect 18647 21984 18972 22012
rect 18647 21981 18659 21984
rect 18601 21975 18659 21981
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 19610 22012 19616 22024
rect 19571 21984 19616 22012
rect 19610 21972 19616 21984
rect 19668 21972 19674 22024
rect 21174 21972 21180 22024
rect 21232 22012 21238 22024
rect 22388 22021 22416 22052
rect 23017 22049 23029 22083
rect 23063 22080 23075 22083
rect 24489 22083 24547 22089
rect 24489 22080 24501 22083
rect 23063 22052 23097 22080
rect 23216 22052 24501 22080
rect 23063 22049 23075 22052
rect 23017 22043 23075 22049
rect 23216 22021 23244 22052
rect 24489 22049 24501 22052
rect 24535 22080 24547 22083
rect 26145 22083 26203 22089
rect 26145 22080 26157 22083
rect 24535 22052 26157 22080
rect 24535 22049 24547 22052
rect 24489 22043 24547 22049
rect 26145 22049 26157 22052
rect 26191 22080 26203 22083
rect 26786 22080 26792 22092
rect 26191 22052 26792 22080
rect 26191 22049 26203 22052
rect 26145 22043 26203 22049
rect 26786 22040 26792 22052
rect 26844 22040 26850 22092
rect 28074 22080 28080 22092
rect 28035 22052 28080 22080
rect 28074 22040 28080 22052
rect 28132 22080 28138 22092
rect 28132 22052 28157 22080
rect 28132 22040 28138 22052
rect 22189 22015 22247 22021
rect 21232 21984 21277 22012
rect 21232 21972 21238 21984
rect 22189 21981 22201 22015
rect 22235 21981 22247 22015
rect 22189 21975 22247 21981
rect 22373 22015 22431 22021
rect 22373 21981 22385 22015
rect 22419 22012 22431 22015
rect 23201 22015 23259 22021
rect 23201 22012 23213 22015
rect 22419 21984 23213 22012
rect 22419 21981 22431 21984
rect 22373 21975 22431 21981
rect 23201 21981 23213 21984
rect 23247 21981 23259 22015
rect 23201 21975 23259 21981
rect 25501 22015 25559 22021
rect 25501 21981 25513 22015
rect 25547 22012 25559 22015
rect 25590 22012 25596 22024
rect 25547 21984 25596 22012
rect 25547 21981 25559 21984
rect 25501 21975 25559 21981
rect 14550 21944 14556 21956
rect 14384 21916 14556 21944
rect 14550 21904 14556 21916
rect 14608 21904 14614 21956
rect 16850 21904 16856 21956
rect 16908 21944 16914 21956
rect 18233 21947 18291 21953
rect 18233 21944 18245 21947
rect 16908 21916 18245 21944
rect 16908 21904 16914 21916
rect 18233 21913 18245 21916
rect 18279 21913 18291 21947
rect 18233 21907 18291 21913
rect 19150 21904 19156 21956
rect 19208 21944 19214 21956
rect 19702 21944 19708 21956
rect 19208 21916 19708 21944
rect 19208 21904 19214 21916
rect 19702 21904 19708 21916
rect 19760 21904 19766 21956
rect 22204 21944 22232 21975
rect 25590 21972 25596 21984
rect 25648 21972 25654 22024
rect 22738 21944 22744 21956
rect 22204 21916 22744 21944
rect 22738 21904 22744 21916
rect 22796 21944 22802 21956
rect 22796 21916 23152 21944
rect 22796 21904 22802 21916
rect 3878 21876 3884 21888
rect 3839 21848 3884 21876
rect 3878 21836 3884 21848
rect 3936 21836 3942 21888
rect 9766 21836 9772 21888
rect 9824 21876 9830 21888
rect 10134 21876 10140 21888
rect 9824 21848 9869 21876
rect 10095 21848 10140 21876
rect 9824 21836 9830 21848
rect 10134 21836 10140 21848
rect 10192 21836 10198 21888
rect 13173 21879 13231 21885
rect 13173 21845 13185 21879
rect 13219 21876 13231 21879
rect 13354 21876 13360 21888
rect 13219 21848 13360 21876
rect 13219 21845 13231 21848
rect 13173 21839 13231 21845
rect 13354 21836 13360 21848
rect 13412 21836 13418 21888
rect 17494 21876 17500 21888
rect 17455 21848 17500 21876
rect 17494 21836 17500 21848
rect 17552 21836 17558 21888
rect 17954 21876 17960 21888
rect 17915 21848 17960 21876
rect 17954 21836 17960 21848
rect 18012 21836 18018 21888
rect 20533 21879 20591 21885
rect 20533 21845 20545 21879
rect 20579 21876 20591 21879
rect 20898 21876 20904 21888
rect 20579 21848 20904 21876
rect 20579 21845 20591 21848
rect 20533 21839 20591 21845
rect 20898 21836 20904 21848
rect 20956 21836 20962 21888
rect 23124 21885 23152 21916
rect 24762 21904 24768 21956
rect 24820 21944 24826 21956
rect 25317 21947 25375 21953
rect 25317 21944 25329 21947
rect 24820 21916 25329 21944
rect 24820 21904 24826 21916
rect 25317 21913 25329 21916
rect 25363 21913 25375 21947
rect 25317 21907 25375 21913
rect 27893 21947 27951 21953
rect 27893 21913 27905 21947
rect 27939 21944 27951 21947
rect 28442 21944 28448 21956
rect 27939 21916 28448 21944
rect 27939 21913 27951 21916
rect 27893 21907 27951 21913
rect 28442 21904 28448 21916
rect 28500 21904 28506 21956
rect 23109 21879 23167 21885
rect 23109 21845 23121 21879
rect 23155 21845 23167 21879
rect 23109 21839 23167 21845
rect 23569 21879 23627 21885
rect 23569 21845 23581 21879
rect 23615 21876 23627 21879
rect 24118 21876 24124 21888
rect 23615 21848 24124 21876
rect 23615 21845 23627 21848
rect 23569 21839 23627 21845
rect 24118 21836 24124 21848
rect 24176 21836 24182 21888
rect 24578 21836 24584 21888
rect 24636 21876 24642 21888
rect 26605 21879 26663 21885
rect 26605 21876 26617 21879
rect 24636 21848 26617 21876
rect 24636 21836 24642 21848
rect 26605 21845 26617 21848
rect 26651 21876 26663 21879
rect 26970 21876 26976 21888
rect 26651 21848 26976 21876
rect 26651 21845 26663 21848
rect 26605 21839 26663 21845
rect 26970 21836 26976 21848
rect 27028 21836 27034 21888
rect 27246 21836 27252 21888
rect 27304 21876 27310 21888
rect 27525 21879 27583 21885
rect 27525 21876 27537 21879
rect 27304 21848 27537 21876
rect 27304 21836 27310 21848
rect 27525 21845 27537 21848
rect 27571 21845 27583 21879
rect 27982 21876 27988 21888
rect 27943 21848 27988 21876
rect 27525 21839 27583 21845
rect 27982 21836 27988 21848
rect 28040 21836 28046 21888
rect 1104 21786 29600 21808
rect 1104 21734 8034 21786
rect 8086 21734 8098 21786
rect 8150 21734 8162 21786
rect 8214 21734 8226 21786
rect 8278 21734 8290 21786
rect 8342 21734 15118 21786
rect 15170 21734 15182 21786
rect 15234 21734 15246 21786
rect 15298 21734 15310 21786
rect 15362 21734 15374 21786
rect 15426 21734 22202 21786
rect 22254 21734 22266 21786
rect 22318 21734 22330 21786
rect 22382 21734 22394 21786
rect 22446 21734 22458 21786
rect 22510 21734 29286 21786
rect 29338 21734 29350 21786
rect 29402 21734 29414 21786
rect 29466 21734 29478 21786
rect 29530 21734 29542 21786
rect 29594 21734 29600 21786
rect 1104 21712 29600 21734
rect 4338 21632 4344 21684
rect 4396 21672 4402 21684
rect 4617 21675 4675 21681
rect 4617 21672 4629 21675
rect 4396 21644 4629 21672
rect 4396 21632 4402 21644
rect 4617 21641 4629 21644
rect 4663 21641 4675 21675
rect 8662 21672 8668 21684
rect 8623 21644 8668 21672
rect 4617 21635 4675 21641
rect 8662 21632 8668 21644
rect 8720 21632 8726 21684
rect 8938 21632 8944 21684
rect 8996 21672 9002 21684
rect 9217 21675 9275 21681
rect 9217 21672 9229 21675
rect 8996 21644 9229 21672
rect 8996 21632 9002 21644
rect 9217 21641 9229 21644
rect 9263 21641 9275 21675
rect 9217 21635 9275 21641
rect 9674 21632 9680 21684
rect 9732 21632 9738 21684
rect 10502 21632 10508 21684
rect 10560 21672 10566 21684
rect 10873 21675 10931 21681
rect 10873 21672 10885 21675
rect 10560 21644 10885 21672
rect 10560 21632 10566 21644
rect 10873 21641 10885 21644
rect 10919 21641 10931 21675
rect 10873 21635 10931 21641
rect 12894 21632 12900 21684
rect 12952 21672 12958 21684
rect 13906 21672 13912 21684
rect 12952 21644 13912 21672
rect 12952 21632 12958 21644
rect 13906 21632 13912 21644
rect 13964 21632 13970 21684
rect 14090 21672 14096 21684
rect 14051 21644 14096 21672
rect 14090 21632 14096 21644
rect 14148 21632 14154 21684
rect 14274 21632 14280 21684
rect 14332 21632 14338 21684
rect 14366 21632 14372 21684
rect 14424 21672 14430 21684
rect 15749 21675 15807 21681
rect 15749 21672 15761 21675
rect 14424 21644 15761 21672
rect 14424 21632 14430 21644
rect 15749 21641 15761 21644
rect 15795 21641 15807 21675
rect 15749 21635 15807 21641
rect 16942 21632 16948 21684
rect 17000 21672 17006 21684
rect 18233 21675 18291 21681
rect 18233 21672 18245 21675
rect 17000 21644 18245 21672
rect 17000 21632 17006 21644
rect 18233 21641 18245 21644
rect 18279 21672 18291 21675
rect 18279 21644 19334 21672
rect 18279 21641 18291 21644
rect 18233 21635 18291 21641
rect 9692 21604 9720 21632
rect 10042 21604 10048 21616
rect 3436 21576 4384 21604
rect 3436 21545 3464 21576
rect 4356 21548 4384 21576
rect 9416 21576 10048 21604
rect 3421 21539 3479 21545
rect 3421 21505 3433 21539
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 4154 21496 4160 21548
rect 4212 21536 4218 21548
rect 4249 21539 4307 21545
rect 4249 21536 4261 21539
rect 4212 21508 4261 21536
rect 4212 21496 4218 21508
rect 4249 21505 4261 21508
rect 4295 21505 4307 21539
rect 4249 21499 4307 21505
rect 4338 21496 4344 21548
rect 4396 21536 4402 21548
rect 9416 21545 9444 21576
rect 10042 21564 10048 21576
rect 10100 21564 10106 21616
rect 12713 21607 12771 21613
rect 12713 21573 12725 21607
rect 12759 21604 12771 21607
rect 14292 21604 14320 21632
rect 14461 21607 14519 21613
rect 14461 21604 14473 21607
rect 12759 21576 14473 21604
rect 12759 21573 12771 21576
rect 12713 21567 12771 21573
rect 14461 21573 14473 21576
rect 14507 21604 14519 21607
rect 15105 21607 15163 21613
rect 15105 21604 15117 21607
rect 14507 21576 15117 21604
rect 14507 21573 14519 21576
rect 14461 21567 14519 21573
rect 15105 21573 15117 21576
rect 15151 21573 15163 21607
rect 15105 21567 15163 21573
rect 15197 21607 15255 21613
rect 15197 21573 15209 21607
rect 15243 21604 15255 21607
rect 15378 21604 15384 21616
rect 15243 21576 15384 21604
rect 15243 21573 15255 21576
rect 15197 21567 15255 21573
rect 15378 21564 15384 21576
rect 15436 21564 15442 21616
rect 17954 21604 17960 21616
rect 16868 21576 17960 21604
rect 4433 21539 4491 21545
rect 4433 21536 4445 21539
rect 4396 21508 4445 21536
rect 4396 21496 4402 21508
rect 4433 21505 4445 21508
rect 4479 21505 4491 21539
rect 4433 21499 4491 21505
rect 9396 21539 9454 21545
rect 9396 21505 9408 21539
rect 9442 21505 9454 21539
rect 9396 21499 9454 21505
rect 9484 21539 9542 21545
rect 9484 21505 9496 21539
rect 9530 21505 9542 21539
rect 9484 21499 9542 21505
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21505 9643 21539
rect 9585 21499 9643 21505
rect 3510 21468 3516 21480
rect 3471 21440 3516 21468
rect 3510 21428 3516 21440
rect 3568 21428 3574 21480
rect 2501 21335 2559 21341
rect 2501 21301 2513 21335
rect 2547 21332 2559 21335
rect 2958 21332 2964 21344
rect 2547 21304 2964 21332
rect 2547 21301 2559 21304
rect 2501 21295 2559 21301
rect 2958 21292 2964 21304
rect 3016 21292 3022 21344
rect 3694 21332 3700 21344
rect 3655 21304 3700 21332
rect 3694 21292 3700 21304
rect 3752 21292 3758 21344
rect 8662 21292 8668 21344
rect 8720 21332 8726 21344
rect 9508 21332 9536 21499
rect 9600 21412 9628 21499
rect 9674 21496 9680 21548
rect 9732 21545 9738 21548
rect 9732 21539 9771 21545
rect 9759 21505 9771 21539
rect 9732 21499 9771 21505
rect 9861 21539 9919 21545
rect 9861 21505 9873 21539
rect 9907 21536 9919 21539
rect 12434 21536 12440 21548
rect 9907 21508 12440 21536
rect 9907 21505 9919 21508
rect 9861 21499 9919 21505
rect 9732 21496 9738 21499
rect 12434 21496 12440 21508
rect 12492 21496 12498 21548
rect 12621 21539 12679 21545
rect 12621 21505 12633 21539
rect 12667 21536 12679 21539
rect 12805 21539 12863 21545
rect 12667 21508 12756 21536
rect 12667 21505 12679 21508
rect 12621 21499 12679 21505
rect 12728 21480 12756 21508
rect 12805 21505 12817 21539
rect 12851 21536 12863 21539
rect 12894 21536 12900 21548
rect 12851 21508 12900 21536
rect 12851 21505 12863 21508
rect 12805 21499 12863 21505
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21505 13323 21539
rect 13265 21499 13323 21505
rect 9692 21440 12434 21468
rect 9582 21360 9588 21412
rect 9640 21360 9646 21412
rect 9692 21332 9720 21440
rect 9766 21360 9772 21412
rect 9824 21400 9830 21412
rect 10321 21403 10379 21409
rect 10321 21400 10333 21403
rect 9824 21372 10333 21400
rect 9824 21360 9830 21372
rect 10321 21369 10333 21372
rect 10367 21369 10379 21403
rect 12406 21400 12434 21440
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 13170 21468 13176 21480
rect 12768 21440 13176 21468
rect 12768 21428 12774 21440
rect 13170 21428 13176 21440
rect 13228 21428 13234 21480
rect 13280 21468 13308 21499
rect 13354 21496 13360 21548
rect 13412 21536 13418 21548
rect 13449 21539 13507 21545
rect 13449 21536 13461 21539
rect 13412 21508 13461 21536
rect 13412 21496 13418 21508
rect 13449 21505 13461 21508
rect 13495 21536 13507 21539
rect 13998 21536 14004 21548
rect 13495 21508 14004 21536
rect 13495 21505 13507 21508
rect 13449 21499 13507 21505
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 14277 21539 14335 21545
rect 14277 21505 14289 21539
rect 14323 21505 14335 21539
rect 14277 21499 14335 21505
rect 13538 21468 13544 21480
rect 13280 21440 13544 21468
rect 13538 21428 13544 21440
rect 13596 21428 13602 21480
rect 14292 21468 14320 21499
rect 14366 21496 14372 21548
rect 14424 21536 14430 21548
rect 14645 21539 14703 21545
rect 14424 21508 14469 21536
rect 14424 21496 14430 21508
rect 14645 21505 14657 21539
rect 14691 21536 14703 21539
rect 14918 21536 14924 21548
rect 14691 21508 14924 21536
rect 14691 21505 14703 21508
rect 14645 21499 14703 21505
rect 14918 21496 14924 21508
rect 14976 21496 14982 21548
rect 15473 21539 15531 21545
rect 15120 21508 15424 21536
rect 15120 21468 15148 21508
rect 14292 21440 15148 21468
rect 15396 21468 15424 21508
rect 15473 21505 15485 21539
rect 15519 21534 15531 21539
rect 16868 21536 16896 21576
rect 17954 21564 17960 21576
rect 18012 21564 18018 21616
rect 18325 21607 18383 21613
rect 18325 21573 18337 21607
rect 18371 21604 18383 21607
rect 18690 21604 18696 21616
rect 18371 21576 18696 21604
rect 18371 21573 18383 21576
rect 18325 21567 18383 21573
rect 18690 21564 18696 21576
rect 18748 21564 18754 21616
rect 19306 21604 19334 21644
rect 19702 21632 19708 21684
rect 19760 21672 19766 21684
rect 21358 21672 21364 21684
rect 19760 21644 21364 21672
rect 19760 21632 19766 21644
rect 21358 21632 21364 21644
rect 21416 21672 21422 21684
rect 21821 21675 21879 21681
rect 21821 21672 21833 21675
rect 21416 21644 21833 21672
rect 21416 21632 21422 21644
rect 21821 21641 21833 21644
rect 21867 21672 21879 21675
rect 24026 21672 24032 21684
rect 21867 21644 24032 21672
rect 21867 21641 21879 21644
rect 21821 21635 21879 21641
rect 24026 21632 24032 21644
rect 24084 21672 24090 21684
rect 27341 21675 27399 21681
rect 27341 21672 27353 21675
rect 24084 21644 27353 21672
rect 24084 21632 24090 21644
rect 27341 21641 27353 21644
rect 27387 21672 27399 21675
rect 27982 21672 27988 21684
rect 27387 21644 27988 21672
rect 27387 21641 27399 21644
rect 27341 21635 27399 21641
rect 27982 21632 27988 21644
rect 28040 21672 28046 21684
rect 28534 21672 28540 21684
rect 28040 21644 28540 21672
rect 28040 21632 28046 21644
rect 28534 21632 28540 21644
rect 28592 21632 28598 21684
rect 23106 21604 23112 21616
rect 19306 21576 20300 21604
rect 23019 21576 23112 21604
rect 17034 21536 17040 21548
rect 15580 21534 16896 21536
rect 15519 21508 16896 21534
rect 16995 21508 17040 21536
rect 15519 21506 15608 21508
rect 15519 21505 15531 21506
rect 15473 21499 15531 21505
rect 17034 21496 17040 21508
rect 17092 21496 17098 21548
rect 15565 21471 15623 21477
rect 15396 21440 15516 21468
rect 15488 21400 15516 21440
rect 15565 21437 15577 21471
rect 15611 21468 15623 21471
rect 16574 21468 16580 21480
rect 15611 21440 16580 21468
rect 15611 21437 15623 21440
rect 15565 21431 15623 21437
rect 16574 21428 16580 21440
rect 16632 21428 16638 21480
rect 17126 21468 17132 21480
rect 17087 21440 17132 21468
rect 17126 21428 17132 21440
rect 17184 21428 17190 21480
rect 17310 21468 17316 21480
rect 17271 21440 17316 21468
rect 17310 21428 17316 21440
rect 17368 21428 17374 21480
rect 17770 21428 17776 21480
rect 17828 21468 17834 21480
rect 20272 21477 20300 21576
rect 20806 21536 20812 21548
rect 20767 21508 20812 21536
rect 20806 21496 20812 21508
rect 20864 21496 20870 21548
rect 20898 21496 20904 21548
rect 20956 21536 20962 21548
rect 20993 21539 21051 21545
rect 20993 21536 21005 21539
rect 20956 21508 21005 21536
rect 20956 21496 20962 21508
rect 20993 21505 21005 21508
rect 21039 21505 21051 21539
rect 20993 21499 21051 21505
rect 21726 21496 21732 21548
rect 21784 21536 21790 21548
rect 23032 21545 23060 21576
rect 23106 21564 23112 21576
rect 23164 21604 23170 21616
rect 26145 21607 26203 21613
rect 23164 21576 24072 21604
rect 23164 21564 23170 21576
rect 24044 21548 24072 21576
rect 26145 21573 26157 21607
rect 26191 21604 26203 21607
rect 27614 21604 27620 21616
rect 26191 21576 27620 21604
rect 26191 21573 26203 21576
rect 26145 21567 26203 21573
rect 27614 21564 27620 21576
rect 27672 21564 27678 21616
rect 22465 21539 22523 21545
rect 22465 21536 22477 21539
rect 21784 21508 22477 21536
rect 21784 21496 21790 21508
rect 22465 21505 22477 21508
rect 22511 21505 22523 21539
rect 22465 21499 22523 21505
rect 23017 21539 23075 21545
rect 23017 21505 23029 21539
rect 23063 21505 23075 21539
rect 23017 21499 23075 21505
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21505 23443 21539
rect 24026 21536 24032 21548
rect 23987 21508 24032 21536
rect 23385 21499 23443 21505
rect 18509 21471 18567 21477
rect 18509 21468 18521 21471
rect 17828 21440 18521 21468
rect 17828 21428 17834 21440
rect 18509 21437 18521 21440
rect 18555 21468 18567 21471
rect 20257 21471 20315 21477
rect 18555 21440 19748 21468
rect 18555 21437 18567 21440
rect 18509 21431 18567 21437
rect 16482 21400 16488 21412
rect 12406 21372 15148 21400
rect 15488 21372 16488 21400
rect 10321 21363 10379 21369
rect 8720 21304 9720 21332
rect 8720 21292 8726 21304
rect 10870 21292 10876 21344
rect 10928 21332 10934 21344
rect 11517 21335 11575 21341
rect 11517 21332 11529 21335
rect 10928 21304 11529 21332
rect 10928 21292 10934 21304
rect 11517 21301 11529 21304
rect 11563 21301 11575 21335
rect 11517 21295 11575 21301
rect 13449 21335 13507 21341
rect 13449 21301 13461 21335
rect 13495 21332 13507 21335
rect 14366 21332 14372 21344
rect 13495 21304 14372 21332
rect 13495 21301 13507 21304
rect 13449 21295 13507 21301
rect 14366 21292 14372 21304
rect 14424 21292 14430 21344
rect 15120 21332 15148 21372
rect 16482 21360 16488 21372
rect 16540 21400 16546 21412
rect 16669 21403 16727 21409
rect 16669 21400 16681 21403
rect 16540 21372 16681 21400
rect 16540 21360 16546 21372
rect 16669 21369 16681 21372
rect 16715 21369 16727 21403
rect 18690 21400 18696 21412
rect 16669 21363 16727 21369
rect 17328 21372 18696 21400
rect 17328 21332 17356 21372
rect 18690 21360 18696 21372
rect 18748 21400 18754 21412
rect 19061 21403 19119 21409
rect 19061 21400 19073 21403
rect 18748 21372 19073 21400
rect 18748 21360 18754 21372
rect 19061 21369 19073 21372
rect 19107 21400 19119 21403
rect 19334 21400 19340 21412
rect 19107 21372 19340 21400
rect 19107 21369 19119 21372
rect 19061 21363 19119 21369
rect 19334 21360 19340 21372
rect 19392 21360 19398 21412
rect 19720 21409 19748 21440
rect 20257 21437 20269 21471
rect 20303 21468 20315 21471
rect 21634 21468 21640 21480
rect 20303 21440 21640 21468
rect 20303 21437 20315 21440
rect 20257 21431 20315 21437
rect 21634 21428 21640 21440
rect 21692 21468 21698 21480
rect 23106 21468 23112 21480
rect 21692 21440 23112 21468
rect 21692 21428 21698 21440
rect 23106 21428 23112 21440
rect 23164 21428 23170 21480
rect 23400 21468 23428 21499
rect 24026 21496 24032 21508
rect 24084 21496 24090 21548
rect 24118 21496 24124 21548
rect 24176 21536 24182 21548
rect 24176 21508 24221 21536
rect 24176 21496 24182 21508
rect 24762 21496 24768 21548
rect 24820 21536 24826 21548
rect 25225 21539 25283 21545
rect 25225 21536 25237 21539
rect 24820 21508 25237 21536
rect 24820 21496 24826 21508
rect 25225 21505 25237 21508
rect 25271 21505 25283 21539
rect 28718 21536 28724 21548
rect 28679 21508 28724 21536
rect 25225 21499 25283 21505
rect 28718 21496 28724 21508
rect 28776 21496 28782 21548
rect 23658 21468 23664 21480
rect 23400 21440 23664 21468
rect 23658 21428 23664 21440
rect 23716 21468 23722 21480
rect 24305 21471 24363 21477
rect 24305 21468 24317 21471
rect 23716 21440 24317 21468
rect 23716 21428 23722 21440
rect 24305 21437 24317 21440
rect 24351 21468 24363 21471
rect 26418 21468 26424 21480
rect 24351 21440 26424 21468
rect 24351 21437 24363 21440
rect 24305 21431 24363 21437
rect 26418 21428 26424 21440
rect 26476 21428 26482 21480
rect 26878 21428 26884 21480
rect 26936 21468 26942 21480
rect 27433 21471 27491 21477
rect 27433 21468 27445 21471
rect 26936 21440 27445 21468
rect 26936 21428 26942 21440
rect 27433 21437 27445 21440
rect 27479 21437 27491 21471
rect 27433 21431 27491 21437
rect 27522 21428 27528 21480
rect 27580 21468 27586 21480
rect 27580 21440 27625 21468
rect 27580 21428 27586 21440
rect 19705 21403 19763 21409
rect 19705 21369 19717 21403
rect 19751 21400 19763 21403
rect 19886 21400 19892 21412
rect 19751 21372 19892 21400
rect 19751 21369 19763 21372
rect 19705 21363 19763 21369
rect 19886 21360 19892 21372
rect 19944 21400 19950 21412
rect 19944 21372 21404 21400
rect 19944 21360 19950 21372
rect 21376 21344 21404 21372
rect 22554 21360 22560 21412
rect 22612 21400 22618 21412
rect 23293 21403 23351 21409
rect 23293 21400 23305 21403
rect 22612 21372 23305 21400
rect 22612 21360 22618 21372
rect 23293 21369 23305 21372
rect 23339 21369 23351 21403
rect 23293 21363 23351 21369
rect 24026 21360 24032 21412
rect 24084 21400 24090 21412
rect 25501 21403 25559 21409
rect 25501 21400 25513 21403
rect 24084 21372 25513 21400
rect 24084 21360 24090 21372
rect 25501 21369 25513 21372
rect 25547 21400 25559 21403
rect 26510 21400 26516 21412
rect 25547 21372 26516 21400
rect 25547 21369 25559 21372
rect 25501 21363 25559 21369
rect 26510 21360 26516 21372
rect 26568 21360 26574 21412
rect 15120 21304 17356 21332
rect 17402 21292 17408 21344
rect 17460 21332 17466 21344
rect 17865 21335 17923 21341
rect 17865 21332 17877 21335
rect 17460 21304 17877 21332
rect 17460 21292 17466 21304
rect 17865 21301 17877 21304
rect 17911 21301 17923 21335
rect 20898 21332 20904 21344
rect 20859 21304 20904 21332
rect 17865 21295 17923 21301
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 21358 21292 21364 21344
rect 21416 21292 21422 21344
rect 23566 21292 23572 21344
rect 23624 21332 23630 21344
rect 24213 21335 24271 21341
rect 24213 21332 24225 21335
rect 23624 21304 24225 21332
rect 23624 21292 23630 21304
rect 24213 21301 24225 21304
rect 24259 21301 24271 21335
rect 24213 21295 24271 21301
rect 26234 21292 26240 21344
rect 26292 21332 26298 21344
rect 26973 21335 27031 21341
rect 26973 21332 26985 21335
rect 26292 21304 26985 21332
rect 26292 21292 26298 21304
rect 26973 21301 26985 21304
rect 27019 21301 27031 21335
rect 26973 21295 27031 21301
rect 1104 21242 29440 21264
rect 1104 21190 4492 21242
rect 4544 21190 4556 21242
rect 4608 21190 4620 21242
rect 4672 21190 4684 21242
rect 4736 21190 4748 21242
rect 4800 21190 11576 21242
rect 11628 21190 11640 21242
rect 11692 21190 11704 21242
rect 11756 21190 11768 21242
rect 11820 21190 11832 21242
rect 11884 21190 18660 21242
rect 18712 21190 18724 21242
rect 18776 21190 18788 21242
rect 18840 21190 18852 21242
rect 18904 21190 18916 21242
rect 18968 21190 25744 21242
rect 25796 21190 25808 21242
rect 25860 21190 25872 21242
rect 25924 21190 25936 21242
rect 25988 21190 26000 21242
rect 26052 21190 29440 21242
rect 1104 21168 29440 21190
rect 9309 21131 9367 21137
rect 9309 21097 9321 21131
rect 9355 21128 9367 21131
rect 9674 21128 9680 21140
rect 9355 21100 9680 21128
rect 9355 21097 9367 21100
rect 9309 21091 9367 21097
rect 9674 21088 9680 21100
rect 9732 21088 9738 21140
rect 10594 21088 10600 21140
rect 10652 21128 10658 21140
rect 11609 21131 11667 21137
rect 11609 21128 11621 21131
rect 10652 21100 11621 21128
rect 10652 21088 10658 21100
rect 11609 21097 11621 21100
rect 11655 21097 11667 21131
rect 11609 21091 11667 21097
rect 12434 21088 12440 21140
rect 12492 21128 12498 21140
rect 13538 21128 13544 21140
rect 12492 21100 12537 21128
rect 13499 21100 13544 21128
rect 12492 21088 12498 21100
rect 13538 21088 13544 21100
rect 13596 21088 13602 21140
rect 16574 21128 16580 21140
rect 16535 21100 16580 21128
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 17126 21088 17132 21140
rect 17184 21128 17190 21140
rect 17221 21131 17279 21137
rect 17221 21128 17233 21131
rect 17184 21100 17233 21128
rect 17184 21088 17190 21100
rect 17221 21097 17233 21100
rect 17267 21097 17279 21131
rect 17221 21091 17279 21097
rect 17310 21088 17316 21140
rect 17368 21128 17374 21140
rect 17865 21131 17923 21137
rect 17865 21128 17877 21131
rect 17368 21100 17877 21128
rect 17368 21088 17374 21100
rect 17865 21097 17877 21100
rect 17911 21128 17923 21131
rect 18322 21128 18328 21140
rect 17911 21100 18328 21128
rect 17911 21097 17923 21100
rect 17865 21091 17923 21097
rect 18322 21088 18328 21100
rect 18380 21088 18386 21140
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 26050 21128 26056 21140
rect 19392 21100 26056 21128
rect 19392 21088 19398 21100
rect 26050 21088 26056 21100
rect 26108 21088 26114 21140
rect 26234 21128 26240 21140
rect 26195 21100 26240 21128
rect 26234 21088 26240 21100
rect 26292 21088 26298 21140
rect 27706 21088 27712 21140
rect 27764 21128 27770 21140
rect 28166 21128 28172 21140
rect 27764 21100 28172 21128
rect 27764 21088 27770 21100
rect 28166 21088 28172 21100
rect 28224 21088 28230 21140
rect 8389 21063 8447 21069
rect 8389 21029 8401 21063
rect 8435 21060 8447 21063
rect 9490 21060 9496 21072
rect 8435 21032 9496 21060
rect 8435 21029 8447 21032
rect 8389 21023 8447 21029
rect 9490 21020 9496 21032
rect 9548 21060 9554 21072
rect 9548 21032 9812 21060
rect 9548 21020 9554 21032
rect 9490 20924 9496 20936
rect 9451 20896 9496 20924
rect 9490 20884 9496 20896
rect 9548 20884 9554 20936
rect 9784 20933 9812 21032
rect 10778 21020 10784 21072
rect 10836 21060 10842 21072
rect 16942 21060 16948 21072
rect 10836 21032 16948 21060
rect 10836 21020 10842 21032
rect 16942 21020 16948 21032
rect 17000 21020 17006 21072
rect 17144 20992 17172 21088
rect 26789 21063 26847 21069
rect 26789 21060 26801 21063
rect 20916 21032 26801 21060
rect 20806 20992 20812 21004
rect 14476 20964 14872 20992
rect 9658 20927 9716 20933
rect 9658 20893 9670 20927
rect 9704 20924 9716 20927
rect 9769 20927 9827 20933
rect 9704 20893 9720 20924
rect 9658 20887 9720 20893
rect 9769 20893 9781 20927
rect 9815 20893 9827 20927
rect 10134 20924 10140 20936
rect 9968 20918 10140 20924
rect 9876 20911 10140 20918
rect 9769 20887 9827 20893
rect 9861 20905 10140 20911
rect 6546 20788 6552 20800
rect 6507 20760 6552 20788
rect 6546 20748 6552 20760
rect 6604 20748 6610 20800
rect 7837 20791 7895 20797
rect 7837 20757 7849 20791
rect 7883 20788 7895 20791
rect 7926 20788 7932 20800
rect 7883 20760 7932 20788
rect 7883 20757 7895 20760
rect 7837 20751 7895 20757
rect 7926 20748 7932 20760
rect 7984 20788 7990 20800
rect 9692 20788 9720 20887
rect 7984 20760 9720 20788
rect 9784 20788 9812 20887
rect 9861 20871 9873 20905
rect 9907 20896 10140 20905
rect 9907 20890 9996 20896
rect 9907 20871 9919 20890
rect 10134 20884 10140 20896
rect 10192 20884 10198 20936
rect 10502 20884 10508 20936
rect 10560 20924 10566 20936
rect 11517 20927 11575 20933
rect 11517 20924 11529 20927
rect 10560 20896 11529 20924
rect 10560 20884 10566 20896
rect 11517 20893 11529 20896
rect 11563 20924 11575 20927
rect 11974 20924 11980 20936
rect 11563 20896 11980 20924
rect 11563 20893 11575 20896
rect 11517 20887 11575 20893
rect 11974 20884 11980 20896
rect 12032 20884 12038 20936
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20893 12495 20927
rect 12618 20924 12624 20936
rect 12579 20896 12624 20924
rect 12437 20887 12495 20893
rect 9861 20865 9919 20871
rect 10870 20856 10876 20868
rect 10428 20828 10876 20856
rect 10428 20788 10456 20828
rect 10870 20816 10876 20828
rect 10928 20816 10934 20868
rect 12452 20856 12480 20887
rect 12618 20884 12624 20896
rect 12676 20884 12682 20936
rect 14090 20884 14096 20936
rect 14148 20924 14154 20936
rect 14272 20927 14330 20933
rect 14272 20924 14284 20927
rect 14148 20896 14284 20924
rect 14148 20884 14154 20896
rect 14272 20893 14284 20896
rect 14318 20924 14330 20927
rect 14476 20924 14504 20964
rect 14642 20924 14648 20936
rect 14318 20896 14504 20924
rect 14603 20896 14648 20924
rect 14318 20893 14330 20896
rect 14272 20887 14330 20893
rect 14642 20884 14648 20896
rect 14700 20884 14706 20936
rect 14737 20927 14795 20933
rect 14737 20893 14749 20927
rect 14783 20893 14795 20927
rect 14737 20887 14795 20893
rect 12452 20828 14136 20856
rect 10594 20788 10600 20800
rect 9784 20760 10456 20788
rect 10555 20760 10600 20788
rect 7984 20748 7990 20760
rect 10594 20748 10600 20760
rect 10652 20748 10658 20800
rect 14108 20797 14136 20828
rect 14182 20816 14188 20868
rect 14240 20856 14246 20868
rect 14366 20856 14372 20868
rect 14240 20828 14372 20856
rect 14240 20816 14246 20828
rect 14366 20816 14372 20828
rect 14424 20816 14430 20868
rect 14461 20859 14519 20865
rect 14461 20825 14473 20859
rect 14507 20825 14519 20859
rect 14461 20819 14519 20825
rect 14093 20791 14151 20797
rect 14093 20757 14105 20791
rect 14139 20757 14151 20791
rect 14093 20751 14151 20757
rect 14274 20748 14280 20800
rect 14332 20788 14338 20800
rect 14476 20788 14504 20819
rect 14550 20816 14556 20868
rect 14608 20856 14614 20868
rect 14752 20856 14780 20887
rect 14608 20828 14780 20856
rect 14844 20856 14872 20964
rect 16592 20964 17172 20992
rect 17236 20964 20812 20992
rect 16390 20924 16396 20936
rect 16351 20896 16396 20924
rect 16390 20884 16396 20896
rect 16448 20884 16454 20936
rect 16592 20933 16620 20964
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20893 16635 20927
rect 16577 20887 16635 20893
rect 16850 20884 16856 20936
rect 16908 20924 16914 20936
rect 17129 20927 17187 20933
rect 17129 20924 17141 20927
rect 16908 20896 17141 20924
rect 16908 20884 16914 20896
rect 17129 20893 17141 20896
rect 17175 20924 17187 20927
rect 17236 20924 17264 20964
rect 17175 20896 17264 20924
rect 17313 20927 17371 20933
rect 17175 20893 17187 20896
rect 17129 20887 17187 20893
rect 17313 20893 17325 20927
rect 17359 20924 17371 20927
rect 17402 20924 17408 20936
rect 17359 20896 17408 20924
rect 17359 20893 17371 20896
rect 17313 20887 17371 20893
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 20732 20933 20760 20964
rect 20806 20952 20812 20964
rect 20864 20952 20870 21004
rect 20916 20933 20944 21032
rect 26789 21029 26801 21032
rect 26835 21029 26847 21063
rect 26789 21023 26847 21029
rect 26970 21020 26976 21072
rect 27028 21020 27034 21072
rect 21082 20952 21088 21004
rect 21140 20992 21146 21004
rect 22557 20995 22615 21001
rect 22557 20992 22569 20995
rect 21140 20964 22569 20992
rect 21140 20952 21146 20964
rect 22557 20961 22569 20964
rect 22603 20992 22615 20995
rect 24578 20992 24584 21004
rect 22603 20964 24584 20992
rect 22603 20961 22615 20964
rect 22557 20955 22615 20961
rect 24578 20952 24584 20964
rect 24636 20952 24642 21004
rect 26053 20995 26111 21001
rect 26053 20961 26065 20995
rect 26099 20992 26111 20995
rect 26418 20992 26424 21004
rect 26099 20964 26424 20992
rect 26099 20961 26111 20964
rect 26053 20955 26111 20961
rect 26418 20952 26424 20964
rect 26476 20992 26482 21004
rect 26694 20992 26700 21004
rect 26476 20964 26700 20992
rect 26476 20952 26482 20964
rect 26694 20952 26700 20964
rect 26752 20952 26758 21004
rect 26988 20992 27016 21020
rect 27433 20995 27491 21001
rect 27433 20992 27445 20995
rect 26988 20964 27445 20992
rect 27433 20961 27445 20964
rect 27479 20961 27491 20995
rect 27706 20992 27712 21004
rect 27667 20964 27712 20992
rect 27433 20955 27491 20961
rect 27706 20952 27712 20964
rect 27764 20952 27770 21004
rect 27985 20995 28043 21001
rect 27985 20961 27997 20995
rect 28031 20992 28043 20995
rect 28074 20992 28080 21004
rect 28031 20964 28080 20992
rect 28031 20961 28043 20964
rect 27985 20955 28043 20961
rect 28074 20952 28080 20964
rect 28132 20952 28138 21004
rect 20717 20927 20775 20933
rect 20717 20893 20729 20927
rect 20763 20893 20775 20927
rect 20717 20887 20775 20893
rect 20901 20927 20959 20933
rect 20901 20893 20913 20927
rect 20947 20893 20959 20927
rect 21634 20924 21640 20936
rect 21595 20896 21640 20924
rect 20901 20887 20959 20893
rect 21634 20884 21640 20896
rect 21692 20884 21698 20936
rect 23382 20924 23388 20936
rect 23343 20896 23388 20924
rect 23382 20884 23388 20896
rect 23440 20884 23446 20936
rect 23569 20927 23627 20933
rect 23569 20893 23581 20927
rect 23615 20924 23627 20927
rect 23658 20924 23664 20936
rect 23615 20896 23664 20924
rect 23615 20893 23627 20896
rect 23569 20887 23627 20893
rect 23658 20884 23664 20896
rect 23716 20884 23722 20936
rect 26329 20927 26387 20933
rect 26329 20893 26341 20927
rect 26375 20924 26387 20927
rect 26510 20924 26516 20936
rect 26375 20896 26516 20924
rect 26375 20893 26387 20896
rect 26329 20887 26387 20893
rect 26510 20884 26516 20896
rect 26568 20884 26574 20936
rect 27614 20933 27620 20936
rect 27592 20927 27620 20933
rect 27592 20893 27604 20927
rect 27592 20887 27620 20893
rect 27614 20884 27620 20887
rect 27672 20884 27678 20936
rect 28258 20884 28264 20936
rect 28316 20924 28322 20936
rect 28445 20927 28503 20933
rect 28445 20924 28457 20927
rect 28316 20896 28457 20924
rect 28316 20884 28322 20896
rect 28445 20893 28457 20896
rect 28491 20893 28503 20927
rect 28445 20887 28503 20893
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 20809 20859 20867 20865
rect 20809 20856 20821 20859
rect 14844 20828 20821 20856
rect 14608 20816 14614 20828
rect 20809 20825 20821 20828
rect 20855 20825 20867 20859
rect 20809 20819 20867 20825
rect 21358 20816 21364 20868
rect 21416 20856 21422 20868
rect 21913 20859 21971 20865
rect 21913 20856 21925 20859
rect 21416 20828 21925 20856
rect 21416 20816 21422 20828
rect 21913 20825 21925 20828
rect 21959 20856 21971 20859
rect 24486 20856 24492 20868
rect 21959 20828 24492 20856
rect 21959 20825 21971 20828
rect 21913 20819 21971 20825
rect 24486 20816 24492 20828
rect 24544 20856 24550 20868
rect 24544 20828 26280 20856
rect 24544 20816 24550 20828
rect 18690 20788 18696 20800
rect 14332 20760 14504 20788
rect 18651 20760 18696 20788
rect 14332 20748 14338 20760
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 19242 20788 19248 20800
rect 19203 20760 19248 20788
rect 19242 20748 19248 20760
rect 19300 20748 19306 20800
rect 23474 20788 23480 20800
rect 23435 20760 23480 20788
rect 23474 20748 23480 20760
rect 23532 20748 23538 20800
rect 23842 20748 23848 20800
rect 23900 20788 23906 20800
rect 24673 20791 24731 20797
rect 24673 20788 24685 20791
rect 23900 20760 24685 20788
rect 23900 20748 23906 20760
rect 24673 20757 24685 20760
rect 24719 20788 24731 20791
rect 24762 20788 24768 20800
rect 24719 20760 24768 20788
rect 24719 20757 24731 20760
rect 24673 20751 24731 20757
rect 24762 20748 24768 20760
rect 24820 20788 24826 20800
rect 25501 20791 25559 20797
rect 25501 20788 25513 20791
rect 24820 20760 25513 20788
rect 24820 20748 24826 20760
rect 25501 20757 25513 20760
rect 25547 20757 25559 20791
rect 25501 20751 25559 20757
rect 26053 20791 26111 20797
rect 26053 20757 26065 20791
rect 26099 20788 26111 20791
rect 26142 20788 26148 20800
rect 26099 20760 26148 20788
rect 26099 20757 26111 20760
rect 26053 20751 26111 20757
rect 26142 20748 26148 20760
rect 26200 20748 26206 20800
rect 26252 20788 26280 20828
rect 27522 20788 27528 20800
rect 26252 20760 27528 20788
rect 27522 20748 27528 20760
rect 27580 20748 27586 20800
rect 27798 20748 27804 20800
rect 27856 20788 27862 20800
rect 28644 20788 28672 20887
rect 27856 20760 28672 20788
rect 27856 20748 27862 20760
rect 1104 20698 29600 20720
rect 1104 20646 8034 20698
rect 8086 20646 8098 20698
rect 8150 20646 8162 20698
rect 8214 20646 8226 20698
rect 8278 20646 8290 20698
rect 8342 20646 15118 20698
rect 15170 20646 15182 20698
rect 15234 20646 15246 20698
rect 15298 20646 15310 20698
rect 15362 20646 15374 20698
rect 15426 20646 22202 20698
rect 22254 20646 22266 20698
rect 22318 20646 22330 20698
rect 22382 20646 22394 20698
rect 22446 20646 22458 20698
rect 22510 20646 29286 20698
rect 29338 20646 29350 20698
rect 29402 20646 29414 20698
rect 29466 20646 29478 20698
rect 29530 20646 29542 20698
rect 29594 20646 29600 20698
rect 1104 20624 29600 20646
rect 1854 20544 1860 20596
rect 1912 20584 1918 20596
rect 1949 20587 2007 20593
rect 1949 20584 1961 20587
rect 1912 20556 1961 20584
rect 1912 20544 1918 20556
rect 1949 20553 1961 20556
rect 1995 20584 2007 20587
rect 8294 20584 8300 20596
rect 1995 20556 8300 20584
rect 1995 20553 2007 20556
rect 1949 20547 2007 20553
rect 8294 20544 8300 20556
rect 8352 20544 8358 20596
rect 9766 20584 9772 20596
rect 9692 20556 9772 20584
rect 4338 20516 4344 20528
rect 3620 20488 4344 20516
rect 3142 20448 3148 20460
rect 3103 20420 3148 20448
rect 3142 20408 3148 20420
rect 3200 20408 3206 20460
rect 3234 20408 3240 20460
rect 3292 20448 3298 20460
rect 3620 20457 3648 20488
rect 4338 20476 4344 20488
rect 4396 20516 4402 20528
rect 9692 20525 9720 20556
rect 9766 20544 9772 20556
rect 9824 20544 9830 20596
rect 11974 20584 11980 20596
rect 11935 20556 11980 20584
rect 11974 20544 11980 20556
rect 12032 20544 12038 20596
rect 12618 20584 12624 20596
rect 12579 20556 12624 20584
rect 12618 20544 12624 20556
rect 12676 20544 12682 20596
rect 14274 20584 14280 20596
rect 13924 20556 14280 20584
rect 4617 20519 4675 20525
rect 4617 20516 4629 20519
rect 4396 20488 4629 20516
rect 4396 20476 4402 20488
rect 4617 20485 4629 20488
rect 4663 20485 4675 20519
rect 4617 20479 4675 20485
rect 9677 20519 9735 20525
rect 9677 20485 9689 20519
rect 9723 20485 9735 20519
rect 9677 20479 9735 20485
rect 3329 20451 3387 20457
rect 3329 20448 3341 20451
rect 3292 20420 3341 20448
rect 3292 20408 3298 20420
rect 3329 20417 3341 20420
rect 3375 20417 3387 20451
rect 3329 20411 3387 20417
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20417 3663 20451
rect 3605 20411 3663 20417
rect 4246 20408 4252 20460
rect 4304 20448 4310 20460
rect 4525 20451 4583 20457
rect 4525 20448 4537 20451
rect 4304 20420 4537 20448
rect 4304 20408 4310 20420
rect 4525 20417 4537 20420
rect 4571 20417 4583 20451
rect 4525 20411 4583 20417
rect 4709 20451 4767 20457
rect 4709 20417 4721 20451
rect 4755 20448 4767 20451
rect 5902 20448 5908 20460
rect 4755 20420 5908 20448
rect 4755 20417 4767 20420
rect 4709 20411 4767 20417
rect 5902 20408 5908 20420
rect 5960 20408 5966 20460
rect 7098 20448 7104 20460
rect 7011 20420 7104 20448
rect 7098 20408 7104 20420
rect 7156 20448 7162 20460
rect 7466 20448 7472 20460
rect 7156 20420 7472 20448
rect 7156 20408 7162 20420
rect 7466 20408 7472 20420
rect 7524 20408 7530 20460
rect 8294 20408 8300 20460
rect 8352 20448 8358 20460
rect 8757 20451 8815 20457
rect 8757 20448 8769 20451
rect 8352 20420 8769 20448
rect 8352 20408 8358 20420
rect 8757 20417 8769 20420
rect 8803 20417 8815 20451
rect 8757 20411 8815 20417
rect 8941 20451 8999 20457
rect 8941 20417 8953 20451
rect 8987 20448 8999 20451
rect 9122 20448 9128 20460
rect 8987 20420 9128 20448
rect 8987 20417 8999 20420
rect 8941 20411 8999 20417
rect 9122 20408 9128 20420
rect 9180 20448 9186 20460
rect 9493 20451 9551 20457
rect 9493 20448 9505 20451
rect 9180 20420 9505 20448
rect 9180 20408 9186 20420
rect 9493 20417 9505 20420
rect 9539 20417 9551 20451
rect 9493 20411 9551 20417
rect 9769 20451 9827 20457
rect 9769 20417 9781 20451
rect 9815 20417 9827 20451
rect 9769 20411 9827 20417
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 10502 20448 10508 20460
rect 9907 20420 10508 20448
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 3513 20383 3571 20389
rect 3513 20349 3525 20383
rect 3559 20380 3571 20383
rect 3878 20380 3884 20392
rect 3559 20352 3884 20380
rect 3559 20349 3571 20352
rect 3513 20343 3571 20349
rect 3878 20340 3884 20352
rect 3936 20340 3942 20392
rect 7006 20340 7012 20392
rect 7064 20380 7070 20392
rect 7193 20383 7251 20389
rect 7193 20380 7205 20383
rect 7064 20352 7205 20380
rect 7064 20340 7070 20352
rect 7193 20349 7205 20352
rect 7239 20380 7251 20383
rect 7282 20380 7288 20392
rect 7239 20352 7288 20380
rect 7239 20349 7251 20352
rect 7193 20343 7251 20349
rect 7282 20340 7288 20352
rect 7340 20340 7346 20392
rect 7374 20340 7380 20392
rect 7432 20380 7438 20392
rect 7561 20383 7619 20389
rect 7561 20380 7573 20383
rect 7432 20352 7573 20380
rect 7432 20340 7438 20352
rect 7561 20349 7573 20352
rect 7607 20349 7619 20383
rect 7561 20343 7619 20349
rect 7926 20340 7932 20392
rect 7984 20380 7990 20392
rect 8573 20383 8631 20389
rect 8573 20380 8585 20383
rect 7984 20352 8585 20380
rect 7984 20340 7990 20352
rect 8573 20349 8585 20352
rect 8619 20380 8631 20383
rect 9784 20380 9812 20411
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 12802 20448 12808 20460
rect 12763 20420 12808 20448
rect 12802 20408 12808 20420
rect 12860 20408 12866 20460
rect 13081 20451 13139 20457
rect 13081 20417 13093 20451
rect 13127 20448 13139 20451
rect 13262 20448 13268 20460
rect 13127 20420 13268 20448
rect 13127 20417 13139 20420
rect 13081 20411 13139 20417
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 13924 20457 13952 20556
rect 14274 20544 14280 20556
rect 14332 20544 14338 20596
rect 16390 20544 16396 20596
rect 16448 20584 16454 20596
rect 16574 20584 16580 20596
rect 16448 20556 16580 20584
rect 16448 20544 16454 20556
rect 16574 20544 16580 20556
rect 16632 20584 16638 20596
rect 16761 20587 16819 20593
rect 16761 20584 16773 20587
rect 16632 20556 16773 20584
rect 16632 20544 16638 20556
rect 16761 20553 16773 20556
rect 16807 20584 16819 20587
rect 17310 20584 17316 20596
rect 16807 20556 17316 20584
rect 16807 20553 16819 20556
rect 16761 20547 16819 20553
rect 17310 20544 17316 20556
rect 17368 20544 17374 20596
rect 17678 20544 17684 20596
rect 17736 20584 17742 20596
rect 17957 20587 18015 20593
rect 17957 20584 17969 20587
rect 17736 20556 17969 20584
rect 17736 20544 17742 20556
rect 17957 20553 17969 20556
rect 18003 20553 18015 20587
rect 25038 20584 25044 20596
rect 24999 20556 25044 20584
rect 17957 20547 18015 20553
rect 25038 20544 25044 20556
rect 25096 20544 25102 20596
rect 14090 20516 14096 20528
rect 14051 20488 14096 20516
rect 14090 20476 14096 20488
rect 14148 20476 14154 20528
rect 20898 20516 20904 20528
rect 14292 20488 20904 20516
rect 13909 20451 13967 20457
rect 13909 20417 13921 20451
rect 13955 20417 13967 20451
rect 14182 20448 14188 20460
rect 14143 20420 14188 20448
rect 13909 20411 13967 20417
rect 14182 20408 14188 20420
rect 14240 20408 14246 20460
rect 14292 20457 14320 20488
rect 20898 20476 20904 20488
rect 20956 20476 20962 20528
rect 23474 20476 23480 20528
rect 23532 20516 23538 20528
rect 25409 20519 25467 20525
rect 25409 20516 25421 20519
rect 23532 20488 25421 20516
rect 23532 20476 23538 20488
rect 25409 20485 25421 20488
rect 25455 20485 25467 20519
rect 25409 20479 25467 20485
rect 25590 20476 25596 20528
rect 25648 20516 25654 20528
rect 26970 20516 26976 20528
rect 25648 20488 26976 20516
rect 25648 20476 25654 20488
rect 26970 20476 26976 20488
rect 27028 20516 27034 20528
rect 27614 20516 27620 20528
rect 27028 20488 27620 20516
rect 27028 20476 27034 20488
rect 27614 20476 27620 20488
rect 27672 20476 27678 20528
rect 14277 20451 14335 20457
rect 14277 20417 14289 20451
rect 14323 20417 14335 20451
rect 14277 20411 14335 20417
rect 18690 20408 18696 20460
rect 18748 20448 18754 20460
rect 19058 20448 19064 20460
rect 18748 20420 19064 20448
rect 18748 20408 18754 20420
rect 19058 20408 19064 20420
rect 19116 20448 19122 20460
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 19116 20420 19257 20448
rect 19116 20408 19122 20420
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20448 19579 20451
rect 19886 20448 19892 20460
rect 19567 20420 19892 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 19886 20408 19892 20420
rect 19944 20448 19950 20460
rect 21634 20448 21640 20460
rect 19944 20420 21640 20448
rect 19944 20408 19950 20420
rect 21634 20408 21640 20420
rect 21692 20448 21698 20460
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 21692 20420 21833 20448
rect 21692 20408 21698 20420
rect 21821 20417 21833 20420
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 23842 20408 23848 20460
rect 23900 20448 23906 20460
rect 24213 20451 24271 20457
rect 24213 20448 24225 20451
rect 23900 20420 24225 20448
rect 23900 20408 23906 20420
rect 24213 20417 24225 20420
rect 24259 20417 24271 20451
rect 24486 20448 24492 20460
rect 24447 20420 24492 20448
rect 24213 20411 24271 20417
rect 24486 20408 24492 20420
rect 24544 20408 24550 20460
rect 25501 20451 25559 20457
rect 25501 20417 25513 20451
rect 25547 20448 25559 20451
rect 26142 20448 26148 20460
rect 25547 20420 26148 20448
rect 25547 20417 25559 20420
rect 25501 20411 25559 20417
rect 26142 20408 26148 20420
rect 26200 20408 26206 20460
rect 8619 20352 9812 20380
rect 19429 20383 19487 20389
rect 8619 20349 8631 20352
rect 8573 20343 8631 20349
rect 19429 20349 19441 20383
rect 19475 20380 19487 20383
rect 20806 20380 20812 20392
rect 19475 20352 20812 20380
rect 19475 20349 19487 20352
rect 19429 20343 19487 20349
rect 20806 20340 20812 20352
rect 20864 20340 20870 20392
rect 23753 20383 23811 20389
rect 23753 20349 23765 20383
rect 23799 20380 23811 20383
rect 24504 20380 24532 20408
rect 23799 20352 24532 20380
rect 24581 20383 24639 20389
rect 23799 20349 23811 20352
rect 23753 20343 23811 20349
rect 24581 20349 24593 20383
rect 24627 20380 24639 20383
rect 24762 20380 24768 20392
rect 24627 20352 24768 20380
rect 24627 20349 24639 20352
rect 24581 20343 24639 20349
rect 24762 20340 24768 20352
rect 24820 20340 24826 20392
rect 25685 20383 25743 20389
rect 25685 20349 25697 20383
rect 25731 20380 25743 20383
rect 26234 20380 26240 20392
rect 25731 20352 26240 20380
rect 25731 20349 25743 20352
rect 25685 20343 25743 20349
rect 26234 20340 26240 20352
rect 26292 20340 26298 20392
rect 1670 20272 1676 20324
rect 1728 20312 1734 20324
rect 2501 20315 2559 20321
rect 2501 20312 2513 20315
rect 1728 20284 2513 20312
rect 1728 20272 1734 20284
rect 2501 20281 2513 20284
rect 2547 20281 2559 20315
rect 2501 20275 2559 20281
rect 3421 20315 3479 20321
rect 3421 20281 3433 20315
rect 3467 20312 3479 20315
rect 4154 20312 4160 20324
rect 3467 20284 4160 20312
rect 3467 20281 3479 20284
rect 3421 20275 3479 20281
rect 4154 20272 4160 20284
rect 4212 20272 4218 20324
rect 19061 20315 19119 20321
rect 8266 20284 10640 20312
rect 3789 20247 3847 20253
rect 3789 20213 3801 20247
rect 3835 20244 3847 20247
rect 3970 20244 3976 20256
rect 3835 20216 3976 20244
rect 3835 20213 3847 20216
rect 3789 20207 3847 20213
rect 3970 20204 3976 20216
rect 4028 20204 4034 20256
rect 5813 20247 5871 20253
rect 5813 20213 5825 20247
rect 5859 20244 5871 20247
rect 6454 20244 6460 20256
rect 5859 20216 6460 20244
rect 5859 20213 5871 20216
rect 5813 20207 5871 20213
rect 6454 20204 6460 20216
rect 6512 20204 6518 20256
rect 6914 20244 6920 20256
rect 6875 20216 6920 20244
rect 6914 20204 6920 20216
rect 6972 20204 6978 20256
rect 7926 20204 7932 20256
rect 7984 20244 7990 20256
rect 8021 20247 8079 20253
rect 8021 20244 8033 20247
rect 7984 20216 8033 20244
rect 7984 20204 7990 20216
rect 8021 20213 8033 20216
rect 8067 20213 8079 20247
rect 8021 20207 8079 20213
rect 8110 20204 8116 20256
rect 8168 20244 8174 20256
rect 8266 20244 8294 20284
rect 8168 20216 8294 20244
rect 8168 20204 8174 20216
rect 9950 20204 9956 20256
rect 10008 20244 10014 20256
rect 10612 20253 10640 20284
rect 19061 20281 19073 20315
rect 19107 20312 19119 20315
rect 21634 20312 21640 20324
rect 19107 20284 21640 20312
rect 19107 20281 19119 20284
rect 19061 20275 19119 20281
rect 21634 20272 21640 20284
rect 21692 20272 21698 20324
rect 23106 20312 23112 20324
rect 23019 20284 23112 20312
rect 23106 20272 23112 20284
rect 23164 20312 23170 20324
rect 28442 20312 28448 20324
rect 23164 20284 28448 20312
rect 23164 20272 23170 20284
rect 28442 20272 28448 20284
rect 28500 20272 28506 20324
rect 10045 20247 10103 20253
rect 10045 20244 10057 20247
rect 10008 20216 10057 20244
rect 10008 20204 10014 20216
rect 10045 20213 10057 20216
rect 10091 20213 10103 20247
rect 10045 20207 10103 20213
rect 10597 20247 10655 20253
rect 10597 20213 10609 20247
rect 10643 20244 10655 20247
rect 10778 20244 10784 20256
rect 10643 20216 10784 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 10778 20204 10784 20216
rect 10836 20204 10842 20256
rect 12989 20247 13047 20253
rect 12989 20213 13001 20247
rect 13035 20244 13047 20247
rect 13354 20244 13360 20256
rect 13035 20216 13360 20244
rect 13035 20213 13047 20216
rect 12989 20207 13047 20213
rect 13354 20204 13360 20216
rect 13412 20204 13418 20256
rect 14461 20247 14519 20253
rect 14461 20213 14473 20247
rect 14507 20244 14519 20247
rect 14550 20244 14556 20256
rect 14507 20216 14556 20244
rect 14507 20213 14519 20216
rect 14461 20207 14519 20213
rect 14550 20204 14556 20216
rect 14608 20204 14614 20256
rect 17497 20247 17555 20253
rect 17497 20213 17509 20247
rect 17543 20244 17555 20247
rect 17770 20244 17776 20256
rect 17543 20216 17776 20244
rect 17543 20213 17555 20216
rect 17497 20207 17555 20213
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 19242 20244 19248 20256
rect 18104 20216 19248 20244
rect 18104 20204 18110 20216
rect 19242 20204 19248 20216
rect 19300 20244 19306 20256
rect 19337 20247 19395 20253
rect 19337 20244 19349 20247
rect 19300 20216 19349 20244
rect 19300 20204 19306 20216
rect 19337 20213 19349 20216
rect 19383 20213 19395 20247
rect 19337 20207 19395 20213
rect 19886 20204 19892 20256
rect 19944 20244 19950 20256
rect 19981 20247 20039 20253
rect 19981 20244 19993 20247
rect 19944 20216 19993 20244
rect 19944 20204 19950 20216
rect 19981 20213 19993 20216
rect 20027 20213 20039 20247
rect 19981 20207 20039 20213
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 20717 20247 20775 20253
rect 20717 20244 20729 20247
rect 20680 20216 20729 20244
rect 20680 20204 20686 20216
rect 20717 20213 20729 20216
rect 20763 20213 20775 20247
rect 20717 20207 20775 20213
rect 25498 20204 25504 20256
rect 25556 20244 25562 20256
rect 26237 20247 26295 20253
rect 26237 20244 26249 20247
rect 25556 20216 26249 20244
rect 25556 20204 25562 20216
rect 26237 20213 26249 20216
rect 26283 20213 26295 20247
rect 26237 20207 26295 20213
rect 27801 20247 27859 20253
rect 27801 20213 27813 20247
rect 27847 20244 27859 20247
rect 27982 20244 27988 20256
rect 27847 20216 27988 20244
rect 27847 20213 27859 20216
rect 27801 20207 27859 20213
rect 27982 20204 27988 20216
rect 28040 20204 28046 20256
rect 28166 20204 28172 20256
rect 28224 20244 28230 20256
rect 28261 20247 28319 20253
rect 28261 20244 28273 20247
rect 28224 20216 28273 20244
rect 28224 20204 28230 20216
rect 28261 20213 28273 20216
rect 28307 20213 28319 20247
rect 28261 20207 28319 20213
rect 1104 20154 29440 20176
rect 1104 20102 4492 20154
rect 4544 20102 4556 20154
rect 4608 20102 4620 20154
rect 4672 20102 4684 20154
rect 4736 20102 4748 20154
rect 4800 20102 11576 20154
rect 11628 20102 11640 20154
rect 11692 20102 11704 20154
rect 11756 20102 11768 20154
rect 11820 20102 11832 20154
rect 11884 20102 18660 20154
rect 18712 20102 18724 20154
rect 18776 20102 18788 20154
rect 18840 20102 18852 20154
rect 18904 20102 18916 20154
rect 18968 20102 25744 20154
rect 25796 20102 25808 20154
rect 25860 20102 25872 20154
rect 25924 20102 25936 20154
rect 25988 20102 26000 20154
rect 26052 20102 29440 20154
rect 1104 20080 29440 20102
rect 3053 20043 3111 20049
rect 3053 20009 3065 20043
rect 3099 20009 3111 20043
rect 3234 20040 3240 20052
rect 3195 20012 3240 20040
rect 3053 20003 3111 20009
rect 3068 19904 3096 20003
rect 3234 20000 3240 20012
rect 3292 20000 3298 20052
rect 5902 20040 5908 20052
rect 5863 20012 5908 20040
rect 5902 20000 5908 20012
rect 5960 20000 5966 20052
rect 6089 20043 6147 20049
rect 6089 20009 6101 20043
rect 6135 20040 6147 20043
rect 6546 20040 6552 20052
rect 6135 20012 6552 20040
rect 6135 20009 6147 20012
rect 6089 20003 6147 20009
rect 3881 19975 3939 19981
rect 3881 19941 3893 19975
rect 3927 19972 3939 19975
rect 4154 19972 4160 19984
rect 3927 19944 4160 19972
rect 3927 19941 3939 19944
rect 3881 19935 3939 19941
rect 4154 19932 4160 19944
rect 4212 19932 4218 19984
rect 5261 19975 5319 19981
rect 5261 19972 5273 19975
rect 4264 19944 5273 19972
rect 4264 19904 4292 19944
rect 5261 19941 5273 19944
rect 5307 19941 5319 19975
rect 5261 19935 5319 19941
rect 6104 19904 6132 20003
rect 6546 20000 6552 20012
rect 6604 20000 6610 20052
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 8294 20040 8300 20052
rect 7064 20012 8156 20040
rect 8255 20012 8300 20040
rect 7064 20000 7070 20012
rect 6454 19972 6460 19984
rect 6196 19944 6460 19972
rect 6196 19913 6224 19944
rect 6454 19932 6460 19944
rect 6512 19972 6518 19984
rect 7834 19972 7840 19984
rect 6512 19944 7840 19972
rect 6512 19932 6518 19944
rect 7834 19932 7840 19944
rect 7892 19932 7898 19984
rect 8128 19972 8156 20012
rect 8294 20000 8300 20012
rect 8352 20040 8358 20052
rect 9125 20043 9183 20049
rect 9125 20040 9137 20043
rect 8352 20012 9137 20040
rect 8352 20000 8358 20012
rect 9125 20009 9137 20012
rect 9171 20009 9183 20043
rect 9950 20040 9956 20052
rect 9911 20012 9956 20040
rect 9125 20003 9183 20009
rect 9950 20000 9956 20012
rect 10008 20000 10014 20052
rect 12894 20000 12900 20052
rect 12952 20040 12958 20052
rect 13538 20040 13544 20052
rect 12952 20012 13544 20040
rect 12952 20000 12958 20012
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 21913 20043 21971 20049
rect 17052 20012 18552 20040
rect 9582 19972 9588 19984
rect 8128 19944 9588 19972
rect 9582 19932 9588 19944
rect 9640 19972 9646 19984
rect 10597 19975 10655 19981
rect 10597 19972 10609 19975
rect 9640 19944 10609 19972
rect 9640 19932 9646 19944
rect 10597 19941 10609 19944
rect 10643 19941 10655 19975
rect 14642 19972 14648 19984
rect 10597 19935 10655 19941
rect 13280 19944 14648 19972
rect 2240 19876 2820 19904
rect 3068 19876 4292 19904
rect 2240 19848 2268 19876
rect 1670 19836 1676 19848
rect 1631 19808 1676 19836
rect 1670 19796 1676 19808
rect 1728 19796 1734 19848
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19836 2191 19839
rect 2222 19836 2228 19848
rect 2179 19808 2228 19836
rect 2179 19805 2191 19808
rect 2133 19799 2191 19805
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 2317 19839 2375 19845
rect 2317 19805 2329 19839
rect 2363 19836 2375 19839
rect 2682 19836 2688 19848
rect 2363 19808 2688 19836
rect 2363 19805 2375 19808
rect 2317 19799 2375 19805
rect 2682 19796 2688 19808
rect 2740 19796 2746 19848
rect 2792 19845 2820 19876
rect 4264 19848 4292 19876
rect 5276 19876 6132 19904
rect 6181 19907 6239 19913
rect 5276 19848 5304 19876
rect 6181 19873 6193 19907
rect 6227 19873 6239 19907
rect 6181 19867 6239 19873
rect 6472 19876 7328 19904
rect 2777 19839 2835 19845
rect 2777 19805 2789 19839
rect 2823 19805 2835 19839
rect 4062 19836 4068 19848
rect 4023 19808 4068 19836
rect 2777 19799 2835 19805
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 4246 19836 4252 19848
rect 4159 19808 4252 19836
rect 4246 19796 4252 19808
rect 4304 19796 4310 19848
rect 4430 19836 4436 19848
rect 4391 19808 4436 19836
rect 4430 19796 4436 19808
rect 4488 19796 4494 19848
rect 4525 19839 4583 19845
rect 4525 19805 4537 19839
rect 4571 19805 4583 19839
rect 4525 19799 4583 19805
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19805 5043 19839
rect 5258 19836 5264 19848
rect 5219 19808 5264 19836
rect 4985 19799 5043 19805
rect 3694 19728 3700 19780
rect 3752 19768 3758 19780
rect 3878 19768 3884 19780
rect 3752 19740 3884 19768
rect 3752 19728 3758 19740
rect 3878 19728 3884 19740
rect 3936 19768 3942 19780
rect 4157 19771 4215 19777
rect 4157 19768 4169 19771
rect 3936 19740 4169 19768
rect 3936 19728 3942 19740
rect 4157 19737 4169 19740
rect 4203 19737 4215 19771
rect 4157 19731 4215 19737
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 2317 19703 2375 19709
rect 2317 19669 2329 19703
rect 2363 19700 2375 19703
rect 4062 19700 4068 19712
rect 2363 19672 4068 19700
rect 2363 19669 2375 19672
rect 2317 19663 2375 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 4540 19700 4568 19799
rect 5000 19768 5028 19799
rect 5258 19796 5264 19808
rect 5316 19796 5322 19848
rect 5445 19839 5503 19845
rect 5445 19805 5457 19839
rect 5491 19836 5503 19839
rect 6196 19836 6224 19867
rect 6472 19845 6500 19876
rect 5491 19808 6224 19836
rect 6457 19839 6515 19845
rect 5491 19805 5503 19808
rect 5445 19799 5503 19805
rect 6457 19805 6469 19839
rect 6503 19805 6515 19839
rect 7098 19836 7104 19848
rect 7059 19808 7104 19836
rect 6457 19799 6515 19805
rect 6472 19768 6500 19799
rect 7098 19796 7104 19808
rect 7156 19796 7162 19848
rect 7300 19845 7328 19876
rect 9858 19864 9864 19916
rect 9916 19864 9922 19916
rect 13280 19913 13308 19944
rect 14642 19932 14648 19944
rect 14700 19932 14706 19984
rect 13265 19907 13323 19913
rect 13265 19873 13277 19907
rect 13311 19873 13323 19907
rect 13265 19867 13323 19873
rect 13449 19907 13507 19913
rect 13449 19873 13461 19907
rect 13495 19904 13507 19907
rect 13538 19904 13544 19916
rect 13495 19876 13544 19904
rect 13495 19873 13507 19876
rect 13449 19867 13507 19873
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 13906 19864 13912 19916
rect 13964 19904 13970 19916
rect 14458 19904 14464 19916
rect 13964 19876 14464 19904
rect 13964 19864 13970 19876
rect 14458 19864 14464 19876
rect 14516 19904 14522 19916
rect 14516 19876 14687 19904
rect 14516 19864 14522 19876
rect 7193 19839 7251 19845
rect 7193 19805 7205 19839
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19836 7343 19839
rect 7374 19836 7380 19848
rect 7331 19808 7380 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 5000 19740 6500 19768
rect 7006 19728 7012 19780
rect 7064 19768 7070 19780
rect 7208 19768 7236 19799
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 9769 19839 9827 19845
rect 9769 19805 9781 19839
rect 9815 19836 9827 19839
rect 9876 19836 9904 19864
rect 9815 19808 9904 19836
rect 10045 19839 10103 19845
rect 9815 19805 9827 19808
rect 9769 19799 9827 19805
rect 10045 19805 10057 19839
rect 10091 19836 10103 19839
rect 10594 19836 10600 19848
rect 10091 19808 10600 19836
rect 10091 19805 10103 19808
rect 10045 19799 10103 19805
rect 10594 19796 10600 19808
rect 10652 19836 10658 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 10652 19808 10916 19836
rect 10652 19796 10658 19808
rect 7064 19740 7236 19768
rect 7064 19728 7070 19740
rect 7466 19728 7472 19780
rect 7524 19768 7530 19780
rect 9677 19771 9735 19777
rect 9677 19768 9689 19771
rect 7524 19740 9689 19768
rect 7524 19728 7530 19740
rect 9677 19737 9689 19740
rect 9723 19737 9735 19771
rect 9677 19731 9735 19737
rect 9858 19728 9864 19780
rect 9916 19768 9922 19780
rect 10137 19771 10195 19777
rect 10137 19768 10149 19771
rect 9916 19740 10149 19768
rect 9916 19728 9922 19740
rect 10137 19737 10149 19740
rect 10183 19737 10195 19771
rect 10778 19768 10784 19780
rect 10739 19740 10784 19768
rect 10137 19731 10195 19737
rect 10778 19728 10784 19740
rect 10836 19728 10842 19780
rect 10888 19712 10916 19808
rect 12820 19808 14289 19836
rect 10965 19771 11023 19777
rect 10965 19737 10977 19771
rect 11011 19768 11023 19771
rect 11514 19768 11520 19780
rect 11011 19740 11520 19768
rect 11011 19737 11023 19740
rect 10965 19731 11023 19737
rect 11514 19728 11520 19740
rect 11572 19728 11578 19780
rect 4706 19700 4712 19712
rect 4540 19672 4712 19700
rect 4706 19660 4712 19672
rect 4764 19700 4770 19712
rect 5718 19700 5724 19712
rect 4764 19672 5724 19700
rect 4764 19660 4770 19672
rect 5718 19660 5724 19672
rect 5776 19660 5782 19712
rect 6917 19703 6975 19709
rect 6917 19669 6929 19703
rect 6963 19700 6975 19703
rect 7282 19700 7288 19712
rect 6963 19672 7288 19700
rect 6963 19669 6975 19672
rect 6917 19663 6975 19669
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 10870 19660 10876 19712
rect 10928 19700 10934 19712
rect 11977 19703 12035 19709
rect 11977 19700 11989 19703
rect 10928 19672 11989 19700
rect 10928 19660 10934 19672
rect 11977 19669 11989 19672
rect 12023 19669 12035 19703
rect 11977 19663 12035 19669
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 12820 19709 12848 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19805 14427 19839
rect 14550 19836 14556 19848
rect 14511 19808 14556 19836
rect 14369 19799 14427 19805
rect 12894 19728 12900 19780
rect 12952 19768 12958 19780
rect 14384 19768 14412 19799
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 14659 19845 14687 19876
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19805 14703 19839
rect 16114 19836 16120 19848
rect 16027 19808 16120 19836
rect 14645 19799 14703 19805
rect 16114 19796 16120 19808
rect 16172 19836 16178 19848
rect 16945 19839 17003 19845
rect 16945 19836 16957 19839
rect 16172 19808 16957 19836
rect 16172 19796 16178 19808
rect 16945 19805 16957 19808
rect 16991 19836 17003 19839
rect 17052 19836 17080 20012
rect 17678 19932 17684 19984
rect 17736 19972 17742 19984
rect 18417 19975 18475 19981
rect 18417 19972 18429 19975
rect 17736 19944 18429 19972
rect 17736 19932 17742 19944
rect 18417 19941 18429 19944
rect 18463 19941 18475 19975
rect 18524 19972 18552 20012
rect 21913 20009 21925 20043
rect 21959 20040 21971 20043
rect 22738 20040 22744 20052
rect 21959 20012 22744 20040
rect 21959 20009 21971 20012
rect 21913 20003 21971 20009
rect 22738 20000 22744 20012
rect 22796 20040 22802 20052
rect 25590 20040 25596 20052
rect 22796 20012 25596 20040
rect 22796 20000 22802 20012
rect 25590 20000 25596 20012
rect 25648 20000 25654 20052
rect 26145 20043 26203 20049
rect 26145 20009 26157 20043
rect 26191 20040 26203 20043
rect 26234 20040 26240 20052
rect 26191 20012 26240 20040
rect 26191 20009 26203 20012
rect 26145 20003 26203 20009
rect 26234 20000 26240 20012
rect 26292 20000 26298 20052
rect 25498 19972 25504 19984
rect 18524 19944 25504 19972
rect 18417 19935 18475 19941
rect 25498 19932 25504 19944
rect 25556 19972 25562 19984
rect 27249 19975 27307 19981
rect 27249 19972 27261 19975
rect 25556 19944 27261 19972
rect 25556 19932 25562 19944
rect 27249 19941 27261 19944
rect 27295 19972 27307 19975
rect 27798 19972 27804 19984
rect 27295 19944 27804 19972
rect 27295 19941 27307 19944
rect 27249 19935 27307 19941
rect 27798 19932 27804 19944
rect 27856 19932 27862 19984
rect 17221 19907 17279 19913
rect 17221 19873 17233 19907
rect 17267 19904 17279 19907
rect 17770 19904 17776 19916
rect 17267 19876 17776 19904
rect 17267 19873 17279 19876
rect 17221 19867 17279 19873
rect 17770 19864 17776 19876
rect 17828 19864 17834 19916
rect 18138 19864 18144 19916
rect 18196 19904 18202 19916
rect 18509 19907 18567 19913
rect 18509 19904 18521 19907
rect 18196 19876 18521 19904
rect 18196 19864 18202 19876
rect 18509 19873 18521 19876
rect 18555 19904 18567 19907
rect 19242 19904 19248 19916
rect 18555 19876 19248 19904
rect 18555 19873 18567 19876
rect 18509 19867 18567 19873
rect 19242 19864 19248 19876
rect 19300 19864 19306 19916
rect 20714 19864 20720 19916
rect 20772 19904 20778 19916
rect 21085 19907 21143 19913
rect 21085 19904 21097 19907
rect 20772 19876 21097 19904
rect 20772 19864 20778 19876
rect 21085 19873 21097 19876
rect 21131 19873 21143 19907
rect 23014 19904 23020 19916
rect 21085 19867 21143 19873
rect 22572 19876 23020 19904
rect 18340 19845 18460 19846
rect 16991 19808 17080 19836
rect 18293 19839 18460 19845
rect 16991 19805 17003 19808
rect 16945 19799 17003 19805
rect 18293 19805 18305 19839
rect 18339 19818 18460 19839
rect 18339 19808 18368 19818
rect 18339 19805 18351 19808
rect 18293 19799 18351 19805
rect 17037 19771 17095 19777
rect 17037 19768 17049 19771
rect 12952 19740 14412 19768
rect 15580 19740 17049 19768
rect 12952 19728 12958 19740
rect 15580 19712 15608 19740
rect 17037 19737 17049 19740
rect 17083 19768 17095 19771
rect 17310 19768 17316 19780
rect 17083 19740 17316 19768
rect 17083 19737 17095 19740
rect 17037 19731 17095 19737
rect 17310 19728 17316 19740
rect 17368 19728 17374 19780
rect 18432 19768 18460 19818
rect 18598 19796 18604 19848
rect 18656 19836 18662 19848
rect 20257 19839 20315 19845
rect 18656 19808 18701 19836
rect 18656 19796 18662 19808
rect 20257 19805 20269 19839
rect 20303 19836 20315 19839
rect 20622 19836 20628 19848
rect 20303 19808 20628 19836
rect 20303 19805 20315 19808
rect 20257 19799 20315 19805
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 20990 19836 20996 19848
rect 20951 19808 20996 19836
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 21269 19839 21327 19845
rect 21269 19805 21281 19839
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 21361 19839 21419 19845
rect 21361 19805 21373 19839
rect 21407 19836 21419 19839
rect 21818 19836 21824 19848
rect 21407 19808 21824 19836
rect 21407 19805 21419 19808
rect 21361 19799 21419 19805
rect 20530 19768 20536 19780
rect 18432 19740 20536 19768
rect 20530 19728 20536 19740
rect 20588 19728 20594 19780
rect 20640 19768 20668 19796
rect 21284 19768 21312 19799
rect 21818 19796 21824 19808
rect 21876 19796 21882 19848
rect 22572 19836 22600 19876
rect 23014 19864 23020 19876
rect 23072 19864 23078 19916
rect 22649 19839 22707 19845
rect 22649 19836 22661 19839
rect 22572 19808 22661 19836
rect 22649 19805 22661 19808
rect 22695 19805 22707 19839
rect 22649 19799 22707 19805
rect 22738 19796 22744 19848
rect 22796 19836 22802 19848
rect 22796 19808 22841 19836
rect 22796 19796 22802 19808
rect 23106 19796 23112 19848
rect 23164 19836 23170 19848
rect 23845 19839 23903 19845
rect 23845 19836 23857 19839
rect 23164 19808 23857 19836
rect 23164 19796 23170 19808
rect 23845 19805 23857 19808
rect 23891 19836 23903 19839
rect 24857 19839 24915 19845
rect 24857 19836 24869 19839
rect 23891 19808 24869 19836
rect 23891 19805 23903 19808
rect 23845 19799 23903 19805
rect 24857 19805 24869 19808
rect 24903 19805 24915 19839
rect 24857 19799 24915 19805
rect 25501 19839 25559 19845
rect 25501 19805 25513 19839
rect 25547 19805 25559 19839
rect 27982 19836 27988 19848
rect 27943 19808 27988 19836
rect 25501 19799 25559 19805
rect 20640 19740 21312 19768
rect 24762 19728 24768 19780
rect 24820 19768 24826 19780
rect 25516 19768 25544 19799
rect 27982 19796 27988 19808
rect 28040 19796 28046 19848
rect 24820 19740 25544 19768
rect 24820 19728 24826 19740
rect 12805 19703 12863 19709
rect 12805 19700 12817 19703
rect 12768 19672 12817 19700
rect 12768 19660 12774 19672
rect 12805 19669 12817 19672
rect 12851 19669 12863 19703
rect 12805 19663 12863 19669
rect 13173 19703 13231 19709
rect 13173 19669 13185 19703
rect 13219 19700 13231 19703
rect 13354 19700 13360 19712
rect 13219 19672 13360 19700
rect 13219 19669 13231 19672
rect 13173 19663 13231 19669
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 14093 19703 14151 19709
rect 14093 19700 14105 19703
rect 13872 19672 14105 19700
rect 13872 19660 13878 19672
rect 14093 19669 14105 19672
rect 14139 19669 14151 19703
rect 15562 19700 15568 19712
rect 15523 19672 15568 19700
rect 14093 19663 14151 19669
rect 15562 19660 15568 19672
rect 15620 19660 15626 19712
rect 16577 19703 16635 19709
rect 16577 19669 16589 19703
rect 16623 19700 16635 19703
rect 16666 19700 16672 19712
rect 16623 19672 16672 19700
rect 16623 19669 16635 19672
rect 16577 19663 16635 19669
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 18138 19700 18144 19712
rect 18099 19672 18144 19700
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 20346 19660 20352 19712
rect 20404 19700 20410 19712
rect 20901 19703 20959 19709
rect 20901 19700 20913 19703
rect 20404 19672 20913 19700
rect 20404 19660 20410 19672
rect 20901 19669 20913 19672
rect 20947 19669 20959 19703
rect 20901 19663 20959 19669
rect 22465 19703 22523 19709
rect 22465 19669 22477 19703
rect 22511 19700 22523 19703
rect 22830 19700 22836 19712
rect 22511 19672 22836 19700
rect 22511 19669 22523 19672
rect 22465 19663 22523 19669
rect 22830 19660 22836 19672
rect 22888 19660 22894 19712
rect 28166 19700 28172 19712
rect 28127 19672 28172 19700
rect 28166 19660 28172 19672
rect 28224 19660 28230 19712
rect 1104 19610 29600 19632
rect 1104 19558 8034 19610
rect 8086 19558 8098 19610
rect 8150 19558 8162 19610
rect 8214 19558 8226 19610
rect 8278 19558 8290 19610
rect 8342 19558 15118 19610
rect 15170 19558 15182 19610
rect 15234 19558 15246 19610
rect 15298 19558 15310 19610
rect 15362 19558 15374 19610
rect 15426 19558 22202 19610
rect 22254 19558 22266 19610
rect 22318 19558 22330 19610
rect 22382 19558 22394 19610
rect 22446 19558 22458 19610
rect 22510 19558 29286 19610
rect 29338 19558 29350 19610
rect 29402 19558 29414 19610
rect 29466 19558 29478 19610
rect 29530 19558 29542 19610
rect 29594 19558 29600 19610
rect 1104 19536 29600 19558
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 3142 19496 3148 19508
rect 2832 19468 3148 19496
rect 2832 19456 2838 19468
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 4058 19499 4116 19505
rect 4058 19465 4070 19499
rect 4104 19496 4116 19499
rect 4430 19496 4436 19508
rect 4104 19468 4436 19496
rect 4104 19465 4116 19468
rect 4058 19459 4116 19465
rect 4430 19456 4436 19468
rect 4488 19456 4494 19508
rect 4706 19496 4712 19508
rect 4667 19468 4712 19496
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 5258 19496 5264 19508
rect 5219 19468 5264 19496
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 6809 19499 6867 19505
rect 6809 19465 6821 19499
rect 6855 19496 6867 19499
rect 6914 19496 6920 19508
rect 6855 19468 6920 19496
rect 6855 19465 6867 19468
rect 6809 19459 6867 19465
rect 6914 19456 6920 19468
rect 6972 19456 6978 19508
rect 10042 19496 10048 19508
rect 10003 19468 10048 19496
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 10229 19499 10287 19505
rect 10229 19465 10241 19499
rect 10275 19496 10287 19499
rect 12066 19496 12072 19508
rect 10275 19468 12072 19496
rect 10275 19465 10287 19468
rect 10229 19459 10287 19465
rect 12066 19456 12072 19468
rect 12124 19456 12130 19508
rect 16114 19496 16120 19508
rect 12406 19468 16120 19496
rect 2406 19428 2412 19440
rect 2367 19400 2412 19428
rect 2406 19388 2412 19400
rect 2464 19388 2470 19440
rect 3973 19431 4031 19437
rect 3973 19397 3985 19431
rect 4019 19428 4031 19431
rect 4246 19428 4252 19440
rect 4019 19400 4252 19428
rect 4019 19397 4031 19400
rect 3973 19391 4031 19397
rect 4246 19388 4252 19400
rect 4304 19388 4310 19440
rect 7009 19431 7067 19437
rect 7009 19397 7021 19431
rect 7055 19428 7067 19431
rect 7650 19428 7656 19440
rect 7055 19400 7656 19428
rect 7055 19397 7067 19400
rect 7009 19391 7067 19397
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 2314 19360 2320 19372
rect 2275 19332 2320 19360
rect 2314 19320 2320 19332
rect 2372 19320 2378 19372
rect 2498 19320 2504 19372
rect 2556 19360 2562 19372
rect 2593 19363 2651 19369
rect 2593 19360 2605 19363
rect 2556 19332 2605 19360
rect 2556 19320 2562 19332
rect 2593 19329 2605 19332
rect 2639 19329 2651 19363
rect 3878 19360 3884 19372
rect 3791 19332 3884 19360
rect 2593 19323 2651 19329
rect 3878 19320 3884 19332
rect 3936 19360 3942 19372
rect 3936 19332 4016 19360
rect 3936 19320 3942 19332
rect 3988 19292 4016 19332
rect 4062 19320 4068 19372
rect 4120 19360 4126 19372
rect 4157 19363 4215 19369
rect 4157 19360 4169 19363
rect 4120 19332 4169 19360
rect 4120 19320 4126 19332
rect 4157 19329 4169 19332
rect 4203 19329 4215 19363
rect 5902 19360 5908 19372
rect 4157 19323 4215 19329
rect 4264 19332 5908 19360
rect 4264 19292 4292 19332
rect 5902 19320 5908 19332
rect 5960 19320 5966 19372
rect 3988 19264 4292 19292
rect 5813 19295 5871 19301
rect 5813 19261 5825 19295
rect 5859 19292 5871 19295
rect 7024 19292 7052 19391
rect 7650 19388 7656 19400
rect 7708 19388 7714 19440
rect 9122 19428 9128 19440
rect 9083 19400 9128 19428
rect 9122 19388 9128 19400
rect 9180 19388 9186 19440
rect 9398 19388 9404 19440
rect 9456 19428 9462 19440
rect 10060 19428 10088 19456
rect 10689 19431 10747 19437
rect 10689 19428 10701 19431
rect 9456 19400 9996 19428
rect 10060 19400 10701 19428
rect 9456 19388 9462 19400
rect 8941 19363 8999 19369
rect 8941 19329 8953 19363
rect 8987 19360 8999 19363
rect 9490 19360 9496 19372
rect 8987 19332 9496 19360
rect 8987 19329 8999 19332
rect 8941 19323 8999 19329
rect 9490 19320 9496 19332
rect 9548 19360 9554 19372
rect 9585 19363 9643 19369
rect 9585 19360 9597 19363
rect 9548 19332 9597 19360
rect 9548 19320 9554 19332
rect 9585 19329 9597 19332
rect 9631 19329 9643 19363
rect 9585 19323 9643 19329
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 9858 19360 9864 19372
rect 9723 19332 9864 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 9968 19360 9996 19400
rect 10689 19397 10701 19400
rect 10735 19397 10747 19431
rect 10689 19391 10747 19397
rect 10048 19363 10106 19369
rect 10048 19360 10060 19363
rect 9968 19332 10060 19360
rect 10048 19329 10060 19332
rect 10094 19360 10106 19363
rect 12406 19360 12434 19468
rect 16114 19456 16120 19468
rect 16172 19456 16178 19508
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19496 16911 19499
rect 17034 19496 17040 19508
rect 16899 19468 17040 19496
rect 16899 19465 16911 19468
rect 16853 19459 16911 19465
rect 17034 19456 17040 19468
rect 17092 19456 17098 19508
rect 17310 19496 17316 19508
rect 17271 19468 17316 19496
rect 17310 19456 17316 19468
rect 17368 19456 17374 19508
rect 19889 19499 19947 19505
rect 19889 19465 19901 19499
rect 19935 19465 19947 19499
rect 20346 19496 20352 19508
rect 20307 19468 20352 19496
rect 19889 19459 19947 19465
rect 18138 19428 18144 19440
rect 14016 19400 18144 19428
rect 13814 19360 13820 19372
rect 10094 19332 12434 19360
rect 13775 19332 13820 19360
rect 10094 19329 10106 19332
rect 10048 19323 10106 19329
rect 13814 19320 13820 19332
rect 13872 19320 13878 19372
rect 14016 19369 14044 19400
rect 18138 19388 18144 19400
rect 18196 19388 18202 19440
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19329 14059 19363
rect 14001 19323 14059 19329
rect 14642 19320 14648 19372
rect 14700 19360 14706 19372
rect 16666 19360 16672 19372
rect 14700 19332 16528 19360
rect 16627 19332 16672 19360
rect 14700 19320 14706 19332
rect 7098 19292 7104 19304
rect 5859 19264 7104 19292
rect 5859 19261 5871 19264
rect 5813 19255 5871 19261
rect 7098 19252 7104 19264
rect 7156 19252 7162 19304
rect 7374 19252 7380 19304
rect 7432 19292 7438 19304
rect 8757 19295 8815 19301
rect 8757 19292 8769 19295
rect 7432 19264 8769 19292
rect 7432 19252 7438 19264
rect 8757 19261 8769 19264
rect 8803 19261 8815 19295
rect 16500 19292 16528 19332
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 16850 19360 16856 19372
rect 16811 19332 16856 19360
rect 16850 19320 16856 19332
rect 16908 19320 16914 19372
rect 19904 19360 19932 19459
rect 20346 19456 20352 19468
rect 20404 19456 20410 19508
rect 27798 19496 27804 19508
rect 27759 19468 27804 19496
rect 27798 19456 27804 19468
rect 27856 19456 27862 19508
rect 20257 19431 20315 19437
rect 20257 19397 20269 19431
rect 20303 19428 20315 19431
rect 20438 19428 20444 19440
rect 20303 19400 20444 19428
rect 20303 19397 20315 19400
rect 20257 19391 20315 19397
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 23474 19428 23480 19440
rect 23435 19400 23480 19428
rect 23474 19388 23480 19400
rect 23532 19388 23538 19440
rect 16960 19332 19932 19360
rect 16960 19292 16988 19332
rect 19978 19320 19984 19372
rect 20036 19360 20042 19372
rect 23106 19360 23112 19372
rect 20036 19332 23112 19360
rect 20036 19320 20042 19332
rect 23106 19320 23112 19332
rect 23164 19320 23170 19372
rect 23198 19320 23204 19372
rect 23256 19360 23262 19372
rect 23293 19363 23351 19369
rect 23293 19360 23305 19363
rect 23256 19332 23305 19360
rect 23256 19320 23262 19332
rect 23293 19329 23305 19332
rect 23339 19329 23351 19363
rect 24578 19360 24584 19372
rect 24539 19332 24584 19360
rect 23293 19323 23351 19329
rect 16500 19264 16988 19292
rect 17957 19295 18015 19301
rect 8757 19255 8815 19261
rect 17957 19261 17969 19295
rect 18003 19292 18015 19295
rect 18046 19292 18052 19304
rect 18003 19264 18052 19292
rect 18003 19261 18015 19264
rect 17957 19255 18015 19261
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 20441 19295 20499 19301
rect 20441 19292 20453 19295
rect 19352 19264 20453 19292
rect 1946 19184 1952 19236
rect 2004 19224 2010 19236
rect 2004 19196 7604 19224
rect 2004 19184 2010 19196
rect 1765 19159 1823 19165
rect 1765 19125 1777 19159
rect 1811 19156 1823 19159
rect 2314 19156 2320 19168
rect 1811 19128 2320 19156
rect 1811 19125 1823 19128
rect 1765 19119 1823 19125
rect 2314 19116 2320 19128
rect 2372 19116 2378 19168
rect 2406 19116 2412 19168
rect 2464 19156 2470 19168
rect 3237 19159 3295 19165
rect 3237 19156 3249 19159
rect 2464 19128 3249 19156
rect 2464 19116 2470 19128
rect 3237 19125 3249 19128
rect 3283 19125 3295 19159
rect 3237 19119 3295 19125
rect 6178 19116 6184 19168
rect 6236 19156 6242 19168
rect 6641 19159 6699 19165
rect 6641 19156 6653 19159
rect 6236 19128 6653 19156
rect 6236 19116 6242 19128
rect 6641 19125 6653 19128
rect 6687 19125 6699 19159
rect 6641 19119 6699 19125
rect 6825 19159 6883 19165
rect 6825 19125 6837 19159
rect 6871 19156 6883 19159
rect 7282 19156 7288 19168
rect 6871 19128 7288 19156
rect 6871 19125 6883 19128
rect 6825 19119 6883 19125
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 7576 19165 7604 19196
rect 10226 19184 10232 19236
rect 10284 19224 10290 19236
rect 10284 19196 12434 19224
rect 10284 19184 10290 19196
rect 7561 19159 7619 19165
rect 7561 19125 7573 19159
rect 7607 19156 7619 19159
rect 7650 19156 7656 19168
rect 7607 19128 7656 19156
rect 7607 19125 7619 19128
rect 7561 19119 7619 19125
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 7926 19116 7932 19168
rect 7984 19156 7990 19168
rect 8202 19156 8208 19168
rect 7984 19128 8208 19156
rect 7984 19116 7990 19128
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 12406 19156 12434 19196
rect 13906 19156 13912 19168
rect 12406 19128 13912 19156
rect 13906 19116 13912 19128
rect 13964 19116 13970 19168
rect 16022 19116 16028 19168
rect 16080 19156 16086 19168
rect 16117 19159 16175 19165
rect 16117 19156 16129 19159
rect 16080 19128 16129 19156
rect 16080 19116 16086 19128
rect 16117 19125 16129 19128
rect 16163 19156 16175 19159
rect 16298 19156 16304 19168
rect 16163 19128 16304 19156
rect 16163 19125 16175 19128
rect 16117 19119 16175 19125
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 16574 19116 16580 19168
rect 16632 19156 16638 19168
rect 16758 19156 16764 19168
rect 16632 19128 16764 19156
rect 16632 19116 16638 19128
rect 16758 19116 16764 19128
rect 16816 19156 16822 19168
rect 19352 19165 19380 19264
rect 20441 19261 20453 19264
rect 20487 19261 20499 19295
rect 20441 19255 20499 19261
rect 20530 19252 20536 19304
rect 20588 19292 20594 19304
rect 23308 19292 23336 19323
rect 24578 19320 24584 19332
rect 24636 19320 24642 19372
rect 28166 19360 28172 19372
rect 27908 19332 28172 19360
rect 23937 19295 23995 19301
rect 23937 19292 23949 19295
rect 20588 19264 22094 19292
rect 23308 19264 23949 19292
rect 20588 19252 20594 19264
rect 19337 19159 19395 19165
rect 19337 19156 19349 19159
rect 16816 19128 19349 19156
rect 16816 19116 16822 19128
rect 19337 19125 19349 19128
rect 19383 19125 19395 19159
rect 19337 19119 19395 19125
rect 21269 19159 21327 19165
rect 21269 19125 21281 19159
rect 21315 19156 21327 19159
rect 21358 19156 21364 19168
rect 21315 19128 21364 19156
rect 21315 19125 21327 19128
rect 21269 19119 21327 19125
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 22066 19156 22094 19264
rect 23937 19261 23949 19264
rect 23983 19261 23995 19295
rect 24762 19292 24768 19304
rect 24723 19264 24768 19292
rect 23937 19255 23995 19261
rect 24762 19252 24768 19264
rect 24820 19252 24826 19304
rect 26326 19292 26332 19304
rect 26287 19264 26332 19292
rect 26326 19252 26332 19264
rect 26384 19292 26390 19304
rect 27706 19292 27712 19304
rect 26384 19264 27712 19292
rect 26384 19252 26390 19264
rect 27706 19252 27712 19264
rect 27764 19292 27770 19304
rect 27908 19301 27936 19332
rect 28166 19320 28172 19332
rect 28224 19320 28230 19372
rect 27893 19295 27951 19301
rect 27893 19292 27905 19295
rect 27764 19264 27905 19292
rect 27764 19252 27770 19264
rect 27893 19261 27905 19264
rect 27939 19261 27951 19295
rect 28074 19292 28080 19304
rect 28035 19264 28080 19292
rect 27893 19255 27951 19261
rect 28074 19252 28080 19264
rect 28132 19252 28138 19304
rect 23106 19156 23112 19168
rect 22066 19128 23112 19156
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 27430 19156 27436 19168
rect 27391 19128 27436 19156
rect 27430 19116 27436 19128
rect 27488 19116 27494 19168
rect 28166 19116 28172 19168
rect 28224 19156 28230 19168
rect 28442 19156 28448 19168
rect 28224 19128 28448 19156
rect 28224 19116 28230 19128
rect 28442 19116 28448 19128
rect 28500 19156 28506 19168
rect 28629 19159 28687 19165
rect 28629 19156 28641 19159
rect 28500 19128 28641 19156
rect 28500 19116 28506 19128
rect 28629 19125 28641 19128
rect 28675 19125 28687 19159
rect 28629 19119 28687 19125
rect 1104 19066 29440 19088
rect 1104 19014 4492 19066
rect 4544 19014 4556 19066
rect 4608 19014 4620 19066
rect 4672 19014 4684 19066
rect 4736 19014 4748 19066
rect 4800 19014 11576 19066
rect 11628 19014 11640 19066
rect 11692 19014 11704 19066
rect 11756 19014 11768 19066
rect 11820 19014 11832 19066
rect 11884 19014 18660 19066
rect 18712 19014 18724 19066
rect 18776 19014 18788 19066
rect 18840 19014 18852 19066
rect 18904 19014 18916 19066
rect 18968 19014 25744 19066
rect 25796 19014 25808 19066
rect 25860 19014 25872 19066
rect 25924 19014 25936 19066
rect 25988 19014 26000 19066
rect 26052 19014 29440 19066
rect 1104 18992 29440 19014
rect 2222 18952 2228 18964
rect 2183 18924 2228 18952
rect 2222 18912 2228 18924
rect 2280 18912 2286 18964
rect 4709 18955 4767 18961
rect 4709 18921 4721 18955
rect 4755 18952 4767 18955
rect 5350 18952 5356 18964
rect 4755 18924 5356 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 5350 18912 5356 18924
rect 5408 18912 5414 18964
rect 7193 18955 7251 18961
rect 7193 18921 7205 18955
rect 7239 18952 7251 18955
rect 7466 18952 7472 18964
rect 7239 18924 7472 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 7466 18912 7472 18924
rect 7524 18912 7530 18964
rect 7837 18955 7895 18961
rect 7837 18921 7849 18955
rect 7883 18952 7895 18955
rect 8386 18952 8392 18964
rect 7883 18924 8392 18952
rect 7883 18921 7895 18924
rect 7837 18915 7895 18921
rect 5169 18887 5227 18893
rect 5169 18884 5181 18887
rect 2424 18856 5181 18884
rect 2424 18828 2452 18856
rect 5169 18853 5181 18856
rect 5215 18853 5227 18887
rect 5169 18847 5227 18853
rect 2406 18816 2412 18828
rect 2240 18788 2412 18816
rect 2240 18757 2268 18788
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 2225 18751 2283 18757
rect 2225 18748 2237 18751
rect 1688 18720 2237 18748
rect 1486 18572 1492 18624
rect 1544 18612 1550 18624
rect 1688 18621 1716 18720
rect 2225 18717 2237 18720
rect 2271 18717 2283 18751
rect 2225 18711 2283 18717
rect 2314 18708 2320 18760
rect 2372 18748 2378 18760
rect 2372 18720 2417 18748
rect 2372 18708 2378 18720
rect 2498 18680 2504 18692
rect 2459 18652 2504 18680
rect 2498 18640 2504 18652
rect 2556 18640 2562 18692
rect 2590 18640 2596 18692
rect 2648 18680 2654 18692
rect 5184 18680 5212 18847
rect 5368 18816 5396 18912
rect 5534 18844 5540 18896
rect 5592 18884 5598 18896
rect 7742 18884 7748 18896
rect 5592 18856 7748 18884
rect 5592 18844 5598 18856
rect 7742 18844 7748 18856
rect 7800 18844 7806 18896
rect 5626 18816 5632 18828
rect 5368 18788 5632 18816
rect 5626 18776 5632 18788
rect 5684 18816 5690 18828
rect 7852 18816 7880 18915
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 9490 18952 9496 18964
rect 9451 18924 9496 18952
rect 9490 18912 9496 18924
rect 9548 18912 9554 18964
rect 9766 18912 9772 18964
rect 9824 18952 9830 18964
rect 10229 18955 10287 18961
rect 10229 18952 10241 18955
rect 9824 18924 10241 18952
rect 9824 18912 9830 18924
rect 10229 18921 10241 18924
rect 10275 18921 10287 18955
rect 15470 18952 15476 18964
rect 15431 18924 15476 18952
rect 10229 18915 10287 18921
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 17862 18952 17868 18964
rect 17823 18924 17868 18952
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 21637 18955 21695 18961
rect 21637 18952 21649 18955
rect 20772 18924 21649 18952
rect 20772 18912 20778 18924
rect 21637 18921 21649 18924
rect 21683 18952 21695 18955
rect 21726 18952 21732 18964
rect 21683 18924 21732 18952
rect 21683 18921 21695 18924
rect 21637 18915 21695 18921
rect 21726 18912 21732 18924
rect 21784 18912 21790 18964
rect 23658 18912 23664 18964
rect 23716 18952 23722 18964
rect 23845 18955 23903 18961
rect 23845 18952 23857 18955
rect 23716 18924 23857 18952
rect 23716 18912 23722 18924
rect 23845 18921 23857 18924
rect 23891 18952 23903 18955
rect 24670 18952 24676 18964
rect 23891 18924 24676 18952
rect 23891 18921 23903 18924
rect 23845 18915 23903 18921
rect 24670 18912 24676 18924
rect 24728 18912 24734 18964
rect 27982 18912 27988 18964
rect 28040 18952 28046 18964
rect 28537 18955 28595 18961
rect 28537 18952 28549 18955
rect 28040 18924 28549 18952
rect 28040 18912 28046 18924
rect 28537 18921 28549 18924
rect 28583 18921 28595 18955
rect 28537 18915 28595 18921
rect 16298 18844 16304 18896
rect 16356 18884 16362 18896
rect 16356 18856 17172 18884
rect 16356 18844 16362 18856
rect 5684 18788 6040 18816
rect 5684 18776 5690 18788
rect 5902 18748 5908 18760
rect 5863 18720 5908 18748
rect 5902 18708 5908 18720
rect 5960 18708 5966 18760
rect 6012 18757 6040 18788
rect 7116 18788 7880 18816
rect 5997 18751 6055 18757
rect 5997 18717 6009 18751
rect 6043 18717 6055 18751
rect 6178 18748 6184 18760
rect 6139 18720 6184 18748
rect 5997 18711 6055 18717
rect 6178 18708 6184 18720
rect 6236 18708 6242 18760
rect 6273 18751 6331 18757
rect 6273 18717 6285 18751
rect 6319 18748 6331 18751
rect 7006 18748 7012 18760
rect 6319 18720 7012 18748
rect 6319 18717 6331 18720
rect 6273 18711 6331 18717
rect 7006 18708 7012 18720
rect 7064 18708 7070 18760
rect 7116 18757 7144 18788
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 15562 18816 15568 18828
rect 8628 18788 15568 18816
rect 8628 18776 8634 18788
rect 15562 18776 15568 18788
rect 15620 18776 15626 18828
rect 16117 18819 16175 18825
rect 16117 18785 16129 18819
rect 16163 18816 16175 18819
rect 16758 18816 16764 18828
rect 16163 18788 16764 18816
rect 16163 18785 16175 18788
rect 16117 18779 16175 18785
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 17144 18825 17172 18856
rect 21082 18844 21088 18896
rect 21140 18884 21146 18896
rect 28074 18884 28080 18896
rect 21140 18856 28080 18884
rect 21140 18844 21146 18856
rect 17129 18819 17187 18825
rect 17129 18785 17141 18819
rect 17175 18785 17187 18819
rect 17129 18779 17187 18785
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18816 17371 18819
rect 17770 18816 17776 18828
rect 17359 18788 17776 18816
rect 17359 18785 17371 18788
rect 17313 18779 17371 18785
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 18104 18788 18429 18816
rect 18104 18776 18110 18788
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 20714 18776 20720 18828
rect 20772 18816 20778 18828
rect 20993 18819 21051 18825
rect 20993 18816 21005 18819
rect 20772 18788 21005 18816
rect 20772 18776 20778 18788
rect 20993 18785 21005 18788
rect 21039 18785 21051 18819
rect 20993 18779 21051 18785
rect 23474 18776 23480 18828
rect 23532 18816 23538 18828
rect 23532 18788 24624 18816
rect 23532 18776 23538 18788
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18717 7159 18751
rect 7101 18711 7159 18717
rect 7285 18751 7343 18757
rect 7285 18717 7297 18751
rect 7331 18748 7343 18751
rect 8202 18748 8208 18760
rect 7331 18720 8208 18748
rect 7331 18717 7343 18720
rect 7285 18711 7343 18717
rect 7300 18680 7328 18711
rect 8202 18708 8208 18720
rect 8260 18748 8266 18760
rect 8297 18751 8355 18757
rect 8297 18748 8309 18751
rect 8260 18720 8309 18748
rect 8260 18708 8266 18720
rect 8297 18717 8309 18720
rect 8343 18748 8355 18751
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 8343 18720 9321 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 9309 18717 9321 18720
rect 9355 18717 9367 18751
rect 9490 18748 9496 18760
rect 9451 18720 9496 18748
rect 9309 18711 9367 18717
rect 9490 18708 9496 18720
rect 9548 18708 9554 18760
rect 14093 18751 14151 18757
rect 14093 18717 14105 18751
rect 14139 18717 14151 18751
rect 14093 18711 14151 18717
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18748 14335 18751
rect 14323 18720 15516 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 14108 18680 14136 18711
rect 14182 18680 14188 18692
rect 2648 18652 2774 18680
rect 5184 18652 7328 18680
rect 14095 18652 14188 18680
rect 2648 18640 2654 18652
rect 1673 18615 1731 18621
rect 1673 18612 1685 18615
rect 1544 18584 1685 18612
rect 1544 18572 1550 18584
rect 1673 18581 1685 18584
rect 1719 18581 1731 18615
rect 2746 18612 2774 18652
rect 14182 18640 14188 18652
rect 14240 18680 14246 18692
rect 15010 18680 15016 18692
rect 14240 18652 15016 18680
rect 14240 18640 14246 18652
rect 15010 18640 15016 18652
rect 15068 18640 15074 18692
rect 5534 18612 5540 18624
rect 2746 18584 5540 18612
rect 1673 18575 1731 18581
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 5718 18612 5724 18624
rect 5679 18584 5724 18612
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 14090 18612 14096 18624
rect 14051 18584 14096 18612
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 15488 18612 15516 18720
rect 15580 18680 15608 18776
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 17034 18748 17040 18760
rect 15979 18720 17040 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 17034 18708 17040 18720
rect 17092 18708 17098 18760
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18748 19763 18751
rect 20625 18751 20683 18757
rect 20625 18748 20637 18751
rect 19751 18720 20637 18748
rect 19751 18717 19763 18720
rect 19705 18711 19763 18717
rect 20625 18717 20637 18720
rect 20671 18748 20683 18751
rect 20806 18748 20812 18760
rect 20671 18720 20812 18748
rect 20671 18717 20683 18720
rect 20625 18711 20683 18717
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 19886 18680 19892 18692
rect 15580 18652 17080 18680
rect 19847 18652 19892 18680
rect 15562 18612 15568 18624
rect 15488 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 15838 18612 15844 18624
rect 15799 18584 15844 18612
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 16669 18615 16727 18621
rect 16669 18581 16681 18615
rect 16715 18612 16727 18615
rect 16850 18612 16856 18624
rect 16715 18584 16856 18612
rect 16715 18581 16727 18584
rect 16669 18575 16727 18581
rect 16850 18572 16856 18584
rect 16908 18572 16914 18624
rect 17052 18621 17080 18652
rect 19886 18640 19892 18652
rect 19944 18640 19950 18692
rect 20717 18683 20775 18689
rect 20717 18649 20729 18683
rect 20763 18680 20775 18683
rect 21100 18680 21128 18711
rect 21450 18708 21456 18760
rect 21508 18748 21514 18760
rect 21821 18751 21879 18757
rect 21821 18748 21833 18751
rect 21508 18720 21833 18748
rect 21508 18708 21514 18720
rect 21821 18717 21833 18720
rect 21867 18717 21879 18751
rect 21821 18711 21879 18717
rect 23198 18708 23204 18760
rect 23256 18748 23262 18760
rect 24596 18757 24624 18788
rect 26234 18776 26240 18828
rect 26292 18816 26298 18828
rect 27908 18825 27936 18856
rect 28074 18844 28080 18856
rect 28132 18844 28138 18896
rect 26697 18819 26755 18825
rect 26697 18816 26709 18819
rect 26292 18788 26709 18816
rect 26292 18776 26298 18788
rect 26697 18785 26709 18788
rect 26743 18785 26755 18819
rect 26697 18779 26755 18785
rect 27893 18819 27951 18825
rect 27893 18785 27905 18819
rect 27939 18785 27951 18819
rect 27893 18779 27951 18785
rect 24397 18751 24455 18757
rect 24397 18748 24409 18751
rect 23256 18720 24409 18748
rect 23256 18708 23262 18720
rect 24397 18717 24409 18720
rect 24443 18717 24455 18751
rect 24397 18711 24455 18717
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 26142 18708 26148 18760
rect 26200 18748 26206 18760
rect 26513 18751 26571 18757
rect 26513 18748 26525 18751
rect 26200 18720 26525 18748
rect 26200 18708 26206 18720
rect 26513 18717 26525 18720
rect 26559 18717 26571 18751
rect 27706 18748 27712 18760
rect 27667 18720 27712 18748
rect 26513 18711 26571 18717
rect 27706 18708 27712 18720
rect 27764 18708 27770 18760
rect 28718 18748 28724 18760
rect 28679 18720 28724 18748
rect 28718 18708 28724 18720
rect 28776 18708 28782 18760
rect 21358 18680 21364 18692
rect 20763 18652 21036 18680
rect 21100 18652 21364 18680
rect 20763 18649 20775 18652
rect 20717 18643 20775 18649
rect 21008 18624 21036 18652
rect 21358 18640 21364 18652
rect 21416 18680 21422 18692
rect 21416 18652 21864 18680
rect 21416 18640 21422 18652
rect 21836 18624 21864 18652
rect 17037 18615 17095 18621
rect 17037 18581 17049 18615
rect 17083 18581 17095 18615
rect 18230 18612 18236 18624
rect 18191 18584 18236 18612
rect 17037 18575 17095 18581
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 18322 18572 18328 18624
rect 18380 18612 18386 18624
rect 18380 18584 18425 18612
rect 18380 18572 18386 18584
rect 19426 18572 19432 18624
rect 19484 18612 19490 18624
rect 19521 18615 19579 18621
rect 19521 18612 19533 18615
rect 19484 18584 19533 18612
rect 19484 18572 19490 18584
rect 19521 18581 19533 18584
rect 19567 18581 19579 18615
rect 20346 18612 20352 18624
rect 20307 18584 20352 18612
rect 19521 18575 19579 18581
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 20809 18615 20867 18621
rect 20809 18581 20821 18615
rect 20855 18612 20867 18615
rect 20898 18612 20904 18624
rect 20855 18584 20904 18612
rect 20855 18581 20867 18584
rect 20809 18575 20867 18581
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 20990 18572 20996 18624
rect 21048 18572 21054 18624
rect 21818 18572 21824 18624
rect 21876 18572 21882 18624
rect 24489 18615 24547 18621
rect 24489 18581 24501 18615
rect 24535 18612 24547 18615
rect 24670 18612 24676 18624
rect 24535 18584 24676 18612
rect 24535 18581 24547 18584
rect 24489 18575 24547 18581
rect 24670 18572 24676 18584
rect 24728 18572 24734 18624
rect 24946 18572 24952 18624
rect 25004 18612 25010 18624
rect 26145 18615 26203 18621
rect 26145 18612 26157 18615
rect 25004 18584 26157 18612
rect 25004 18572 25010 18584
rect 26145 18581 26157 18584
rect 26191 18581 26203 18615
rect 26145 18575 26203 18581
rect 26605 18615 26663 18621
rect 26605 18581 26617 18615
rect 26651 18612 26663 18615
rect 27062 18612 27068 18624
rect 26651 18584 27068 18612
rect 26651 18581 26663 18584
rect 26605 18575 26663 18581
rect 27062 18572 27068 18584
rect 27120 18572 27126 18624
rect 27154 18572 27160 18624
rect 27212 18612 27218 18624
rect 27341 18615 27399 18621
rect 27341 18612 27353 18615
rect 27212 18584 27353 18612
rect 27212 18572 27218 18584
rect 27341 18581 27353 18584
rect 27387 18581 27399 18615
rect 27341 18575 27399 18581
rect 27801 18615 27859 18621
rect 27801 18581 27813 18615
rect 27847 18612 27859 18615
rect 28166 18612 28172 18624
rect 27847 18584 28172 18612
rect 27847 18581 27859 18584
rect 27801 18575 27859 18581
rect 28166 18572 28172 18584
rect 28224 18572 28230 18624
rect 1104 18522 29600 18544
rect 1104 18470 8034 18522
rect 8086 18470 8098 18522
rect 8150 18470 8162 18522
rect 8214 18470 8226 18522
rect 8278 18470 8290 18522
rect 8342 18470 15118 18522
rect 15170 18470 15182 18522
rect 15234 18470 15246 18522
rect 15298 18470 15310 18522
rect 15362 18470 15374 18522
rect 15426 18470 22202 18522
rect 22254 18470 22266 18522
rect 22318 18470 22330 18522
rect 22382 18470 22394 18522
rect 22446 18470 22458 18522
rect 22510 18470 29286 18522
rect 29338 18470 29350 18522
rect 29402 18470 29414 18522
rect 29466 18470 29478 18522
rect 29530 18470 29542 18522
rect 29594 18470 29600 18522
rect 1104 18448 29600 18470
rect 2498 18368 2504 18420
rect 2556 18408 2562 18420
rect 6914 18408 6920 18420
rect 2556 18380 6920 18408
rect 2556 18368 2562 18380
rect 2225 18343 2283 18349
rect 2225 18309 2237 18343
rect 2271 18340 2283 18343
rect 2590 18340 2596 18352
rect 2271 18312 2596 18340
rect 2271 18309 2283 18312
rect 2225 18303 2283 18309
rect 2590 18300 2596 18312
rect 2648 18300 2654 18352
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 4080 18281 4108 18380
rect 6914 18368 6920 18380
rect 6972 18368 6978 18420
rect 8386 18368 8392 18420
rect 8444 18408 8450 18420
rect 9125 18411 9183 18417
rect 9125 18408 9137 18411
rect 8444 18380 9137 18408
rect 8444 18368 8450 18380
rect 9125 18377 9137 18380
rect 9171 18408 9183 18411
rect 9490 18408 9496 18420
rect 9171 18380 9496 18408
rect 9171 18377 9183 18380
rect 9125 18371 9183 18377
rect 9490 18368 9496 18380
rect 9548 18368 9554 18420
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 9953 18411 10011 18417
rect 9953 18408 9965 18411
rect 9732 18380 9965 18408
rect 9732 18368 9738 18380
rect 9953 18377 9965 18380
rect 9999 18408 10011 18411
rect 10410 18408 10416 18420
rect 9999 18380 10416 18408
rect 9999 18377 10011 18380
rect 9953 18371 10011 18377
rect 10410 18368 10416 18380
rect 10468 18368 10474 18420
rect 14461 18411 14519 18417
rect 14461 18408 14473 18411
rect 13188 18380 14473 18408
rect 4982 18340 4988 18352
rect 4895 18312 4988 18340
rect 4982 18300 4988 18312
rect 5040 18340 5046 18352
rect 5166 18340 5172 18352
rect 5040 18312 5172 18340
rect 5040 18300 5046 18312
rect 5166 18300 5172 18312
rect 5224 18300 5230 18352
rect 7282 18340 7288 18352
rect 6748 18312 7288 18340
rect 6748 18281 6776 18312
rect 7282 18300 7288 18312
rect 7340 18300 7346 18352
rect 11974 18340 11980 18352
rect 11808 18312 11980 18340
rect 1857 18275 1915 18281
rect 1857 18272 1869 18275
rect 1636 18244 1869 18272
rect 1636 18232 1642 18244
rect 1857 18241 1869 18244
rect 1903 18241 1915 18275
rect 1857 18235 1915 18241
rect 4065 18275 4123 18281
rect 4065 18241 4077 18275
rect 4111 18241 4123 18275
rect 4065 18235 4123 18241
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18241 6791 18275
rect 6733 18235 6791 18241
rect 6917 18275 6975 18281
rect 6917 18241 6929 18275
rect 6963 18272 6975 18275
rect 7466 18272 7472 18284
rect 6963 18244 7472 18272
rect 6963 18241 6975 18244
rect 6917 18235 6975 18241
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 7650 18272 7656 18284
rect 7611 18244 7656 18272
rect 7650 18232 7656 18244
rect 7708 18232 7714 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7760 18244 7849 18272
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18204 4031 18207
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 4019 18176 6837 18204
rect 4019 18173 4031 18176
rect 3973 18167 4031 18173
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6825 18167 6883 18173
rect 4982 18096 4988 18148
rect 5040 18136 5046 18148
rect 7760 18136 7788 18244
rect 7837 18241 7849 18244
rect 7883 18272 7895 18275
rect 8297 18275 8355 18281
rect 8297 18272 8309 18275
rect 7883 18244 8309 18272
rect 7883 18241 7895 18244
rect 7837 18235 7895 18241
rect 8297 18241 8309 18244
rect 8343 18272 8355 18275
rect 8386 18272 8392 18284
rect 8343 18244 8392 18272
rect 8343 18241 8355 18244
rect 8297 18235 8355 18241
rect 8386 18232 8392 18244
rect 8444 18272 8450 18284
rect 8570 18272 8576 18284
rect 8444 18244 8576 18272
rect 8444 18232 8450 18244
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 11808 18281 11836 18312
rect 11974 18300 11980 18312
rect 12032 18300 12038 18352
rect 11793 18275 11851 18281
rect 11793 18241 11805 18275
rect 11839 18241 11851 18275
rect 12066 18272 12072 18284
rect 12027 18244 12072 18272
rect 11793 18235 11851 18241
rect 12066 18232 12072 18244
rect 12124 18232 12130 18284
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 12618 18204 12624 18216
rect 11931 18176 12624 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 5040 18108 7788 18136
rect 5040 18096 5046 18108
rect 9214 18096 9220 18148
rect 9272 18136 9278 18148
rect 11977 18139 12035 18145
rect 9272 18108 11744 18136
rect 9272 18096 9278 18108
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 4433 18071 4491 18077
rect 4433 18068 4445 18071
rect 4396 18040 4445 18068
rect 4396 18028 4402 18040
rect 4433 18037 4445 18040
rect 4479 18037 4491 18071
rect 5258 18068 5264 18080
rect 5219 18040 5264 18068
rect 4433 18031 4491 18037
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 7742 18068 7748 18080
rect 7703 18040 7748 18068
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 9950 18028 9956 18080
rect 10008 18068 10014 18080
rect 10413 18071 10471 18077
rect 10413 18068 10425 18071
rect 10008 18040 10425 18068
rect 10008 18028 10014 18040
rect 10413 18037 10425 18040
rect 10459 18068 10471 18071
rect 10870 18068 10876 18080
rect 10459 18040 10876 18068
rect 10459 18037 10471 18040
rect 10413 18031 10471 18037
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11609 18071 11667 18077
rect 11609 18068 11621 18071
rect 11112 18040 11621 18068
rect 11112 18028 11118 18040
rect 11609 18037 11621 18040
rect 11655 18037 11667 18071
rect 11716 18068 11744 18108
rect 11977 18105 11989 18139
rect 12023 18136 12035 18139
rect 13188 18136 13216 18380
rect 14461 18377 14473 18380
rect 14507 18377 14519 18411
rect 14461 18371 14519 18377
rect 15562 18368 15568 18420
rect 15620 18408 15626 18420
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 15620 18380 16681 18408
rect 15620 18368 15626 18380
rect 16669 18377 16681 18380
rect 16715 18377 16727 18411
rect 17770 18408 17776 18420
rect 17731 18380 17776 18408
rect 16669 18371 16727 18377
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 20533 18411 20591 18417
rect 20533 18408 20545 18411
rect 18380 18380 20545 18408
rect 18380 18368 18386 18380
rect 20533 18377 20545 18380
rect 20579 18377 20591 18411
rect 20533 18371 20591 18377
rect 27706 18368 27712 18420
rect 27764 18408 27770 18420
rect 28169 18411 28227 18417
rect 28169 18408 28181 18411
rect 27764 18380 28181 18408
rect 27764 18368 27770 18380
rect 28169 18377 28181 18380
rect 28215 18377 28227 18411
rect 28169 18371 28227 18377
rect 13262 18300 13268 18352
rect 13320 18340 13326 18352
rect 14737 18343 14795 18349
rect 14737 18340 14749 18343
rect 13320 18312 14749 18340
rect 13320 18300 13326 18312
rect 14737 18309 14749 18312
rect 14783 18309 14795 18343
rect 14737 18303 14795 18309
rect 14829 18343 14887 18349
rect 14829 18309 14841 18343
rect 14875 18340 14887 18343
rect 15470 18340 15476 18352
rect 14875 18312 15476 18340
rect 14875 18309 14887 18312
rect 14829 18303 14887 18309
rect 15470 18300 15476 18312
rect 15528 18300 15534 18352
rect 18138 18340 18144 18352
rect 17052 18312 18144 18340
rect 14642 18272 14648 18284
rect 14603 18244 14648 18272
rect 14642 18232 14648 18244
rect 14700 18232 14706 18284
rect 15010 18272 15016 18284
rect 14971 18244 15016 18272
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 16850 18272 16856 18284
rect 16811 18244 16856 18272
rect 16850 18232 16856 18244
rect 16908 18232 16914 18284
rect 17052 18281 17080 18312
rect 18138 18300 18144 18312
rect 18196 18340 18202 18352
rect 18233 18343 18291 18349
rect 18233 18340 18245 18343
rect 18196 18312 18245 18340
rect 18196 18300 18202 18312
rect 18233 18309 18245 18312
rect 18279 18340 18291 18343
rect 19978 18340 19984 18352
rect 18279 18312 19984 18340
rect 18279 18309 18291 18312
rect 18233 18303 18291 18309
rect 19978 18300 19984 18312
rect 20036 18300 20042 18352
rect 20806 18340 20812 18352
rect 20732 18312 20812 18340
rect 17037 18275 17095 18281
rect 17037 18241 17049 18275
rect 17083 18241 17095 18275
rect 17037 18235 17095 18241
rect 17129 18275 17187 18281
rect 17129 18241 17141 18275
rect 17175 18272 17187 18275
rect 20346 18272 20352 18284
rect 17175 18244 20352 18272
rect 17175 18241 17187 18244
rect 17129 18235 17187 18241
rect 20346 18232 20352 18244
rect 20404 18232 20410 18284
rect 20732 18281 20760 18312
rect 20806 18300 20812 18312
rect 20864 18300 20870 18352
rect 23106 18300 23112 18352
rect 23164 18340 23170 18352
rect 23477 18343 23535 18349
rect 23477 18340 23489 18343
rect 23164 18312 23489 18340
rect 23164 18300 23170 18312
rect 23477 18309 23489 18312
rect 23523 18309 23535 18343
rect 23477 18303 23535 18309
rect 23661 18343 23719 18349
rect 23661 18309 23673 18343
rect 23707 18340 23719 18343
rect 24946 18340 24952 18352
rect 23707 18312 24952 18340
rect 23707 18309 23719 18312
rect 23661 18303 23719 18309
rect 24946 18300 24952 18312
rect 25004 18300 25010 18352
rect 26510 18300 26516 18352
rect 26568 18340 26574 18352
rect 26568 18312 27292 18340
rect 26568 18300 26574 18312
rect 20717 18275 20775 18281
rect 20717 18241 20729 18275
rect 20763 18241 20775 18275
rect 20717 18235 20775 18241
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 21177 18275 21235 18281
rect 21177 18272 21189 18275
rect 20956 18244 21189 18272
rect 20956 18232 20962 18244
rect 21177 18241 21189 18244
rect 21223 18272 21235 18275
rect 21450 18272 21456 18284
rect 21223 18244 21456 18272
rect 21223 18241 21235 18244
rect 21177 18235 21235 18241
rect 21450 18232 21456 18244
rect 21508 18232 21514 18284
rect 27154 18272 27160 18284
rect 27115 18244 27160 18272
rect 27154 18232 27160 18244
rect 27212 18232 27218 18284
rect 27264 18281 27292 18312
rect 27249 18275 27307 18281
rect 27249 18241 27261 18275
rect 27295 18272 27307 18275
rect 27522 18272 27528 18284
rect 27295 18244 27528 18272
rect 27295 18241 27307 18244
rect 27249 18235 27307 18241
rect 27522 18232 27528 18244
rect 27580 18232 27586 18284
rect 14366 18204 14372 18216
rect 12023 18108 13216 18136
rect 13832 18176 14372 18204
rect 12023 18105 12035 18108
rect 11977 18099 12035 18105
rect 13832 18068 13860 18176
rect 14366 18164 14372 18176
rect 14424 18204 14430 18216
rect 14424 18176 14596 18204
rect 14424 18164 14430 18176
rect 14568 18136 14596 18176
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 16942 18204 16948 18216
rect 16632 18176 16948 18204
rect 16632 18164 16638 18176
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 20806 18204 20812 18216
rect 20767 18176 20812 18204
rect 20806 18164 20812 18176
rect 20864 18164 20870 18216
rect 23750 18204 23756 18216
rect 23711 18176 23756 18204
rect 23750 18164 23756 18176
rect 23808 18164 23814 18216
rect 26694 18164 26700 18216
rect 26752 18204 26758 18216
rect 26973 18207 27031 18213
rect 26973 18204 26985 18207
rect 26752 18176 26985 18204
rect 26752 18164 26758 18176
rect 26973 18173 26985 18176
rect 27019 18173 27031 18207
rect 26973 18167 27031 18173
rect 23201 18139 23259 18145
rect 23201 18136 23213 18139
rect 14568 18108 23213 18136
rect 23201 18105 23213 18108
rect 23247 18105 23259 18139
rect 23201 18099 23259 18105
rect 11716 18040 13860 18068
rect 11609 18031 11667 18037
rect 13998 18028 14004 18080
rect 14056 18068 14062 18080
rect 14274 18068 14280 18080
rect 14056 18040 14280 18068
rect 14056 18028 14062 18040
rect 14274 18028 14280 18040
rect 14332 18028 14338 18080
rect 16117 18071 16175 18077
rect 16117 18037 16129 18071
rect 16163 18068 16175 18071
rect 16758 18068 16764 18080
rect 16163 18040 16764 18068
rect 16163 18037 16175 18040
rect 16117 18031 16175 18037
rect 16758 18028 16764 18040
rect 16816 18068 16822 18080
rect 17310 18068 17316 18080
rect 16816 18040 17316 18068
rect 16816 18028 16822 18040
rect 17310 18028 17316 18040
rect 17368 18028 17374 18080
rect 19886 18028 19892 18080
rect 19944 18068 19950 18080
rect 19981 18071 20039 18077
rect 19981 18068 19993 18071
rect 19944 18040 19993 18068
rect 19944 18028 19950 18040
rect 19981 18037 19993 18040
rect 20027 18037 20039 18071
rect 21082 18068 21088 18080
rect 21043 18040 21088 18068
rect 19981 18031 20039 18037
rect 21082 18028 21088 18040
rect 21140 18028 21146 18080
rect 27062 18068 27068 18080
rect 27023 18040 27068 18068
rect 27062 18028 27068 18040
rect 27120 18028 27126 18080
rect 1104 17978 29440 18000
rect 1104 17926 4492 17978
rect 4544 17926 4556 17978
rect 4608 17926 4620 17978
rect 4672 17926 4684 17978
rect 4736 17926 4748 17978
rect 4800 17926 11576 17978
rect 11628 17926 11640 17978
rect 11692 17926 11704 17978
rect 11756 17926 11768 17978
rect 11820 17926 11832 17978
rect 11884 17926 18660 17978
rect 18712 17926 18724 17978
rect 18776 17926 18788 17978
rect 18840 17926 18852 17978
rect 18904 17926 18916 17978
rect 18968 17926 25744 17978
rect 25796 17926 25808 17978
rect 25860 17926 25872 17978
rect 25924 17926 25936 17978
rect 25988 17926 26000 17978
rect 26052 17926 29440 17978
rect 1104 17904 29440 17926
rect 4356 17836 6960 17864
rect 1578 17796 1584 17808
rect 1539 17768 1584 17796
rect 1578 17756 1584 17768
rect 1636 17756 1642 17808
rect 4154 17796 4160 17808
rect 4115 17768 4160 17796
rect 4154 17756 4160 17768
rect 4212 17756 4218 17808
rect 4356 17669 4384 17836
rect 5258 17756 5264 17808
rect 5316 17796 5322 17808
rect 6546 17796 6552 17808
rect 5316 17768 6552 17796
rect 5316 17756 5322 17768
rect 6546 17756 6552 17768
rect 6604 17756 6610 17808
rect 6932 17796 6960 17836
rect 7006 17824 7012 17876
rect 7064 17864 7070 17876
rect 10965 17867 11023 17873
rect 10965 17864 10977 17867
rect 7064 17836 10977 17864
rect 7064 17824 7070 17836
rect 10965 17833 10977 17836
rect 11011 17833 11023 17867
rect 10965 17827 11023 17833
rect 11882 17824 11888 17876
rect 11940 17864 11946 17876
rect 11974 17864 11980 17876
rect 11940 17836 11980 17864
rect 11940 17824 11946 17836
rect 11974 17824 11980 17836
rect 12032 17864 12038 17876
rect 13814 17864 13820 17876
rect 12032 17836 13820 17864
rect 12032 17824 12038 17836
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 17770 17824 17776 17876
rect 17828 17864 17834 17876
rect 17865 17867 17923 17873
rect 17865 17864 17877 17867
rect 17828 17836 17877 17864
rect 17828 17824 17834 17836
rect 17865 17833 17877 17836
rect 17911 17833 17923 17867
rect 17865 17827 17923 17833
rect 18046 17824 18052 17876
rect 18104 17864 18110 17876
rect 18601 17867 18659 17873
rect 18601 17864 18613 17867
rect 18104 17836 18613 17864
rect 18104 17824 18110 17836
rect 18601 17833 18613 17836
rect 18647 17833 18659 17867
rect 18601 17827 18659 17833
rect 10594 17796 10600 17808
rect 6932 17768 10600 17796
rect 10594 17756 10600 17768
rect 10652 17756 10658 17808
rect 13173 17799 13231 17805
rect 13173 17765 13185 17799
rect 13219 17796 13231 17799
rect 13538 17796 13544 17808
rect 13219 17768 13544 17796
rect 13219 17765 13231 17768
rect 13173 17759 13231 17765
rect 13538 17756 13544 17768
rect 13596 17756 13602 17808
rect 16669 17799 16727 17805
rect 16669 17765 16681 17799
rect 16715 17765 16727 17799
rect 16669 17759 16727 17765
rect 6457 17731 6515 17737
rect 6457 17697 6469 17731
rect 6503 17728 6515 17731
rect 7101 17731 7159 17737
rect 7101 17728 7113 17731
rect 6503 17700 7113 17728
rect 6503 17697 6515 17700
rect 6457 17691 6515 17697
rect 7101 17697 7113 17700
rect 7147 17697 7159 17731
rect 7282 17728 7288 17740
rect 7243 17700 7288 17728
rect 7101 17691 7159 17697
rect 7282 17688 7288 17700
rect 7340 17688 7346 17740
rect 7377 17731 7435 17737
rect 7377 17697 7389 17731
rect 7423 17728 7435 17731
rect 7742 17728 7748 17740
rect 7423 17700 7748 17728
rect 7423 17697 7435 17700
rect 7377 17691 7435 17697
rect 7742 17688 7748 17700
rect 7800 17728 7806 17740
rect 11054 17728 11060 17740
rect 7800 17700 9628 17728
rect 11015 17700 11060 17728
rect 7800 17688 7806 17700
rect 4341 17663 4399 17669
rect 4341 17629 4353 17663
rect 4387 17629 4399 17663
rect 4341 17623 4399 17629
rect 4430 17620 4436 17672
rect 4488 17660 4494 17672
rect 4617 17663 4675 17669
rect 4617 17660 4629 17663
rect 4488 17632 4629 17660
rect 4488 17620 4494 17632
rect 4617 17629 4629 17632
rect 4663 17629 4675 17663
rect 5718 17660 5724 17672
rect 5679 17632 5724 17660
rect 4617 17623 4675 17629
rect 5718 17620 5724 17632
rect 5776 17620 5782 17672
rect 6362 17660 6368 17672
rect 6323 17632 6368 17660
rect 6362 17620 6368 17632
rect 6420 17620 6426 17672
rect 6546 17660 6552 17672
rect 6507 17632 6552 17660
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 7193 17663 7251 17669
rect 7193 17629 7205 17663
rect 7239 17660 7251 17663
rect 7466 17660 7472 17672
rect 7239 17632 7472 17660
rect 7239 17629 7251 17632
rect 7193 17623 7251 17629
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 7650 17620 7656 17672
rect 7708 17660 7714 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7708 17632 8217 17660
rect 7708 17620 7714 17632
rect 8205 17629 8217 17632
rect 8251 17660 8263 17663
rect 9030 17660 9036 17672
rect 8251 17632 9036 17660
rect 8251 17629 8263 17632
rect 8205 17623 8263 17629
rect 9030 17620 9036 17632
rect 9088 17620 9094 17672
rect 9488 17663 9546 17669
rect 9488 17660 9500 17663
rect 9416 17632 9500 17660
rect 2222 17552 2228 17604
rect 2280 17592 2286 17604
rect 4249 17595 4307 17601
rect 4249 17592 4261 17595
rect 2280 17564 4261 17592
rect 2280 17552 2286 17564
rect 4249 17561 4261 17564
rect 4295 17561 4307 17595
rect 4249 17555 4307 17561
rect 4985 17595 5043 17601
rect 4985 17561 4997 17595
rect 5031 17592 5043 17595
rect 5166 17592 5172 17604
rect 5031 17564 5172 17592
rect 5031 17561 5043 17564
rect 4985 17555 5043 17561
rect 5166 17552 5172 17564
rect 5224 17592 5230 17604
rect 7098 17592 7104 17604
rect 5224 17564 7104 17592
rect 5224 17552 5230 17564
rect 7098 17552 7104 17564
rect 7156 17552 7162 17604
rect 8386 17592 8392 17604
rect 8347 17564 8392 17592
rect 8386 17552 8392 17564
rect 8444 17552 8450 17604
rect 2866 17484 2872 17536
rect 2924 17524 2930 17536
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 2924 17496 5825 17524
rect 2924 17484 2930 17496
rect 5813 17493 5825 17496
rect 5859 17493 5871 17527
rect 7558 17524 7564 17536
rect 7519 17496 7564 17524
rect 5813 17487 5871 17493
rect 7558 17484 7564 17496
rect 7616 17484 7622 17536
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7984 17496 8033 17524
rect 7984 17484 7990 17496
rect 8021 17493 8033 17496
rect 8067 17493 8079 17527
rect 9306 17524 9312 17536
rect 9267 17496 9312 17524
rect 8021 17487 8079 17493
rect 9306 17484 9312 17496
rect 9364 17484 9370 17536
rect 9416 17524 9444 17632
rect 9488 17629 9500 17632
rect 9534 17629 9546 17663
rect 9600 17660 9628 17700
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 16574 17728 16580 17740
rect 16040 17700 16580 17728
rect 9805 17663 9863 17669
rect 9805 17660 9817 17663
rect 9600 17632 9817 17660
rect 9488 17623 9546 17629
rect 9805 17629 9817 17632
rect 9851 17629 9863 17663
rect 9805 17623 9863 17629
rect 9950 17620 9956 17672
rect 10008 17660 10014 17672
rect 10781 17663 10839 17669
rect 10008 17632 10053 17660
rect 10008 17620 10014 17632
rect 10781 17629 10793 17663
rect 10827 17629 10839 17663
rect 10781 17623 10839 17629
rect 9582 17592 9588 17604
rect 9543 17564 9588 17592
rect 9582 17552 9588 17564
rect 9640 17552 9646 17604
rect 9674 17552 9680 17604
rect 9732 17592 9738 17604
rect 10796 17592 10824 17623
rect 10870 17620 10876 17672
rect 10928 17660 10934 17672
rect 10928 17632 10973 17660
rect 10928 17620 10934 17632
rect 12802 17620 12808 17672
rect 12860 17660 12866 17672
rect 13081 17663 13139 17669
rect 13081 17660 13093 17663
rect 12860 17632 13093 17660
rect 12860 17620 12866 17632
rect 13081 17629 13093 17632
rect 13127 17629 13139 17663
rect 13262 17660 13268 17672
rect 13223 17632 13268 17660
rect 13081 17623 13139 17629
rect 13262 17620 13268 17632
rect 13320 17620 13326 17672
rect 13357 17663 13415 17669
rect 13357 17629 13369 17663
rect 13403 17660 13415 17663
rect 14090 17660 14096 17672
rect 13403 17632 14096 17660
rect 13403 17629 13415 17632
rect 13357 17623 13415 17629
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14274 17660 14280 17672
rect 14235 17632 14280 17660
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 16040 17669 16068 17700
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17629 16083 17663
rect 16025 17623 16083 17629
rect 16209 17663 16267 17669
rect 16209 17629 16221 17663
rect 16255 17660 16267 17663
rect 16684 17660 16712 17759
rect 17126 17728 17132 17740
rect 17087 17700 17132 17728
rect 17126 17688 17132 17700
rect 17184 17688 17190 17740
rect 17313 17731 17371 17737
rect 17313 17697 17325 17731
rect 17359 17728 17371 17731
rect 17788 17728 17816 17824
rect 17359 17700 17816 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 16255 17632 16712 17660
rect 16255 17629 16267 17632
rect 16209 17623 16267 17629
rect 14458 17592 14464 17604
rect 9732 17564 9777 17592
rect 10796 17564 11652 17592
rect 14419 17564 14464 17592
rect 9732 17552 9738 17564
rect 9766 17524 9772 17536
rect 9416 17496 9772 17524
rect 9766 17484 9772 17496
rect 9824 17524 9830 17536
rect 10686 17524 10692 17536
rect 9824 17496 10692 17524
rect 9824 17484 9830 17496
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 11624 17533 11652 17564
rect 14458 17552 14464 17564
rect 14516 17552 14522 17604
rect 15565 17595 15623 17601
rect 15565 17561 15577 17595
rect 15611 17592 15623 17595
rect 16298 17592 16304 17604
rect 15611 17564 16304 17592
rect 15611 17561 15623 17564
rect 15565 17555 15623 17561
rect 16298 17552 16304 17564
rect 16356 17592 16362 17604
rect 17037 17595 17095 17601
rect 17037 17592 17049 17595
rect 16356 17564 17049 17592
rect 16356 17552 16362 17564
rect 17037 17561 17049 17564
rect 17083 17561 17095 17595
rect 18616 17592 18644 17827
rect 18690 17824 18696 17876
rect 18748 17864 18754 17876
rect 23382 17864 23388 17876
rect 18748 17836 23388 17864
rect 18748 17824 18754 17836
rect 23382 17824 23388 17836
rect 23440 17824 23446 17876
rect 26973 17867 27031 17873
rect 26973 17833 26985 17867
rect 27019 17864 27031 17867
rect 27798 17864 27804 17876
rect 27019 17836 27804 17864
rect 27019 17833 27031 17836
rect 26973 17827 27031 17833
rect 27798 17824 27804 17836
rect 27856 17824 27862 17876
rect 28718 17864 28724 17876
rect 28679 17836 28724 17864
rect 28718 17824 28724 17836
rect 28776 17824 28782 17876
rect 19242 17756 19248 17808
rect 19300 17796 19306 17808
rect 20533 17799 20591 17805
rect 20533 17796 20545 17799
rect 19300 17768 20545 17796
rect 19300 17756 19306 17768
rect 20533 17765 20545 17768
rect 20579 17765 20591 17799
rect 22373 17799 22431 17805
rect 22373 17796 22385 17799
rect 20533 17759 20591 17765
rect 22066 17768 22385 17796
rect 19334 17660 19340 17672
rect 19295 17632 19340 17660
rect 19334 17620 19340 17632
rect 19392 17620 19398 17672
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 21637 17663 21695 17669
rect 21637 17629 21649 17663
rect 21683 17660 21695 17663
rect 21726 17660 21732 17672
rect 21683 17632 21732 17660
rect 21683 17629 21695 17632
rect 21637 17623 21695 17629
rect 19720 17592 19748 17623
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17660 21879 17663
rect 21867 17632 21901 17660
rect 21867 17629 21879 17632
rect 21821 17623 21879 17629
rect 18616 17564 19748 17592
rect 17037 17555 17095 17561
rect 21542 17552 21548 17604
rect 21600 17592 21606 17604
rect 21836 17592 21864 17623
rect 22066 17592 22094 17768
rect 22373 17765 22385 17768
rect 22419 17796 22431 17799
rect 28350 17796 28356 17808
rect 22419 17768 28356 17796
rect 22419 17765 22431 17768
rect 22373 17759 22431 17765
rect 28350 17756 28356 17768
rect 28408 17756 28414 17808
rect 25409 17731 25467 17737
rect 25409 17728 25421 17731
rect 24780 17700 25421 17728
rect 24578 17620 24584 17672
rect 24636 17660 24642 17672
rect 24780 17669 24808 17700
rect 25409 17697 25421 17700
rect 25455 17697 25467 17731
rect 25409 17691 25467 17697
rect 27617 17731 27675 17737
rect 27617 17697 27629 17731
rect 27663 17728 27675 17731
rect 27890 17728 27896 17740
rect 27663 17700 27896 17728
rect 27663 17697 27675 17700
rect 27617 17691 27675 17697
rect 27890 17688 27896 17700
rect 27948 17688 27954 17740
rect 24765 17663 24823 17669
rect 24765 17660 24777 17663
rect 24636 17632 24777 17660
rect 24636 17620 24642 17632
rect 24765 17629 24777 17632
rect 24811 17629 24823 17663
rect 24946 17660 24952 17672
rect 24907 17632 24952 17660
rect 24765 17623 24823 17629
rect 24946 17620 24952 17632
rect 25004 17620 25010 17672
rect 27709 17663 27767 17669
rect 27709 17629 27721 17663
rect 27755 17660 27767 17663
rect 27798 17660 27804 17672
rect 27755 17632 27804 17660
rect 27755 17629 27767 17632
rect 27709 17623 27767 17629
rect 27798 17620 27804 17632
rect 27856 17620 27862 17672
rect 21600 17564 22094 17592
rect 21600 17552 21606 17564
rect 11609 17527 11667 17533
rect 11609 17493 11621 17527
rect 11655 17524 11667 17527
rect 12158 17524 12164 17536
rect 11655 17496 12164 17524
rect 11655 17493 11667 17496
rect 11609 17487 11667 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12894 17524 12900 17536
rect 12855 17496 12900 17524
rect 12894 17484 12900 17496
rect 12952 17484 12958 17536
rect 14090 17524 14096 17536
rect 14051 17496 14096 17524
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 15838 17484 15844 17536
rect 15896 17524 15902 17536
rect 16117 17527 16175 17533
rect 16117 17524 16129 17527
rect 15896 17496 16129 17524
rect 15896 17484 15902 17496
rect 16117 17493 16129 17496
rect 16163 17524 16175 17527
rect 16574 17524 16580 17536
rect 16163 17496 16580 17524
rect 16163 17493 16175 17496
rect 16117 17487 16175 17493
rect 16574 17484 16580 17496
rect 16632 17484 16638 17536
rect 21726 17524 21732 17536
rect 21687 17496 21732 17524
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 24486 17484 24492 17536
rect 24544 17524 24550 17536
rect 24765 17527 24823 17533
rect 24765 17524 24777 17527
rect 24544 17496 24777 17524
rect 24544 17484 24550 17496
rect 24765 17493 24777 17496
rect 24811 17493 24823 17527
rect 26326 17524 26332 17536
rect 26287 17496 26332 17524
rect 24765 17487 24823 17493
rect 26326 17484 26332 17496
rect 26384 17524 26390 17536
rect 26970 17524 26976 17536
rect 26384 17496 26976 17524
rect 26384 17484 26390 17496
rect 26970 17484 26976 17496
rect 27028 17524 27034 17536
rect 27801 17527 27859 17533
rect 27801 17524 27813 17527
rect 27028 17496 27813 17524
rect 27028 17484 27034 17496
rect 27801 17493 27813 17496
rect 27847 17493 27859 17527
rect 27801 17487 27859 17493
rect 28169 17527 28227 17533
rect 28169 17493 28181 17527
rect 28215 17524 28227 17527
rect 28350 17524 28356 17536
rect 28215 17496 28356 17524
rect 28215 17493 28227 17496
rect 28169 17487 28227 17493
rect 28350 17484 28356 17496
rect 28408 17484 28414 17536
rect 1104 17434 29600 17456
rect 1104 17382 8034 17434
rect 8086 17382 8098 17434
rect 8150 17382 8162 17434
rect 8214 17382 8226 17434
rect 8278 17382 8290 17434
rect 8342 17382 15118 17434
rect 15170 17382 15182 17434
rect 15234 17382 15246 17434
rect 15298 17382 15310 17434
rect 15362 17382 15374 17434
rect 15426 17382 22202 17434
rect 22254 17382 22266 17434
rect 22318 17382 22330 17434
rect 22382 17382 22394 17434
rect 22446 17382 22458 17434
rect 22510 17382 29286 17434
rect 29338 17382 29350 17434
rect 29402 17382 29414 17434
rect 29466 17382 29478 17434
rect 29530 17382 29542 17434
rect 29594 17382 29600 17434
rect 1104 17360 29600 17382
rect 4801 17323 4859 17329
rect 4801 17289 4813 17323
rect 4847 17320 4859 17323
rect 4982 17320 4988 17332
rect 4847 17292 4988 17320
rect 4847 17289 4859 17292
rect 4801 17283 4859 17289
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 7561 17323 7619 17329
rect 7561 17320 7573 17323
rect 6972 17292 7573 17320
rect 6972 17280 6978 17292
rect 7561 17289 7573 17292
rect 7607 17289 7619 17323
rect 12894 17320 12900 17332
rect 7561 17283 7619 17289
rect 11992 17292 12900 17320
rect 9306 17212 9312 17264
rect 9364 17252 9370 17264
rect 9858 17252 9864 17264
rect 9364 17224 9628 17252
rect 9819 17224 9864 17252
rect 9364 17212 9370 17224
rect 1762 17144 1768 17196
rect 1820 17184 1826 17196
rect 2133 17187 2191 17193
rect 2133 17184 2145 17187
rect 1820 17156 2145 17184
rect 1820 17144 1826 17156
rect 2133 17153 2145 17156
rect 2179 17153 2191 17187
rect 2133 17147 2191 17153
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17184 7619 17187
rect 7650 17184 7656 17196
rect 7607 17156 7656 17184
rect 7607 17153 7619 17156
rect 7561 17147 7619 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17153 7803 17187
rect 9490 17184 9496 17196
rect 9451 17156 9496 17184
rect 7745 17147 7803 17153
rect 2225 17119 2283 17125
rect 2225 17085 2237 17119
rect 2271 17116 2283 17119
rect 5810 17116 5816 17128
rect 2271 17088 5816 17116
rect 2271 17085 2283 17088
rect 2225 17079 2283 17085
rect 5810 17076 5816 17088
rect 5868 17076 5874 17128
rect 7760 17116 7788 17147
rect 9490 17144 9496 17156
rect 9548 17144 9554 17196
rect 9600 17193 9628 17224
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 10042 17212 10048 17264
rect 10100 17212 10106 17264
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 9769 17187 9827 17193
rect 9769 17153 9781 17187
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17184 10011 17187
rect 10060 17184 10088 17212
rect 11882 17184 11888 17196
rect 9999 17156 10088 17184
rect 11843 17156 11888 17184
rect 9999 17153 10011 17156
rect 9953 17147 10011 17153
rect 7926 17116 7932 17128
rect 7760 17088 7932 17116
rect 7926 17076 7932 17088
rect 7984 17116 7990 17128
rect 9784 17116 9812 17147
rect 11882 17144 11888 17156
rect 11940 17144 11946 17196
rect 11992 17193 12020 17292
rect 12894 17280 12900 17292
rect 12952 17280 12958 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17289 13231 17323
rect 13173 17283 13231 17289
rect 13188 17252 13216 17283
rect 14642 17280 14648 17332
rect 14700 17320 14706 17332
rect 15194 17320 15200 17332
rect 14700 17292 15200 17320
rect 14700 17280 14706 17292
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 16761 17323 16819 17329
rect 16761 17289 16773 17323
rect 16807 17320 16819 17323
rect 17126 17320 17132 17332
rect 16807 17292 17132 17320
rect 16807 17289 16819 17292
rect 16761 17283 16819 17289
rect 17126 17280 17132 17292
rect 17184 17280 17190 17332
rect 21266 17320 21272 17332
rect 21227 17292 21272 17320
rect 21266 17280 21272 17292
rect 21324 17320 21330 17332
rect 22002 17320 22008 17332
rect 21324 17292 22008 17320
rect 21324 17280 21330 17292
rect 22002 17280 22008 17292
rect 22060 17280 22066 17332
rect 23382 17320 23388 17332
rect 23343 17292 23388 17320
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 27890 17280 27896 17332
rect 27948 17320 27954 17332
rect 28261 17323 28319 17329
rect 28261 17320 28273 17323
rect 27948 17292 28273 17320
rect 27948 17280 27954 17292
rect 28261 17289 28273 17292
rect 28307 17289 28319 17323
rect 28261 17283 28319 17289
rect 12084 17224 13216 17252
rect 20349 17255 20407 17261
rect 12084 17193 12112 17224
rect 20349 17221 20361 17255
rect 20395 17252 20407 17255
rect 23750 17252 23756 17264
rect 20395 17224 23756 17252
rect 20395 17221 20407 17224
rect 20349 17215 20407 17221
rect 23750 17212 23756 17224
rect 23808 17252 23814 17264
rect 24121 17255 24179 17261
rect 24121 17252 24133 17255
rect 23808 17224 24133 17252
rect 23808 17212 23814 17224
rect 24121 17221 24133 17224
rect 24167 17221 24179 17255
rect 24121 17215 24179 17221
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 12069 17187 12127 17193
rect 12069 17153 12081 17187
rect 12115 17153 12127 17187
rect 12069 17147 12127 17153
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17153 12311 17187
rect 12253 17147 12311 17153
rect 7984 17088 9812 17116
rect 10045 17119 10103 17125
rect 7984 17076 7990 17088
rect 10045 17085 10057 17119
rect 10091 17116 10103 17119
rect 12268 17116 12296 17147
rect 12986 17144 12992 17196
rect 13044 17184 13050 17196
rect 13357 17187 13415 17193
rect 13357 17184 13369 17187
rect 13044 17156 13369 17184
rect 13044 17144 13050 17156
rect 13357 17153 13369 17156
rect 13403 17184 13415 17187
rect 13633 17187 13691 17193
rect 13403 17156 13584 17184
rect 13403 17153 13415 17156
rect 13357 17147 13415 17153
rect 10091 17088 12296 17116
rect 13449 17119 13507 17125
rect 10091 17085 10103 17088
rect 10045 17079 10103 17085
rect 13449 17085 13461 17119
rect 13495 17085 13507 17119
rect 13556 17116 13584 17156
rect 13633 17153 13645 17187
rect 13679 17184 13691 17187
rect 13906 17184 13912 17196
rect 13679 17156 13912 17184
rect 13679 17153 13691 17156
rect 13633 17147 13691 17153
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 19334 17184 19340 17196
rect 19295 17156 19340 17184
rect 19334 17144 19340 17156
rect 19392 17144 19398 17196
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 15470 17116 15476 17128
rect 13556 17088 15476 17116
rect 13449 17079 13507 17085
rect 6457 17051 6515 17057
rect 6457 17017 6469 17051
rect 6503 17048 6515 17051
rect 6546 17048 6552 17060
rect 6503 17020 6552 17048
rect 6503 17017 6515 17020
rect 6457 17011 6515 17017
rect 6546 17008 6552 17020
rect 6604 17048 6610 17060
rect 8481 17051 8539 17057
rect 8481 17048 8493 17051
rect 6604 17020 8493 17048
rect 6604 17008 6610 17020
rect 8481 17017 8493 17020
rect 8527 17048 8539 17051
rect 8570 17048 8576 17060
rect 8527 17020 8576 17048
rect 8527 17017 8539 17020
rect 8481 17011 8539 17017
rect 8570 17008 8576 17020
rect 8628 17008 8634 17060
rect 13464 17048 13492 17079
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 18414 17076 18420 17128
rect 18472 17116 18478 17128
rect 19536 17116 19564 17147
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 21726 17184 21732 17196
rect 20772 17156 21732 17184
rect 20772 17144 20778 17156
rect 21726 17144 21732 17156
rect 21784 17184 21790 17196
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 21784 17156 21833 17184
rect 21784 17144 21790 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 22002 17144 22008 17196
rect 22060 17184 22066 17196
rect 22097 17187 22155 17193
rect 22097 17184 22109 17187
rect 22060 17156 22109 17184
rect 22060 17144 22066 17156
rect 22097 17153 22109 17156
rect 22143 17153 22155 17187
rect 22097 17147 22155 17153
rect 22554 17144 22560 17196
rect 22612 17184 22618 17196
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 22612 17156 22845 17184
rect 22612 17144 22618 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 23109 17187 23167 17193
rect 23109 17153 23121 17187
rect 23155 17153 23167 17187
rect 23109 17147 23167 17153
rect 18472 17088 19564 17116
rect 18472 17076 18478 17088
rect 21174 17076 21180 17128
rect 21232 17116 21238 17128
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 21232 17088 21925 17116
rect 21232 17076 21238 17088
rect 21913 17085 21925 17088
rect 21959 17085 21971 17119
rect 23124 17116 23152 17147
rect 23198 17144 23204 17196
rect 23256 17184 23262 17196
rect 27246 17184 27252 17196
rect 23256 17156 23301 17184
rect 27207 17156 27252 17184
rect 23256 17144 23262 17156
rect 27246 17144 27252 17156
rect 27304 17144 27310 17196
rect 27341 17187 27399 17193
rect 27341 17153 27353 17187
rect 27387 17184 27399 17187
rect 27522 17184 27528 17196
rect 27387 17156 27528 17184
rect 27387 17153 27399 17156
rect 27341 17147 27399 17153
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 23566 17116 23572 17128
rect 23124 17088 23572 17116
rect 21913 17079 21971 17085
rect 23566 17076 23572 17088
rect 23624 17076 23630 17128
rect 26326 17116 26332 17128
rect 24136 17088 26332 17116
rect 13814 17048 13820 17060
rect 13464 17020 13820 17048
rect 13814 17008 13820 17020
rect 13872 17048 13878 17060
rect 15562 17048 15568 17060
rect 13872 17020 15568 17048
rect 13872 17008 13878 17020
rect 15562 17008 15568 17020
rect 15620 17008 15626 17060
rect 17218 17008 17224 17060
rect 17276 17048 17282 17060
rect 24136 17048 24164 17088
rect 26326 17076 26332 17088
rect 26384 17076 26390 17128
rect 27065 17119 27123 17125
rect 27065 17085 27077 17119
rect 27111 17116 27123 17119
rect 27614 17116 27620 17128
rect 27111 17088 27620 17116
rect 27111 17085 27123 17088
rect 27065 17079 27123 17085
rect 27614 17076 27620 17088
rect 27672 17076 27678 17128
rect 24302 17048 24308 17060
rect 17276 17020 24164 17048
rect 24263 17020 24308 17048
rect 17276 17008 17282 17020
rect 24302 17008 24308 17020
rect 24360 17008 24366 17060
rect 1857 16983 1915 16989
rect 1857 16949 1869 16983
rect 1903 16980 1915 16983
rect 1946 16980 1952 16992
rect 1903 16952 1952 16980
rect 1903 16949 1915 16952
rect 1857 16943 1915 16949
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 5810 16980 5816 16992
rect 5723 16952 5816 16980
rect 5810 16940 5816 16952
rect 5868 16980 5874 16992
rect 6362 16980 6368 16992
rect 5868 16952 6368 16980
rect 5868 16940 5874 16952
rect 6362 16940 6368 16952
rect 6420 16980 6426 16992
rect 7101 16983 7159 16989
rect 7101 16980 7113 16983
rect 6420 16952 7113 16980
rect 6420 16940 6426 16952
rect 7101 16949 7113 16952
rect 7147 16980 7159 16983
rect 9030 16980 9036 16992
rect 7147 16952 9036 16980
rect 7147 16949 7159 16952
rect 7101 16943 7159 16949
rect 9030 16940 9036 16952
rect 9088 16980 9094 16992
rect 9582 16980 9588 16992
rect 9088 16952 9588 16980
rect 9088 16940 9094 16952
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 10597 16983 10655 16989
rect 10597 16949 10609 16983
rect 10643 16980 10655 16983
rect 10686 16980 10692 16992
rect 10643 16952 10692 16980
rect 10643 16949 10655 16952
rect 10597 16943 10655 16949
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 11422 16940 11428 16992
rect 11480 16980 11486 16992
rect 11609 16983 11667 16989
rect 11609 16980 11621 16983
rect 11480 16952 11621 16980
rect 11480 16940 11486 16952
rect 11609 16949 11621 16952
rect 11655 16949 11667 16983
rect 11609 16943 11667 16949
rect 13633 16983 13691 16989
rect 13633 16949 13645 16983
rect 13679 16980 13691 16983
rect 14090 16980 14096 16992
rect 13679 16952 14096 16980
rect 13679 16949 13691 16952
rect 13633 16943 13691 16949
rect 14090 16940 14096 16952
rect 14148 16980 14154 16992
rect 14274 16980 14280 16992
rect 14148 16952 14280 16980
rect 14148 16940 14154 16952
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 21634 16940 21640 16992
rect 21692 16980 21698 16992
rect 21821 16983 21879 16989
rect 21821 16980 21833 16983
rect 21692 16952 21833 16980
rect 21692 16940 21698 16952
rect 21821 16949 21833 16952
rect 21867 16949 21879 16983
rect 21821 16943 21879 16949
rect 22281 16983 22339 16989
rect 22281 16949 22293 16983
rect 22327 16980 22339 16983
rect 22646 16980 22652 16992
rect 22327 16952 22652 16980
rect 22327 16949 22339 16952
rect 22281 16943 22339 16949
rect 22646 16940 22652 16952
rect 22704 16940 22710 16992
rect 22922 16980 22928 16992
rect 22883 16952 22928 16980
rect 22922 16940 22928 16952
rect 22980 16940 22986 16992
rect 26786 16940 26792 16992
rect 26844 16980 26850 16992
rect 27157 16983 27215 16989
rect 27157 16980 27169 16983
rect 26844 16952 27169 16980
rect 26844 16940 26850 16952
rect 27157 16949 27169 16952
rect 27203 16949 27215 16983
rect 27157 16943 27215 16949
rect 1104 16890 29440 16912
rect 1104 16838 4492 16890
rect 4544 16838 4556 16890
rect 4608 16838 4620 16890
rect 4672 16838 4684 16890
rect 4736 16838 4748 16890
rect 4800 16838 11576 16890
rect 11628 16838 11640 16890
rect 11692 16838 11704 16890
rect 11756 16838 11768 16890
rect 11820 16838 11832 16890
rect 11884 16838 18660 16890
rect 18712 16838 18724 16890
rect 18776 16838 18788 16890
rect 18840 16838 18852 16890
rect 18904 16838 18916 16890
rect 18968 16838 25744 16890
rect 25796 16838 25808 16890
rect 25860 16838 25872 16890
rect 25924 16838 25936 16890
rect 25988 16838 26000 16890
rect 26052 16838 29440 16890
rect 1104 16816 29440 16838
rect 1762 16776 1768 16788
rect 1723 16748 1768 16776
rect 1762 16736 1768 16748
rect 1820 16736 1826 16788
rect 2866 16776 2872 16788
rect 2827 16748 2872 16776
rect 2866 16736 2872 16748
rect 2924 16736 2930 16788
rect 5166 16776 5172 16788
rect 5127 16748 5172 16776
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 7006 16736 7012 16788
rect 7064 16776 7070 16788
rect 7193 16779 7251 16785
rect 7193 16776 7205 16779
rect 7064 16748 7205 16776
rect 7064 16736 7070 16748
rect 7193 16745 7205 16748
rect 7239 16745 7251 16779
rect 7193 16739 7251 16745
rect 7929 16779 7987 16785
rect 7929 16745 7941 16779
rect 7975 16776 7987 16779
rect 8386 16776 8392 16788
rect 7975 16748 8392 16776
rect 7975 16745 7987 16748
rect 7929 16739 7987 16745
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 9490 16776 9496 16788
rect 9451 16748 9496 16776
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 9677 16779 9735 16785
rect 9677 16745 9689 16779
rect 9723 16776 9735 16779
rect 9858 16776 9864 16788
rect 9723 16748 9864 16776
rect 9723 16745 9735 16748
rect 9677 16739 9735 16745
rect 9858 16736 9864 16748
rect 9916 16736 9922 16788
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10321 16779 10379 16785
rect 10321 16776 10333 16779
rect 10100 16748 10333 16776
rect 10100 16736 10106 16748
rect 10321 16745 10333 16748
rect 10367 16745 10379 16779
rect 12618 16776 12624 16788
rect 12579 16748 12624 16776
rect 10321 16739 10379 16745
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 13906 16736 13912 16788
rect 13964 16776 13970 16788
rect 13964 16748 19288 16776
rect 13964 16736 13970 16748
rect 2222 16640 2228 16652
rect 2183 16612 2228 16640
rect 2222 16600 2228 16612
rect 2280 16600 2286 16652
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 9033 16643 9091 16649
rect 9033 16640 9045 16643
rect 8628 16612 9045 16640
rect 8628 16600 8634 16612
rect 9033 16609 9045 16612
rect 9079 16640 9091 16643
rect 9876 16640 9904 16736
rect 10594 16668 10600 16720
rect 10652 16708 10658 16720
rect 11517 16711 11575 16717
rect 11517 16708 11529 16711
rect 10652 16680 11529 16708
rect 10652 16668 10658 16680
rect 11517 16677 11529 16680
rect 11563 16677 11575 16711
rect 17218 16708 17224 16720
rect 11517 16671 11575 16677
rect 12406 16680 17224 16708
rect 12406 16640 12434 16680
rect 17218 16668 17224 16680
rect 17276 16668 17282 16720
rect 18138 16708 18144 16720
rect 18099 16680 18144 16708
rect 18138 16668 18144 16680
rect 18196 16708 18202 16720
rect 19150 16708 19156 16720
rect 18196 16680 19156 16708
rect 18196 16668 18202 16680
rect 19150 16668 19156 16680
rect 19208 16668 19214 16720
rect 19260 16708 19288 16748
rect 19334 16736 19340 16788
rect 19392 16776 19398 16788
rect 19797 16779 19855 16785
rect 19797 16776 19809 16779
rect 19392 16748 19809 16776
rect 19392 16736 19398 16748
rect 19797 16745 19809 16748
rect 19843 16745 19855 16779
rect 19797 16739 19855 16745
rect 20346 16736 20352 16788
rect 20404 16776 20410 16788
rect 21269 16779 21327 16785
rect 21269 16776 21281 16779
rect 20404 16748 21281 16776
rect 20404 16736 20410 16748
rect 21269 16745 21281 16748
rect 21315 16745 21327 16779
rect 26418 16776 26424 16788
rect 21269 16739 21327 16745
rect 23216 16748 26424 16776
rect 20714 16708 20720 16720
rect 19260 16680 20720 16708
rect 20714 16668 20720 16680
rect 20772 16708 20778 16720
rect 22922 16708 22928 16720
rect 20772 16680 21036 16708
rect 20772 16668 20778 16680
rect 9079 16612 12434 16640
rect 13081 16643 13139 16649
rect 9079 16609 9091 16612
rect 9033 16603 9091 16609
rect 13081 16609 13093 16643
rect 13127 16640 13139 16643
rect 13170 16640 13176 16652
rect 13127 16612 13176 16640
rect 13127 16609 13139 16612
rect 13081 16603 13139 16609
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 14829 16643 14887 16649
rect 14829 16640 14841 16643
rect 13596 16612 14841 16640
rect 13596 16600 13602 16612
rect 14829 16609 14841 16612
rect 14875 16609 14887 16643
rect 20898 16640 20904 16652
rect 14829 16603 14887 16609
rect 19996 16612 20904 16640
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16572 2191 16575
rect 2406 16572 2412 16584
rect 2179 16544 2412 16572
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 2406 16532 2412 16544
rect 2464 16572 2470 16584
rect 2866 16572 2872 16584
rect 2464 16544 2872 16572
rect 2464 16532 2470 16544
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 11422 16532 11428 16584
rect 11480 16572 11486 16584
rect 11701 16575 11759 16581
rect 11701 16572 11713 16575
rect 11480 16544 11713 16572
rect 11480 16532 11486 16544
rect 11701 16541 11713 16544
rect 11747 16541 11759 16575
rect 11882 16572 11888 16584
rect 11843 16544 11888 16572
rect 11701 16535 11759 16541
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 11977 16575 12035 16581
rect 11977 16541 11989 16575
rect 12023 16572 12035 16575
rect 12158 16572 12164 16584
rect 12023 16544 12164 16572
rect 12023 16541 12035 16544
rect 11977 16535 12035 16541
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 12618 16532 12624 16584
rect 12676 16572 12682 16584
rect 12802 16572 12808 16584
rect 12676 16544 12808 16572
rect 12676 16532 12682 16544
rect 12802 16532 12808 16544
rect 12860 16532 12866 16584
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16541 13047 16575
rect 12989 16535 13047 16541
rect 9858 16504 9864 16516
rect 9819 16476 9864 16504
rect 9858 16464 9864 16476
rect 9916 16464 9922 16516
rect 13004 16504 13032 16535
rect 13262 16532 13268 16584
rect 13320 16572 13326 16584
rect 18230 16572 18236 16584
rect 13320 16544 18236 16572
rect 13320 16532 13326 16544
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 19610 16532 19616 16584
rect 19668 16572 19674 16584
rect 19996 16581 20024 16612
rect 20898 16600 20904 16612
rect 20956 16600 20962 16652
rect 19705 16575 19763 16581
rect 19705 16572 19717 16575
rect 19668 16544 19717 16572
rect 19668 16532 19674 16544
rect 19705 16541 19717 16544
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 20622 16532 20628 16584
rect 20680 16572 20686 16584
rect 21008 16581 21036 16680
rect 21100 16680 22928 16708
rect 21100 16581 21128 16680
rect 22922 16668 22928 16680
rect 22980 16668 22986 16720
rect 23109 16643 23167 16649
rect 23109 16609 23121 16643
rect 23155 16640 23167 16643
rect 23216 16640 23244 16748
rect 26418 16736 26424 16748
rect 26476 16736 26482 16788
rect 27430 16736 27436 16788
rect 27488 16776 27494 16788
rect 27801 16779 27859 16785
rect 27801 16776 27813 16779
rect 27488 16748 27813 16776
rect 27488 16736 27494 16748
rect 27801 16745 27813 16748
rect 27847 16745 27859 16779
rect 27801 16739 27859 16745
rect 26786 16708 26792 16720
rect 25240 16680 26792 16708
rect 23155 16612 23244 16640
rect 23293 16643 23351 16649
rect 23155 16609 23167 16612
rect 23109 16603 23167 16609
rect 23293 16609 23305 16643
rect 23339 16640 23351 16643
rect 23750 16640 23756 16652
rect 23339 16612 23756 16640
rect 23339 16609 23351 16612
rect 23293 16603 23351 16609
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 25240 16649 25268 16680
rect 26786 16668 26792 16680
rect 26844 16668 26850 16720
rect 25225 16643 25283 16649
rect 25225 16609 25237 16643
rect 25271 16609 25283 16643
rect 25225 16603 25283 16609
rect 25409 16643 25467 16649
rect 25409 16609 25421 16643
rect 25455 16640 25467 16643
rect 26234 16640 26240 16652
rect 25455 16612 26240 16640
rect 25455 16609 25467 16612
rect 25409 16603 25467 16609
rect 26234 16600 26240 16612
rect 26292 16640 26298 16652
rect 27065 16643 27123 16649
rect 27065 16640 27077 16643
rect 26292 16612 27077 16640
rect 26292 16600 26298 16612
rect 27065 16609 27077 16612
rect 27111 16640 27123 16643
rect 27246 16640 27252 16652
rect 27111 16612 27252 16640
rect 27111 16609 27123 16612
rect 27065 16603 27123 16609
rect 27246 16600 27252 16612
rect 27304 16600 27310 16652
rect 27614 16640 27620 16652
rect 27527 16612 27620 16640
rect 27614 16600 27620 16612
rect 27672 16640 27678 16652
rect 28074 16640 28080 16652
rect 27672 16612 28080 16640
rect 27672 16600 27678 16612
rect 28074 16600 28080 16612
rect 28132 16600 28138 16652
rect 20809 16575 20867 16581
rect 20809 16572 20821 16575
rect 20680 16544 20821 16572
rect 20680 16532 20686 16544
rect 20809 16541 20821 16544
rect 20855 16541 20867 16575
rect 20809 16535 20867 16541
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 21085 16575 21143 16581
rect 21085 16541 21097 16575
rect 21131 16541 21143 16575
rect 21358 16572 21364 16584
rect 21319 16544 21364 16572
rect 21085 16535 21143 16541
rect 21358 16532 21364 16544
rect 21416 16572 21422 16584
rect 21821 16575 21879 16581
rect 21821 16572 21833 16575
rect 21416 16544 21833 16572
rect 21416 16532 21422 16544
rect 21821 16541 21833 16544
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 23017 16575 23075 16581
rect 23017 16541 23029 16575
rect 23063 16572 23075 16575
rect 23382 16572 23388 16584
rect 23063 16544 23388 16572
rect 23063 16541 23075 16544
rect 23017 16535 23075 16541
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 23566 16532 23572 16584
rect 23624 16572 23630 16584
rect 25133 16575 25191 16581
rect 25133 16572 25145 16575
rect 23624 16544 25145 16572
rect 23624 16532 23630 16544
rect 25133 16541 25145 16544
rect 25179 16541 25191 16575
rect 25133 16535 25191 16541
rect 25314 16532 25320 16584
rect 25372 16572 25378 16584
rect 25372 16544 26648 16572
rect 25372 16532 25378 16544
rect 14645 16507 14703 16513
rect 14645 16504 14657 16507
rect 13004 16476 14657 16504
rect 14645 16473 14657 16476
rect 14691 16504 14703 16507
rect 16482 16504 16488 16516
rect 14691 16476 16488 16504
rect 14691 16473 14703 16476
rect 14645 16467 14703 16473
rect 16482 16464 16488 16476
rect 16540 16464 16546 16516
rect 18598 16464 18604 16516
rect 18656 16504 18662 16516
rect 19242 16504 19248 16516
rect 18656 16476 19248 16504
rect 18656 16464 18662 16476
rect 19242 16464 19248 16476
rect 19300 16504 19306 16516
rect 22554 16504 22560 16516
rect 19300 16476 22560 16504
rect 19300 16464 19306 16476
rect 22554 16464 22560 16476
rect 22612 16464 22618 16516
rect 9661 16439 9719 16445
rect 9661 16405 9673 16439
rect 9707 16436 9719 16439
rect 10042 16436 10048 16448
rect 9707 16408 10048 16436
rect 9707 16405 9719 16408
rect 9661 16399 9719 16405
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 14277 16439 14335 16445
rect 14277 16436 14289 16439
rect 13872 16408 14289 16436
rect 13872 16396 13878 16408
rect 14277 16405 14289 16408
rect 14323 16436 14335 16439
rect 14550 16436 14556 16448
rect 14323 16408 14556 16436
rect 14323 16405 14335 16408
rect 14277 16399 14335 16405
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 14737 16439 14795 16445
rect 14737 16405 14749 16439
rect 14783 16436 14795 16439
rect 15194 16436 15200 16448
rect 14783 16408 15200 16436
rect 14783 16405 14795 16408
rect 14737 16399 14795 16405
rect 15194 16396 15200 16408
rect 15252 16436 15258 16448
rect 16390 16436 16396 16448
rect 15252 16408 16396 16436
rect 15252 16396 15258 16408
rect 16390 16396 16396 16408
rect 16448 16396 16454 16448
rect 17310 16396 17316 16448
rect 17368 16436 17374 16448
rect 17497 16439 17555 16445
rect 17497 16436 17509 16439
rect 17368 16408 17509 16436
rect 17368 16396 17374 16408
rect 17497 16405 17509 16408
rect 17543 16405 17555 16439
rect 17497 16399 17555 16405
rect 22094 16396 22100 16448
rect 22152 16436 22158 16448
rect 22649 16439 22707 16445
rect 22649 16436 22661 16439
rect 22152 16408 22661 16436
rect 22152 16396 22158 16408
rect 22649 16405 22661 16408
rect 22695 16405 22707 16439
rect 24762 16436 24768 16448
rect 24723 16408 24768 16436
rect 22649 16399 22707 16405
rect 24762 16396 24768 16408
rect 24820 16396 24826 16448
rect 26418 16436 26424 16448
rect 26379 16408 26424 16436
rect 26418 16396 26424 16408
rect 26476 16396 26482 16448
rect 26620 16436 26648 16544
rect 27430 16532 27436 16584
rect 27488 16572 27494 16584
rect 27893 16575 27951 16581
rect 27893 16572 27905 16575
rect 27488 16544 27905 16572
rect 27488 16532 27494 16544
rect 27893 16541 27905 16544
rect 27939 16541 27951 16575
rect 28718 16572 28724 16584
rect 28679 16544 28724 16572
rect 27893 16535 27951 16541
rect 28718 16532 28724 16544
rect 28776 16532 28782 16584
rect 26786 16504 26792 16516
rect 26747 16476 26792 16504
rect 26786 16464 26792 16476
rect 26844 16464 26850 16516
rect 26881 16507 26939 16513
rect 26881 16473 26893 16507
rect 26927 16504 26939 16507
rect 27338 16504 27344 16516
rect 26927 16476 27344 16504
rect 26927 16473 26939 16476
rect 26881 16467 26939 16473
rect 27338 16464 27344 16476
rect 27396 16504 27402 16516
rect 27617 16507 27675 16513
rect 27617 16504 27629 16507
rect 27396 16476 27629 16504
rect 27396 16464 27402 16476
rect 27617 16473 27629 16476
rect 27663 16473 27675 16507
rect 27617 16467 27675 16473
rect 28537 16439 28595 16445
rect 28537 16436 28549 16439
rect 26620 16408 28549 16436
rect 28537 16405 28549 16408
rect 28583 16405 28595 16439
rect 28537 16399 28595 16405
rect 1104 16346 29600 16368
rect 1104 16294 8034 16346
rect 8086 16294 8098 16346
rect 8150 16294 8162 16346
rect 8214 16294 8226 16346
rect 8278 16294 8290 16346
rect 8342 16294 15118 16346
rect 15170 16294 15182 16346
rect 15234 16294 15246 16346
rect 15298 16294 15310 16346
rect 15362 16294 15374 16346
rect 15426 16294 22202 16346
rect 22254 16294 22266 16346
rect 22318 16294 22330 16346
rect 22382 16294 22394 16346
rect 22446 16294 22458 16346
rect 22510 16294 29286 16346
rect 29338 16294 29350 16346
rect 29402 16294 29414 16346
rect 29466 16294 29478 16346
rect 29530 16294 29542 16346
rect 29594 16294 29600 16346
rect 1104 16272 29600 16294
rect 9030 16192 9036 16244
rect 9088 16232 9094 16244
rect 9217 16235 9275 16241
rect 9217 16232 9229 16235
rect 9088 16204 9229 16232
rect 9088 16192 9094 16204
rect 9217 16201 9229 16204
rect 9263 16232 9275 16235
rect 9858 16232 9864 16244
rect 9263 16204 9864 16232
rect 9263 16201 9275 16204
rect 9217 16195 9275 16201
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 10042 16232 10048 16244
rect 9955 16204 10048 16232
rect 10042 16192 10048 16204
rect 10100 16232 10106 16244
rect 10410 16232 10416 16244
rect 10100 16204 10416 16232
rect 10100 16192 10106 16204
rect 10410 16192 10416 16204
rect 10468 16232 10474 16244
rect 10962 16232 10968 16244
rect 10468 16204 10968 16232
rect 10468 16192 10474 16204
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 12584 16204 14596 16232
rect 12584 16192 12590 16204
rect 3786 16164 3792 16176
rect 3747 16136 3792 16164
rect 3786 16124 3792 16136
rect 3844 16124 3850 16176
rect 3970 16164 3976 16176
rect 3931 16136 3976 16164
rect 3970 16124 3976 16136
rect 4028 16124 4034 16176
rect 13170 16164 13176 16176
rect 12820 16136 13176 16164
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16096 1458 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 1452 16068 2053 16096
rect 1452 16056 1458 16068
rect 2041 16065 2053 16068
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 4062 16056 4068 16108
rect 4120 16096 4126 16108
rect 6730 16096 6736 16108
rect 4120 16068 4165 16096
rect 6691 16068 6736 16096
rect 4120 16056 4126 16068
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16096 6883 16099
rect 6914 16096 6920 16108
rect 6871 16068 6920 16096
rect 6871 16065 6883 16068
rect 6825 16059 6883 16065
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7009 16099 7067 16105
rect 7009 16065 7021 16099
rect 7055 16065 7067 16099
rect 7009 16059 7067 16065
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16065 7159 16099
rect 7101 16059 7159 16065
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16096 7619 16099
rect 7742 16096 7748 16108
rect 7607 16068 7748 16096
rect 7607 16065 7619 16068
rect 7561 16059 7619 16065
rect 5534 15988 5540 16040
rect 5592 16028 5598 16040
rect 7024 16028 7052 16059
rect 5592 16000 7052 16028
rect 7116 16028 7144 16059
rect 7742 16056 7748 16068
rect 7800 16056 7806 16108
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16096 11943 16099
rect 11974 16096 11980 16108
rect 11931 16068 11980 16096
rect 11931 16065 11943 16068
rect 11885 16059 11943 16065
rect 11974 16056 11980 16068
rect 12032 16056 12038 16108
rect 12069 16099 12127 16105
rect 12069 16065 12081 16099
rect 12115 16096 12127 16099
rect 12618 16096 12624 16108
rect 12115 16068 12624 16096
rect 12115 16065 12127 16068
rect 12069 16059 12127 16065
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 12820 16105 12848 16136
rect 13170 16124 13176 16136
rect 13228 16124 13234 16176
rect 14568 16164 14596 16204
rect 14918 16192 14924 16244
rect 14976 16232 14982 16244
rect 15105 16235 15163 16241
rect 15105 16232 15117 16235
rect 14976 16204 15117 16232
rect 14976 16192 14982 16204
rect 15105 16201 15117 16204
rect 15151 16232 15163 16235
rect 16206 16232 16212 16244
rect 15151 16204 16212 16232
rect 15151 16201 15163 16204
rect 15105 16195 15163 16201
rect 16206 16192 16212 16204
rect 16264 16192 16270 16244
rect 16574 16192 16580 16244
rect 16632 16232 16638 16244
rect 17129 16235 17187 16241
rect 17129 16232 17141 16235
rect 16632 16204 17141 16232
rect 16632 16192 16638 16204
rect 17129 16201 17141 16204
rect 17175 16201 17187 16235
rect 17129 16195 17187 16201
rect 18230 16192 18236 16244
rect 18288 16232 18294 16244
rect 20165 16235 20223 16241
rect 20165 16232 20177 16235
rect 18288 16204 20177 16232
rect 18288 16192 18294 16204
rect 20165 16201 20177 16204
rect 20211 16201 20223 16235
rect 20165 16195 20223 16201
rect 22833 16235 22891 16241
rect 22833 16201 22845 16235
rect 22879 16232 22891 16235
rect 22922 16232 22928 16244
rect 22879 16204 22928 16232
rect 22879 16201 22891 16204
rect 22833 16195 22891 16201
rect 22922 16192 22928 16204
rect 22980 16192 22986 16244
rect 23477 16235 23535 16241
rect 23477 16201 23489 16235
rect 23523 16232 23535 16235
rect 23658 16232 23664 16244
rect 23523 16204 23664 16232
rect 23523 16201 23535 16204
rect 23477 16195 23535 16201
rect 23658 16192 23664 16204
rect 23716 16192 23722 16244
rect 24026 16192 24032 16244
rect 24084 16232 24090 16244
rect 24121 16235 24179 16241
rect 24121 16232 24133 16235
rect 24084 16204 24133 16232
rect 24084 16192 24090 16204
rect 24121 16201 24133 16204
rect 24167 16201 24179 16235
rect 24121 16195 24179 16201
rect 24489 16235 24547 16241
rect 24489 16201 24501 16235
rect 24535 16232 24547 16235
rect 25038 16232 25044 16244
rect 24535 16204 25044 16232
rect 24535 16201 24547 16204
rect 24489 16195 24547 16201
rect 25038 16192 25044 16204
rect 25096 16192 25102 16244
rect 27062 16192 27068 16244
rect 27120 16232 27126 16244
rect 27341 16235 27399 16241
rect 27341 16232 27353 16235
rect 27120 16204 27353 16232
rect 27120 16192 27126 16204
rect 27341 16201 27353 16204
rect 27387 16201 27399 16235
rect 27341 16195 27399 16201
rect 15010 16164 15016 16176
rect 14568 16136 15016 16164
rect 15010 16124 15016 16136
rect 15068 16124 15074 16176
rect 17037 16167 17095 16173
rect 17037 16133 17049 16167
rect 17083 16164 17095 16167
rect 17218 16164 17224 16176
rect 17083 16136 17224 16164
rect 17083 16133 17095 16136
rect 17037 16127 17095 16133
rect 17218 16124 17224 16136
rect 17276 16124 17282 16176
rect 24762 16164 24768 16176
rect 18708 16136 24768 16164
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16065 12863 16099
rect 13262 16096 13268 16108
rect 12805 16059 12863 16065
rect 13004 16068 13268 16096
rect 12894 16028 12900 16040
rect 7116 16000 12900 16028
rect 5592 15988 5598 16000
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 7466 15960 7472 15972
rect 1627 15932 7472 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 7466 15920 7472 15932
rect 7524 15920 7530 15972
rect 7650 15960 7656 15972
rect 7611 15932 7656 15960
rect 7650 15920 7656 15932
rect 7708 15920 7714 15972
rect 7742 15920 7748 15972
rect 7800 15960 7806 15972
rect 8297 15963 8355 15969
rect 8297 15960 8309 15963
rect 7800 15932 8309 15960
rect 7800 15920 7806 15932
rect 8297 15929 8309 15932
rect 8343 15960 8355 15963
rect 10778 15960 10784 15972
rect 8343 15932 10784 15960
rect 8343 15929 8355 15932
rect 8297 15923 8355 15929
rect 10778 15920 10784 15932
rect 10836 15960 10842 15972
rect 12802 15960 12808 15972
rect 10836 15932 12808 15960
rect 10836 15920 10842 15932
rect 12802 15920 12808 15932
rect 12860 15920 12866 15972
rect 13004 15960 13032 16068
rect 13262 16056 13268 16068
rect 13320 16056 13326 16108
rect 13538 16056 13544 16108
rect 13596 16096 13602 16108
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 13596 16068 13737 16096
rect 13596 16056 13602 16068
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 13906 16096 13912 16108
rect 13867 16068 13912 16096
rect 13725 16059 13783 16065
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 15997 13139 16031
rect 13740 16028 13768 16059
rect 13906 16056 13912 16068
rect 13964 16056 13970 16108
rect 18414 16096 18420 16108
rect 15212 16068 18420 16096
rect 15212 16037 15240 16068
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 18598 16096 18604 16108
rect 18559 16068 18604 16096
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 18708 16105 18736 16136
rect 24762 16124 24768 16136
rect 24820 16124 24826 16176
rect 28169 16167 28227 16173
rect 28169 16133 28181 16167
rect 28215 16133 28227 16167
rect 28169 16127 28227 16133
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16065 18751 16099
rect 18693 16059 18751 16065
rect 18877 16099 18935 16105
rect 18877 16065 18889 16099
rect 18923 16096 18935 16099
rect 19058 16096 19064 16108
rect 18923 16068 19064 16096
rect 18923 16065 18935 16068
rect 18877 16059 18935 16065
rect 19058 16056 19064 16068
rect 19116 16096 19122 16108
rect 19337 16099 19395 16105
rect 19337 16096 19349 16099
rect 19116 16068 19349 16096
rect 19116 16056 19122 16068
rect 19337 16065 19349 16068
rect 19383 16065 19395 16099
rect 19337 16059 19395 16065
rect 20346 16056 20352 16108
rect 20404 16096 20410 16108
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 20404 16068 20545 16096
rect 20404 16056 20410 16068
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 21358 16056 21364 16108
rect 21416 16096 21422 16108
rect 22741 16099 22799 16105
rect 22741 16096 22753 16099
rect 21416 16068 22753 16096
rect 21416 16056 21422 16068
rect 22741 16065 22753 16068
rect 22787 16065 22799 16099
rect 22741 16059 22799 16065
rect 22925 16099 22983 16105
rect 22925 16065 22937 16099
rect 22971 16096 22983 16099
rect 23014 16096 23020 16108
rect 22971 16068 23020 16096
rect 22971 16065 22983 16068
rect 22925 16059 22983 16065
rect 15197 16031 15255 16037
rect 15197 16028 15209 16031
rect 13740 16000 15209 16028
rect 13081 15991 13139 15997
rect 15197 15997 15209 16000
rect 15243 15997 15255 16031
rect 17310 16028 17316 16040
rect 17271 16000 17316 16028
rect 15197 15991 15255 15997
rect 12912 15932 13032 15960
rect 13096 15960 13124 15991
rect 17310 15988 17316 16000
rect 17368 15988 17374 16040
rect 18138 15988 18144 16040
rect 18196 16028 18202 16040
rect 18233 16031 18291 16037
rect 18233 16028 18245 16031
rect 18196 16000 18245 16028
rect 18196 15988 18202 16000
rect 18233 15997 18245 16000
rect 18279 15997 18291 16031
rect 18233 15991 18291 15997
rect 18509 16031 18567 16037
rect 18509 15997 18521 16031
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 13541 15963 13599 15969
rect 13541 15960 13553 15963
rect 13096 15932 13553 15960
rect 4065 15895 4123 15901
rect 4065 15861 4077 15895
rect 4111 15892 4123 15895
rect 5258 15892 5264 15904
rect 4111 15864 5264 15892
rect 4111 15861 4123 15864
rect 4065 15855 4123 15861
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 6178 15852 6184 15904
rect 6236 15892 6242 15904
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 6236 15864 6561 15892
rect 6236 15852 6242 15864
rect 6549 15861 6561 15864
rect 6595 15861 6607 15895
rect 6549 15855 6607 15861
rect 11885 15895 11943 15901
rect 11885 15861 11897 15895
rect 11931 15892 11943 15895
rect 11974 15892 11980 15904
rect 11931 15864 11980 15892
rect 11931 15861 11943 15864
rect 11885 15855 11943 15861
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 12912 15901 12940 15932
rect 13541 15929 13553 15932
rect 13587 15929 13599 15963
rect 13541 15923 13599 15929
rect 14476 15932 15056 15960
rect 14476 15904 14504 15932
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15861 12955 15895
rect 12897 15855 12955 15861
rect 12986 15852 12992 15904
rect 13044 15892 13050 15904
rect 13909 15895 13967 15901
rect 13044 15864 13089 15892
rect 13044 15852 13050 15864
rect 13909 15861 13921 15895
rect 13955 15892 13967 15895
rect 14458 15892 14464 15904
rect 13955 15864 14464 15892
rect 13955 15861 13967 15864
rect 13909 15855 13967 15861
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 14642 15892 14648 15904
rect 14603 15864 14648 15892
rect 14642 15852 14648 15864
rect 14700 15852 14706 15904
rect 15028 15892 15056 15932
rect 16206 15920 16212 15972
rect 16264 15960 16270 15972
rect 16669 15963 16727 15969
rect 16669 15960 16681 15963
rect 16264 15932 16681 15960
rect 16264 15920 16270 15932
rect 16669 15929 16681 15932
rect 16715 15929 16727 15963
rect 18524 15960 18552 15991
rect 19150 15988 19156 16040
rect 19208 16028 19214 16040
rect 20625 16031 20683 16037
rect 19208 16000 19748 16028
rect 19208 15988 19214 16000
rect 19610 15960 19616 15972
rect 16669 15923 16727 15929
rect 18156 15932 19616 15960
rect 18156 15892 18184 15932
rect 19610 15920 19616 15932
rect 19668 15920 19674 15972
rect 15028 15864 18184 15892
rect 19720 15892 19748 16000
rect 20625 15997 20637 16031
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 20717 16031 20775 16037
rect 20717 15997 20729 16031
rect 20763 15997 20775 16031
rect 22756 16028 22784 16059
rect 23014 16056 23020 16068
rect 23072 16056 23078 16108
rect 24302 16056 24308 16108
rect 24360 16096 24366 16108
rect 27433 16099 27491 16105
rect 24360 16068 24716 16096
rect 24360 16056 24366 16068
rect 23658 16028 23664 16040
rect 22756 16000 23664 16028
rect 20717 15991 20775 15997
rect 20530 15920 20536 15972
rect 20588 15960 20594 15972
rect 20640 15960 20668 15991
rect 20588 15932 20668 15960
rect 20588 15920 20594 15932
rect 20732 15892 20760 15991
rect 23658 15988 23664 16000
rect 23716 15988 23722 16040
rect 24688 16037 24716 16068
rect 27433 16065 27445 16099
rect 27479 16096 27491 16099
rect 27706 16096 27712 16108
rect 27479 16068 27712 16096
rect 27479 16065 27491 16068
rect 27433 16059 27491 16065
rect 27706 16056 27712 16068
rect 27764 16096 27770 16108
rect 28184 16096 28212 16127
rect 28350 16096 28356 16108
rect 27764 16068 28212 16096
rect 28311 16068 28356 16096
rect 27764 16056 27770 16068
rect 28350 16056 28356 16068
rect 28408 16056 28414 16108
rect 28445 16099 28503 16105
rect 28445 16065 28457 16099
rect 28491 16065 28503 16099
rect 28445 16059 28503 16065
rect 24581 16031 24639 16037
rect 24581 15997 24593 16031
rect 24627 15997 24639 16031
rect 24581 15991 24639 15997
rect 24673 16031 24731 16037
rect 24673 15997 24685 16031
rect 24719 15997 24731 16031
rect 24673 15991 24731 15997
rect 24596 15960 24624 15991
rect 27246 15988 27252 16040
rect 27304 16028 27310 16040
rect 27525 16031 27583 16037
rect 27525 16028 27537 16031
rect 27304 16000 27537 16028
rect 27304 15988 27310 16000
rect 27525 15997 27537 16000
rect 27571 15997 27583 16031
rect 27525 15991 27583 15997
rect 28074 15988 28080 16040
rect 28132 16028 28138 16040
rect 28169 16031 28227 16037
rect 28169 16028 28181 16031
rect 28132 16000 28181 16028
rect 28132 15988 28138 16000
rect 28169 15997 28181 16000
rect 28215 15997 28227 16031
rect 28169 15991 28227 15997
rect 28258 15988 28264 16040
rect 28316 16028 28322 16040
rect 28460 16028 28488 16059
rect 28316 16000 28488 16028
rect 28316 15988 28322 16000
rect 24596 15932 25452 15960
rect 25424 15904 25452 15932
rect 21821 15895 21879 15901
rect 21821 15892 21833 15895
rect 19720 15864 21833 15892
rect 21821 15861 21833 15864
rect 21867 15861 21879 15895
rect 21821 15855 21879 15861
rect 25406 15852 25412 15904
rect 25464 15892 25470 15904
rect 26973 15895 27031 15901
rect 26973 15892 26985 15895
rect 25464 15864 26985 15892
rect 25464 15852 25470 15864
rect 26973 15861 26985 15864
rect 27019 15861 27031 15895
rect 26973 15855 27031 15861
rect 1104 15802 29440 15824
rect 1104 15750 4492 15802
rect 4544 15750 4556 15802
rect 4608 15750 4620 15802
rect 4672 15750 4684 15802
rect 4736 15750 4748 15802
rect 4800 15750 11576 15802
rect 11628 15750 11640 15802
rect 11692 15750 11704 15802
rect 11756 15750 11768 15802
rect 11820 15750 11832 15802
rect 11884 15750 18660 15802
rect 18712 15750 18724 15802
rect 18776 15750 18788 15802
rect 18840 15750 18852 15802
rect 18904 15750 18916 15802
rect 18968 15750 25744 15802
rect 25796 15750 25808 15802
rect 25860 15750 25872 15802
rect 25924 15750 25936 15802
rect 25988 15750 26000 15802
rect 26052 15750 29440 15802
rect 1104 15728 29440 15750
rect 4614 15648 4620 15700
rect 4672 15688 4678 15700
rect 4801 15691 4859 15697
rect 4801 15688 4813 15691
rect 4672 15660 4813 15688
rect 4672 15648 4678 15660
rect 4801 15657 4813 15660
rect 4847 15688 4859 15691
rect 5166 15688 5172 15700
rect 4847 15660 5172 15688
rect 4847 15657 4859 15660
rect 4801 15651 4859 15657
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 5626 15688 5632 15700
rect 5587 15660 5632 15688
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 9732 15660 10149 15688
rect 9732 15648 9738 15660
rect 10137 15657 10149 15660
rect 10183 15657 10195 15691
rect 16390 15688 16396 15700
rect 16351 15660 16396 15688
rect 10137 15651 10195 15657
rect 16390 15648 16396 15660
rect 16448 15648 16454 15700
rect 16482 15648 16488 15700
rect 16540 15688 16546 15700
rect 17865 15691 17923 15697
rect 17865 15688 17877 15691
rect 16540 15660 17877 15688
rect 16540 15648 16546 15660
rect 17865 15657 17877 15660
rect 17911 15657 17923 15691
rect 17865 15651 17923 15657
rect 19610 15648 19616 15700
rect 19668 15688 19674 15700
rect 19886 15688 19892 15700
rect 19668 15660 19892 15688
rect 19668 15648 19674 15660
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20254 15648 20260 15700
rect 20312 15688 20318 15700
rect 20349 15691 20407 15697
rect 20349 15688 20361 15691
rect 20312 15660 20361 15688
rect 20312 15648 20318 15660
rect 20349 15657 20361 15660
rect 20395 15657 20407 15691
rect 20349 15651 20407 15657
rect 22465 15691 22523 15697
rect 22465 15657 22477 15691
rect 22511 15688 22523 15691
rect 23014 15688 23020 15700
rect 22511 15660 23020 15688
rect 22511 15657 22523 15660
rect 22465 15651 22523 15657
rect 23014 15648 23020 15660
rect 23072 15648 23078 15700
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 23477 15691 23535 15697
rect 23477 15688 23489 15691
rect 23440 15660 23489 15688
rect 23440 15648 23446 15660
rect 23477 15657 23489 15660
rect 23523 15657 23535 15691
rect 28718 15688 28724 15700
rect 28679 15660 28724 15688
rect 23477 15651 23535 15657
rect 28718 15648 28724 15660
rect 28776 15648 28782 15700
rect 15289 15623 15347 15629
rect 15289 15589 15301 15623
rect 15335 15620 15347 15623
rect 15562 15620 15568 15632
rect 15335 15592 15568 15620
rect 15335 15589 15347 15592
rect 15289 15583 15347 15589
rect 15562 15580 15568 15592
rect 15620 15580 15626 15632
rect 18046 15620 18052 15632
rect 17052 15592 18052 15620
rect 6178 15552 6184 15564
rect 6139 15524 6184 15552
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 14642 15512 14648 15564
rect 14700 15552 14706 15564
rect 17052 15561 17080 15592
rect 18046 15580 18052 15592
rect 18104 15580 18110 15632
rect 15381 15555 15439 15561
rect 15381 15552 15393 15555
rect 14700 15524 15393 15552
rect 14700 15512 14706 15524
rect 15381 15521 15393 15524
rect 15427 15521 15439 15555
rect 15381 15515 15439 15521
rect 17037 15555 17095 15561
rect 17037 15521 17049 15555
rect 17083 15521 17095 15555
rect 23032 15552 23060 15648
rect 24578 15580 24584 15632
rect 24636 15580 24642 15632
rect 23382 15552 23388 15564
rect 23032 15524 23388 15552
rect 17037 15515 17095 15521
rect 23382 15512 23388 15524
rect 23440 15512 23446 15564
rect 23934 15512 23940 15564
rect 23992 15552 23998 15564
rect 24596 15552 24624 15580
rect 25869 15555 25927 15561
rect 25869 15552 25881 15555
rect 23992 15524 25881 15552
rect 23992 15512 23998 15524
rect 3786 15484 3792 15496
rect 3747 15456 3792 15484
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 4062 15484 4068 15496
rect 4023 15456 4068 15484
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 6454 15484 6460 15496
rect 6415 15456 6460 15484
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 10686 15444 10692 15496
rect 10744 15484 10750 15496
rect 11241 15487 11299 15493
rect 11241 15484 11253 15487
rect 10744 15456 11253 15484
rect 10744 15444 10750 15456
rect 11241 15453 11253 15456
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 15197 15487 15255 15493
rect 15197 15453 15209 15487
rect 15243 15453 15255 15487
rect 15470 15484 15476 15496
rect 15431 15456 15476 15484
rect 15197 15447 15255 15453
rect 3881 15419 3939 15425
rect 3881 15385 3893 15419
rect 3927 15416 3939 15419
rect 3970 15416 3976 15428
rect 3927 15388 3976 15416
rect 3927 15385 3939 15388
rect 3881 15379 3939 15385
rect 3970 15376 3976 15388
rect 4028 15376 4034 15428
rect 4249 15419 4307 15425
rect 4249 15385 4261 15419
rect 4295 15416 4307 15419
rect 5166 15416 5172 15428
rect 4295 15388 5172 15416
rect 4295 15385 4307 15388
rect 4249 15379 4307 15385
rect 5166 15376 5172 15388
rect 5224 15376 5230 15428
rect 15212 15416 15240 15447
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 16666 15484 16672 15496
rect 15580 15456 16672 15484
rect 15580 15416 15608 15456
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 16761 15487 16819 15493
rect 16761 15453 16773 15487
rect 16807 15484 16819 15487
rect 17402 15484 17408 15496
rect 16807 15456 17408 15484
rect 16807 15453 16819 15456
rect 16761 15447 16819 15453
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15484 18107 15487
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 18095 15456 19257 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 19245 15453 19257 15456
rect 19291 15484 19303 15487
rect 21358 15484 21364 15496
rect 19291 15456 21364 15484
rect 19291 15453 19303 15456
rect 19245 15447 19303 15453
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15484 24639 15487
rect 25038 15484 25044 15496
rect 24627 15456 25044 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 25038 15444 25044 15456
rect 25096 15444 25102 15496
rect 25240 15493 25268 15524
rect 25869 15521 25881 15524
rect 25915 15521 25927 15555
rect 25869 15515 25927 15521
rect 25225 15487 25283 15493
rect 25225 15453 25237 15487
rect 25271 15453 25283 15487
rect 25406 15484 25412 15496
rect 25367 15456 25412 15484
rect 25225 15447 25283 15453
rect 25406 15444 25412 15456
rect 25464 15444 25470 15496
rect 27246 15484 27252 15496
rect 27207 15456 27252 15484
rect 27246 15444 27252 15456
rect 27304 15444 27310 15496
rect 15212 15388 15608 15416
rect 15657 15419 15715 15425
rect 15657 15385 15669 15419
rect 15703 15416 15715 15419
rect 17954 15416 17960 15428
rect 15703 15388 17960 15416
rect 15703 15385 15715 15388
rect 15657 15379 15715 15385
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 18230 15416 18236 15428
rect 18191 15388 18236 15416
rect 18230 15376 18236 15388
rect 18288 15376 18294 15428
rect 9306 15308 9312 15360
rect 9364 15348 9370 15360
rect 10689 15351 10747 15357
rect 10689 15348 10701 15351
rect 9364 15320 10701 15348
rect 9364 15308 9370 15320
rect 10689 15317 10701 15320
rect 10735 15317 10747 15351
rect 12158 15348 12164 15360
rect 12119 15320 12164 15348
rect 10689 15311 10747 15317
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 13906 15308 13912 15360
rect 13964 15348 13970 15360
rect 15010 15348 15016 15360
rect 13964 15320 15016 15348
rect 13964 15308 13970 15320
rect 15010 15308 15016 15320
rect 15068 15348 15074 15360
rect 16758 15348 16764 15360
rect 15068 15320 16764 15348
rect 15068 15308 15074 15320
rect 16758 15308 16764 15320
rect 16816 15308 16822 15360
rect 16853 15351 16911 15357
rect 16853 15317 16865 15351
rect 16899 15348 16911 15351
rect 17218 15348 17224 15360
rect 16899 15320 17224 15348
rect 16899 15317 16911 15320
rect 16853 15311 16911 15317
rect 17218 15308 17224 15320
rect 17276 15308 17282 15360
rect 19058 15308 19064 15360
rect 19116 15348 19122 15360
rect 23934 15348 23940 15360
rect 19116 15320 23940 15348
rect 19116 15308 19122 15320
rect 23934 15308 23940 15320
rect 23992 15308 23998 15360
rect 24578 15308 24584 15360
rect 24636 15348 24642 15360
rect 24673 15351 24731 15357
rect 24673 15348 24685 15351
rect 24636 15320 24685 15348
rect 24636 15308 24642 15320
rect 24673 15317 24685 15320
rect 24719 15317 24731 15351
rect 24673 15311 24731 15317
rect 24854 15308 24860 15360
rect 24912 15348 24918 15360
rect 25225 15351 25283 15357
rect 25225 15348 25237 15351
rect 24912 15320 25237 15348
rect 24912 15308 24918 15320
rect 25225 15317 25237 15320
rect 25271 15317 25283 15351
rect 27522 15348 27528 15360
rect 27483 15320 27528 15348
rect 25225 15311 25283 15317
rect 27522 15308 27528 15320
rect 27580 15308 27586 15360
rect 1104 15258 29600 15280
rect 1104 15206 8034 15258
rect 8086 15206 8098 15258
rect 8150 15206 8162 15258
rect 8214 15206 8226 15258
rect 8278 15206 8290 15258
rect 8342 15206 15118 15258
rect 15170 15206 15182 15258
rect 15234 15206 15246 15258
rect 15298 15206 15310 15258
rect 15362 15206 15374 15258
rect 15426 15206 22202 15258
rect 22254 15206 22266 15258
rect 22318 15206 22330 15258
rect 22382 15206 22394 15258
rect 22446 15206 22458 15258
rect 22510 15206 29286 15258
rect 29338 15206 29350 15258
rect 29402 15206 29414 15258
rect 29466 15206 29478 15258
rect 29530 15206 29542 15258
rect 29594 15206 29600 15258
rect 1104 15184 29600 15206
rect 3789 15147 3847 15153
rect 3789 15113 3801 15147
rect 3835 15144 3847 15147
rect 4062 15144 4068 15156
rect 3835 15116 4068 15144
rect 3835 15113 3847 15116
rect 3789 15107 3847 15113
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 5445 15147 5503 15153
rect 5092 15116 5396 15144
rect 5092 15085 5120 15116
rect 5077 15079 5135 15085
rect 5077 15045 5089 15079
rect 5123 15045 5135 15079
rect 5077 15039 5135 15045
rect 5166 15036 5172 15088
rect 5224 15076 5230 15088
rect 5277 15079 5335 15085
rect 5277 15076 5289 15079
rect 5224 15048 5289 15076
rect 5224 15036 5230 15048
rect 5277 15045 5289 15048
rect 5323 15045 5335 15079
rect 5368 15076 5396 15116
rect 5445 15113 5457 15147
rect 5491 15144 5503 15147
rect 5534 15144 5540 15156
rect 5491 15116 5540 15144
rect 5491 15113 5503 15116
rect 5445 15107 5503 15113
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 6457 15147 6515 15153
rect 6457 15113 6469 15147
rect 6503 15144 6515 15147
rect 6730 15144 6736 15156
rect 6503 15116 6736 15144
rect 6503 15113 6515 15116
rect 6457 15107 6515 15113
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 9674 15104 9680 15156
rect 9732 15104 9738 15156
rect 11885 15147 11943 15153
rect 11885 15113 11897 15147
rect 11931 15144 11943 15147
rect 11974 15144 11980 15156
rect 11931 15116 11980 15144
rect 11931 15113 11943 15116
rect 11885 15107 11943 15113
rect 11974 15104 11980 15116
rect 12032 15104 12038 15156
rect 13446 15104 13452 15156
rect 13504 15144 13510 15156
rect 16758 15144 16764 15156
rect 13504 15116 14412 15144
rect 16719 15116 16764 15144
rect 13504 15104 13510 15116
rect 5626 15076 5632 15088
rect 5368 15048 5632 15076
rect 5277 15039 5335 15045
rect 5626 15036 5632 15048
rect 5684 15036 5690 15088
rect 7466 15036 7472 15088
rect 7524 15076 7530 15088
rect 7561 15079 7619 15085
rect 7561 15076 7573 15079
rect 7524 15048 7573 15076
rect 7524 15036 7530 15048
rect 7561 15045 7573 15048
rect 7607 15045 7619 15079
rect 9692 15076 9720 15104
rect 9766 15076 9772 15088
rect 9679 15048 9772 15076
rect 7561 15039 7619 15045
rect 9766 15036 9772 15048
rect 9824 15076 9830 15088
rect 9861 15079 9919 15085
rect 9861 15076 9873 15079
rect 9824 15048 9873 15076
rect 9824 15036 9830 15048
rect 9861 15045 9873 15048
rect 9907 15045 9919 15079
rect 9861 15039 9919 15045
rect 12894 15036 12900 15088
rect 12952 15076 12958 15088
rect 13633 15079 13691 15085
rect 13633 15076 13645 15079
rect 12952 15048 13645 15076
rect 12952 15036 12958 15048
rect 13633 15045 13645 15048
rect 13679 15045 13691 15079
rect 13633 15039 13691 15045
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 15008 3847 15011
rect 4338 15008 4344 15020
rect 3835 14980 4344 15008
rect 3835 14977 3847 14980
rect 3789 14971 3847 14977
rect 3620 14940 3648 14971
rect 4338 14968 4344 14980
rect 4396 14968 4402 15020
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 15008 4675 15011
rect 6825 15011 6883 15017
rect 6825 15008 6837 15011
rect 4663 14980 6837 15008
rect 4663 14977 4675 14980
rect 4617 14971 4675 14977
rect 6825 14977 6837 14980
rect 6871 15008 6883 15011
rect 7098 15008 7104 15020
rect 6871 14980 7104 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 7929 15011 7987 15017
rect 7929 14977 7941 15011
rect 7975 15008 7987 15011
rect 9122 15008 9128 15020
rect 7975 14980 9128 15008
rect 7975 14977 7987 14980
rect 7929 14971 7987 14977
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 9674 15008 9680 15020
rect 9635 14980 9680 15008
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 9953 15011 10011 15017
rect 9953 14977 9965 15011
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 10091 14980 10180 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 4525 14943 4583 14949
rect 3620 14912 4292 14940
rect 4264 14881 4292 14912
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 4890 14940 4896 14952
rect 4571 14912 4896 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14909 6975 14943
rect 9968 14940 9996 14971
rect 6917 14903 6975 14909
rect 9646 14912 9996 14940
rect 4249 14875 4307 14881
rect 4249 14841 4261 14875
rect 4295 14841 4307 14875
rect 5350 14872 5356 14884
rect 4249 14835 4307 14841
rect 4632 14844 5356 14872
rect 4632 14816 4660 14844
rect 5350 14832 5356 14844
rect 5408 14832 5414 14884
rect 6932 14872 6960 14903
rect 7558 14872 7564 14884
rect 6932 14844 7564 14872
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 4614 14804 4620 14816
rect 4575 14776 4620 14804
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 5074 14764 5080 14816
rect 5132 14804 5138 14816
rect 5258 14804 5264 14816
rect 5132 14776 5264 14804
rect 5132 14764 5138 14776
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 9217 14807 9275 14813
rect 9217 14773 9229 14807
rect 9263 14804 9275 14807
rect 9306 14804 9312 14816
rect 9263 14776 9312 14804
rect 9263 14773 9275 14776
rect 9217 14767 9275 14773
rect 9306 14764 9312 14776
rect 9364 14804 9370 14816
rect 9646 14804 9674 14912
rect 10152 14872 10180 14980
rect 10594 14968 10600 15020
rect 10652 15008 10658 15020
rect 10689 15011 10747 15017
rect 10689 15008 10701 15011
rect 10652 14980 10701 15008
rect 10652 14968 10658 14980
rect 10689 14977 10701 14980
rect 10735 14977 10747 15011
rect 10689 14971 10747 14977
rect 10781 15011 10839 15017
rect 10781 14977 10793 15011
rect 10827 14977 10839 15011
rect 10781 14971 10839 14977
rect 10226 14900 10232 14952
rect 10284 14940 10290 14952
rect 10796 14940 10824 14971
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10928 14980 10977 15008
rect 10928 14968 10934 14980
rect 10965 14977 10977 14980
rect 11011 14977 11023 15011
rect 10965 14971 11023 14977
rect 11422 14968 11428 15020
rect 11480 15008 11486 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11480 14980 11713 15008
rect 11480 14968 11486 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 15008 12035 15011
rect 12986 15008 12992 15020
rect 12023 14980 12992 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12986 14968 12992 14980
rect 13044 14968 13050 15020
rect 13538 15008 13544 15020
rect 13499 14980 13544 15008
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 13998 15008 14004 15020
rect 13959 14980 14004 15008
rect 13998 14968 14004 14980
rect 14056 14968 14062 15020
rect 14384 15017 14412 15116
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 17129 15147 17187 15153
rect 17129 15113 17141 15147
rect 17175 15144 17187 15147
rect 18230 15144 18236 15156
rect 17175 15116 18236 15144
rect 17175 15113 17187 15116
rect 17129 15107 17187 15113
rect 18230 15104 18236 15116
rect 18288 15104 18294 15156
rect 21266 15144 21272 15156
rect 20732 15116 21272 15144
rect 15105 15079 15163 15085
rect 15105 15045 15117 15079
rect 15151 15076 15163 15079
rect 17586 15076 17592 15088
rect 15151 15048 17592 15076
rect 15151 15045 15163 15048
rect 15105 15039 15163 15045
rect 14369 15011 14427 15017
rect 14369 14977 14381 15011
rect 14415 14977 14427 15011
rect 14369 14971 14427 14977
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 15008 14611 15011
rect 14642 15008 14648 15020
rect 14599 14980 14648 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 14642 14968 14648 14980
rect 14700 14968 14706 15020
rect 10284 14912 10824 14940
rect 10284 14900 10290 14912
rect 12158 14900 12164 14952
rect 12216 14940 12222 14952
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 12216 14912 14105 14940
rect 12216 14900 12222 14912
rect 14093 14909 14105 14912
rect 14139 14940 14151 14943
rect 15120 14940 15148 15039
rect 17586 15036 17592 15048
rect 17644 15036 17650 15088
rect 20073 15079 20131 15085
rect 20073 15045 20085 15079
rect 20119 15076 20131 15079
rect 20732 15076 20760 15116
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 24489 15147 24547 15153
rect 24489 15113 24501 15147
rect 24535 15144 24547 15147
rect 24762 15144 24768 15156
rect 24535 15116 24768 15144
rect 24535 15113 24547 15116
rect 24489 15107 24547 15113
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 27338 15144 27344 15156
rect 27299 15116 27344 15144
rect 27338 15104 27344 15116
rect 27396 15104 27402 15156
rect 20119 15048 20760 15076
rect 20119 15045 20131 15048
rect 20073 15039 20131 15045
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17402 15008 17408 15020
rect 17267 14980 17408 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 17402 14968 17408 14980
rect 17460 14968 17466 15020
rect 17954 15008 17960 15020
rect 17915 14980 17960 15008
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 15008 18291 15011
rect 18414 15008 18420 15020
rect 18279 14980 18420 15008
rect 18279 14977 18291 14980
rect 18233 14971 18291 14977
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 20254 14968 20260 15020
rect 20312 15008 20318 15020
rect 20732 15017 20760 15048
rect 20806 15036 20812 15088
rect 20864 15076 20870 15088
rect 20864 15048 20944 15076
rect 20864 15036 20870 15048
rect 20916 15017 20944 15048
rect 20625 15011 20683 15017
rect 20625 15008 20637 15011
rect 20312 14980 20637 15008
rect 20312 14968 20318 14980
rect 20625 14977 20637 14980
rect 20671 14977 20683 15011
rect 20625 14971 20683 14977
rect 20717 15011 20775 15017
rect 20717 14977 20729 15011
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 15008 20959 15011
rect 21634 15008 21640 15020
rect 20947 14980 21640 15008
rect 20947 14977 20959 14980
rect 20901 14971 20959 14977
rect 21634 14968 21640 14980
rect 21692 14968 21698 15020
rect 24302 14968 24308 15020
rect 24360 15008 24366 15020
rect 24360 14980 24716 15008
rect 24360 14968 24366 14980
rect 17310 14940 17316 14952
rect 14139 14912 15148 14940
rect 17223 14912 17316 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 17310 14900 17316 14912
rect 17368 14940 17374 14952
rect 18785 14943 18843 14949
rect 18785 14940 18797 14943
rect 17368 14912 18797 14940
rect 17368 14900 17374 14912
rect 18785 14909 18797 14912
rect 18831 14909 18843 14943
rect 18785 14903 18843 14909
rect 20809 14943 20867 14949
rect 20809 14909 20821 14943
rect 20855 14909 20867 14943
rect 21082 14940 21088 14952
rect 21043 14912 21088 14940
rect 20809 14903 20867 14909
rect 10686 14872 10692 14884
rect 10152 14844 10692 14872
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 18046 14872 18052 14884
rect 18007 14844 18052 14872
rect 18046 14832 18052 14844
rect 18104 14832 18110 14884
rect 20622 14832 20628 14884
rect 20680 14872 20686 14884
rect 20824 14872 20852 14903
rect 21082 14900 21088 14912
rect 21140 14900 21146 14952
rect 24688 14949 24716 14980
rect 27338 14968 27344 15020
rect 27396 15008 27402 15020
rect 28169 15011 28227 15017
rect 28169 15008 28181 15011
rect 27396 14980 28181 15008
rect 27396 14968 27402 14980
rect 28169 14977 28181 14980
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 24581 14943 24639 14949
rect 24581 14909 24593 14943
rect 24627 14909 24639 14943
rect 24581 14903 24639 14909
rect 24673 14943 24731 14949
rect 24673 14909 24685 14943
rect 24719 14940 24731 14943
rect 25498 14940 25504 14952
rect 24719 14912 25504 14940
rect 24719 14909 24731 14912
rect 24673 14903 24731 14909
rect 24302 14872 24308 14884
rect 20680 14844 20852 14872
rect 21008 14844 24308 14872
rect 20680 14832 20686 14844
rect 9364 14776 9674 14804
rect 9364 14764 9370 14776
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 10229 14807 10287 14813
rect 10229 14804 10241 14807
rect 10192 14776 10241 14804
rect 10192 14764 10198 14776
rect 10229 14773 10241 14776
rect 10275 14773 10287 14807
rect 10962 14804 10968 14816
rect 10923 14776 10968 14804
rect 10229 14767 10287 14773
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 11517 14807 11575 14813
rect 11517 14804 11529 14807
rect 11388 14776 11529 14804
rect 11388 14764 11394 14776
rect 11517 14773 11529 14776
rect 11563 14773 11575 14807
rect 11517 14767 11575 14773
rect 15654 14764 15660 14816
rect 15712 14804 15718 14816
rect 16298 14804 16304 14816
rect 15712 14776 16304 14804
rect 15712 14764 15718 14776
rect 16298 14764 16304 14776
rect 16356 14804 16362 14816
rect 21008 14804 21036 14844
rect 24302 14832 24308 14844
rect 24360 14832 24366 14884
rect 24596 14872 24624 14903
rect 25498 14900 25504 14912
rect 25556 14900 25562 14952
rect 27430 14940 27436 14952
rect 27391 14912 27436 14940
rect 27430 14900 27436 14912
rect 27488 14900 27494 14952
rect 27522 14900 27528 14952
rect 27580 14940 27586 14952
rect 27580 14912 27625 14940
rect 27580 14900 27586 14912
rect 25222 14872 25228 14884
rect 24596 14844 25228 14872
rect 25222 14832 25228 14844
rect 25280 14872 25286 14884
rect 26973 14875 27031 14881
rect 26973 14872 26985 14875
rect 25280 14844 26985 14872
rect 25280 14832 25286 14844
rect 26973 14841 26985 14844
rect 27019 14841 27031 14875
rect 26973 14835 27031 14841
rect 16356 14776 21036 14804
rect 16356 14764 16362 14776
rect 23566 14764 23572 14816
rect 23624 14804 23630 14816
rect 24121 14807 24179 14813
rect 24121 14804 24133 14807
rect 23624 14776 24133 14804
rect 23624 14764 23630 14776
rect 24121 14773 24133 14776
rect 24167 14773 24179 14807
rect 24121 14767 24179 14773
rect 28258 14764 28264 14816
rect 28316 14804 28322 14816
rect 28353 14807 28411 14813
rect 28353 14804 28365 14807
rect 28316 14776 28365 14804
rect 28316 14764 28322 14776
rect 28353 14773 28365 14776
rect 28399 14773 28411 14807
rect 28353 14767 28411 14773
rect 1104 14714 29440 14736
rect 1104 14662 4492 14714
rect 4544 14662 4556 14714
rect 4608 14662 4620 14714
rect 4672 14662 4684 14714
rect 4736 14662 4748 14714
rect 4800 14662 11576 14714
rect 11628 14662 11640 14714
rect 11692 14662 11704 14714
rect 11756 14662 11768 14714
rect 11820 14662 11832 14714
rect 11884 14662 18660 14714
rect 18712 14662 18724 14714
rect 18776 14662 18788 14714
rect 18840 14662 18852 14714
rect 18904 14662 18916 14714
rect 18968 14662 25744 14714
rect 25796 14662 25808 14714
rect 25860 14662 25872 14714
rect 25924 14662 25936 14714
rect 25988 14662 26000 14714
rect 26052 14662 29440 14714
rect 1104 14640 29440 14662
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 4982 14600 4988 14612
rect 4396 14572 4988 14600
rect 4396 14560 4402 14572
rect 4982 14560 4988 14572
rect 5040 14600 5046 14612
rect 5261 14603 5319 14609
rect 5261 14600 5273 14603
rect 5040 14572 5273 14600
rect 5040 14560 5046 14572
rect 5261 14569 5273 14572
rect 5307 14569 5319 14603
rect 5261 14563 5319 14569
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 6914 14600 6920 14612
rect 6595 14572 6920 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 7558 14600 7564 14612
rect 7423 14572 7564 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 7558 14560 7564 14572
rect 7616 14560 7622 14612
rect 9490 14600 9496 14612
rect 9403 14572 9496 14600
rect 9490 14560 9496 14572
rect 9548 14600 9554 14612
rect 10226 14600 10232 14612
rect 9548 14572 10232 14600
rect 9548 14560 9554 14572
rect 10226 14560 10232 14572
rect 10284 14560 10290 14612
rect 10689 14603 10747 14609
rect 10689 14569 10701 14603
rect 10735 14600 10747 14603
rect 10870 14600 10876 14612
rect 10735 14572 10876 14600
rect 10735 14569 10747 14572
rect 10689 14563 10747 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13596 14572 14105 14600
rect 13596 14560 13602 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 14093 14563 14151 14569
rect 18233 14603 18291 14609
rect 18233 14569 18245 14603
rect 18279 14569 18291 14603
rect 18414 14600 18420 14612
rect 18375 14572 18420 14600
rect 18233 14563 18291 14569
rect 6822 14532 6828 14544
rect 2240 14504 6828 14532
rect 2240 14473 2268 14504
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 14369 14535 14427 14541
rect 14369 14501 14381 14535
rect 14415 14532 14427 14535
rect 18248 14532 18276 14563
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 19242 14560 19248 14612
rect 19300 14600 19306 14612
rect 19705 14603 19763 14609
rect 19705 14600 19717 14603
rect 19300 14572 19717 14600
rect 19300 14560 19306 14572
rect 19705 14569 19717 14572
rect 19751 14569 19763 14603
rect 19705 14563 19763 14569
rect 19797 14603 19855 14609
rect 19797 14569 19809 14603
rect 19843 14600 19855 14603
rect 21545 14603 21603 14609
rect 21545 14600 21557 14603
rect 19843 14572 21557 14600
rect 19843 14569 19855 14572
rect 19797 14563 19855 14569
rect 21545 14569 21557 14572
rect 21591 14569 21603 14603
rect 21545 14563 21603 14569
rect 23201 14603 23259 14609
rect 23201 14569 23213 14603
rect 23247 14600 23259 14603
rect 23934 14600 23940 14612
rect 23247 14572 23940 14600
rect 23247 14569 23259 14572
rect 23201 14563 23259 14569
rect 23934 14560 23940 14572
rect 23992 14560 23998 14612
rect 24302 14560 24308 14612
rect 24360 14600 24366 14612
rect 26142 14600 26148 14612
rect 24360 14572 26148 14600
rect 24360 14560 24366 14572
rect 26142 14560 26148 14572
rect 26200 14600 26206 14612
rect 26881 14603 26939 14609
rect 26881 14600 26893 14603
rect 26200 14572 26893 14600
rect 26200 14560 26206 14572
rect 26881 14569 26893 14572
rect 26927 14600 26939 14603
rect 27798 14600 27804 14612
rect 26927 14572 27804 14600
rect 26927 14569 26939 14572
rect 26881 14563 26939 14569
rect 27798 14560 27804 14572
rect 27856 14560 27862 14612
rect 19260 14532 19288 14560
rect 22738 14532 22744 14544
rect 14415 14504 19288 14532
rect 20640 14504 22744 14532
rect 14415 14501 14427 14504
rect 14369 14495 14427 14501
rect 20640 14476 20668 14504
rect 22738 14492 22744 14504
rect 22796 14492 22802 14544
rect 27338 14532 27344 14544
rect 23676 14504 27344 14532
rect 2225 14467 2283 14473
rect 2225 14433 2237 14467
rect 2271 14433 2283 14467
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 2225 14427 2283 14433
rect 4356 14436 5365 14464
rect 2130 14396 2136 14408
rect 2091 14368 2136 14396
rect 2130 14356 2136 14368
rect 2188 14396 2194 14408
rect 4356 14405 4384 14436
rect 5353 14433 5365 14436
rect 5399 14464 5411 14467
rect 5399 14436 7144 14464
rect 5399 14433 5411 14436
rect 5353 14427 5411 14433
rect 7116 14408 7144 14436
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 9640 14436 10456 14464
rect 9640 14424 9646 14436
rect 4341 14399 4399 14405
rect 2188 14368 2774 14396
rect 2188 14356 2194 14368
rect 2746 14328 2774 14368
rect 4341 14365 4353 14399
rect 4387 14365 4399 14399
rect 4522 14396 4528 14408
rect 4483 14368 4528 14396
rect 4341 14359 4399 14365
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 4890 14396 4896 14408
rect 4672 14368 4896 14396
rect 4672 14356 4678 14368
rect 4890 14356 4896 14368
rect 4948 14396 4954 14408
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 4948 14368 5089 14396
rect 4948 14356 4954 14368
rect 5077 14365 5089 14368
rect 5123 14365 5135 14399
rect 5077 14359 5135 14365
rect 5169 14399 5227 14405
rect 5169 14365 5181 14399
rect 5215 14396 5227 14399
rect 5258 14396 5264 14408
rect 5215 14368 5264 14396
rect 5215 14365 5227 14368
rect 5169 14359 5227 14365
rect 5258 14356 5264 14368
rect 5316 14356 5322 14408
rect 6454 14396 6460 14408
rect 6367 14368 6460 14396
rect 6454 14356 6460 14368
rect 6512 14356 6518 14408
rect 6549 14399 6607 14405
rect 6549 14365 6561 14399
rect 6595 14396 6607 14399
rect 6638 14396 6644 14408
rect 6595 14368 6644 14396
rect 6595 14365 6607 14368
rect 6549 14359 6607 14365
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 7098 14396 7104 14408
rect 7011 14368 7104 14396
rect 7098 14356 7104 14368
rect 7156 14396 7162 14408
rect 9674 14396 9680 14408
rect 7156 14368 9680 14396
rect 7156 14356 7162 14368
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 10134 14396 10140 14408
rect 10095 14368 10140 14396
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 10428 14405 10456 14436
rect 10962 14424 10968 14476
rect 11020 14464 11026 14476
rect 19886 14464 19892 14476
rect 11020 14436 14596 14464
rect 19847 14436 19892 14464
rect 11020 14424 11026 14436
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 2869 14331 2927 14337
rect 2869 14328 2881 14331
rect 2746 14300 2881 14328
rect 2869 14297 2881 14300
rect 2915 14328 2927 14331
rect 6472 14328 6500 14356
rect 8021 14331 8079 14337
rect 8021 14328 8033 14331
rect 2915 14300 8033 14328
rect 2915 14297 2927 14300
rect 2869 14291 2927 14297
rect 8021 14297 8033 14300
rect 8067 14297 8079 14331
rect 8021 14291 8079 14297
rect 9125 14331 9183 14337
rect 9125 14297 9137 14331
rect 9171 14297 9183 14331
rect 9306 14328 9312 14340
rect 9267 14300 9312 14328
rect 9125 14291 9183 14297
rect 1765 14263 1823 14269
rect 1765 14229 1777 14263
rect 1811 14260 1823 14263
rect 1854 14260 1860 14272
rect 1811 14232 1860 14260
rect 1811 14229 1823 14232
rect 1765 14223 1823 14229
rect 1854 14220 1860 14232
rect 1912 14220 1918 14272
rect 4157 14263 4215 14269
rect 4157 14229 4169 14263
rect 4203 14260 4215 14263
rect 4246 14260 4252 14272
rect 4203 14232 4252 14260
rect 4203 14229 4215 14232
rect 4157 14223 4215 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 6178 14260 6184 14272
rect 6139 14232 6184 14260
rect 6178 14220 6184 14232
rect 6236 14220 6242 14272
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 7834 14260 7840 14272
rect 7607 14232 7840 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 9140 14260 9168 14291
rect 9306 14288 9312 14300
rect 9364 14288 9370 14340
rect 10244 14328 10272 14359
rect 10502 14356 10508 14408
rect 10560 14396 10566 14408
rect 11330 14396 11336 14408
rect 10560 14368 10605 14396
rect 11291 14368 11336 14396
rect 10560 14356 10566 14368
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 11606 14396 11612 14408
rect 11567 14368 11612 14396
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 14274 14396 14280 14408
rect 14235 14368 14280 14396
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 14568 14405 14596 14436
rect 19886 14424 19892 14436
rect 19944 14424 19950 14476
rect 20622 14464 20628 14476
rect 20535 14436 20628 14464
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 20809 14467 20867 14473
rect 20809 14433 20821 14467
rect 20855 14464 20867 14467
rect 21726 14464 21732 14476
rect 20855 14436 21732 14464
rect 20855 14433 20867 14436
rect 20809 14427 20867 14433
rect 21726 14424 21732 14436
rect 21784 14424 21790 14476
rect 23676 14464 23704 14504
rect 27338 14492 27344 14504
rect 27396 14492 27402 14544
rect 22066 14436 23704 14464
rect 23753 14467 23811 14473
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14365 14611 14399
rect 15562 14396 15568 14408
rect 15523 14368 15568 14396
rect 14553 14359 14611 14365
rect 11974 14328 11980 14340
rect 10244 14300 11980 14328
rect 11974 14288 11980 14300
rect 12032 14328 12038 14340
rect 12069 14331 12127 14337
rect 12069 14328 12081 14331
rect 12032 14300 12081 14328
rect 12032 14288 12038 14300
rect 12069 14297 12081 14300
rect 12115 14297 12127 14331
rect 14476 14328 14504 14359
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14365 15991 14399
rect 15933 14359 15991 14365
rect 14642 14328 14648 14340
rect 14476 14300 14648 14328
rect 12069 14291 12127 14297
rect 14642 14288 14648 14300
rect 14700 14288 14706 14340
rect 15470 14288 15476 14340
rect 15528 14328 15534 14340
rect 15948 14328 15976 14359
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 17865 14399 17923 14405
rect 17865 14396 17877 14399
rect 17092 14368 17877 14396
rect 17092 14356 17098 14368
rect 17865 14365 17877 14368
rect 17911 14365 17923 14399
rect 17865 14359 17923 14365
rect 18233 14399 18291 14405
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 18279 14368 19625 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 19613 14365 19625 14368
rect 19659 14396 19671 14399
rect 20898 14396 20904 14408
rect 19659 14368 20576 14396
rect 20859 14368 20904 14396
rect 19659 14365 19671 14368
rect 19613 14359 19671 14365
rect 15528 14300 15976 14328
rect 15528 14288 15534 14300
rect 17310 14288 17316 14340
rect 17368 14328 17374 14340
rect 17405 14331 17463 14337
rect 17405 14328 17417 14331
rect 17368 14300 17417 14328
rect 17368 14288 17374 14300
rect 17405 14297 17417 14300
rect 17451 14297 17463 14331
rect 17880 14328 17908 14359
rect 20441 14331 20499 14337
rect 20441 14328 20453 14331
rect 17880 14300 20453 14328
rect 17405 14291 17463 14297
rect 20441 14297 20453 14300
rect 20487 14297 20499 14331
rect 20548 14328 20576 14368
rect 20898 14356 20904 14368
rect 20956 14396 20962 14408
rect 22066 14396 22094 14436
rect 23753 14433 23765 14467
rect 23799 14464 23811 14467
rect 24397 14467 24455 14473
rect 24397 14464 24409 14467
rect 23799 14436 24409 14464
rect 23799 14433 23811 14436
rect 23753 14427 23811 14433
rect 24397 14433 24409 14436
rect 24443 14464 24455 14467
rect 24762 14464 24768 14476
rect 24443 14436 24768 14464
rect 24443 14433 24455 14436
rect 24397 14427 24455 14433
rect 24762 14424 24768 14436
rect 24820 14424 24826 14476
rect 25038 14464 25044 14476
rect 24999 14436 25044 14464
rect 25038 14424 25044 14436
rect 25096 14424 25102 14476
rect 20956 14368 22094 14396
rect 23661 14399 23719 14405
rect 20956 14356 20962 14368
rect 23661 14365 23673 14399
rect 23707 14365 23719 14399
rect 23661 14359 23719 14365
rect 23845 14399 23903 14405
rect 23845 14365 23857 14399
rect 23891 14396 23903 14399
rect 23934 14396 23940 14408
rect 23891 14368 23940 14396
rect 23891 14365 23903 14368
rect 23845 14359 23903 14365
rect 20806 14328 20812 14340
rect 20548 14300 20812 14328
rect 20441 14291 20499 14297
rect 20806 14288 20812 14300
rect 20864 14288 20870 14340
rect 21082 14288 21088 14340
rect 21140 14328 21146 14340
rect 21513 14331 21571 14337
rect 21513 14328 21525 14331
rect 21140 14300 21525 14328
rect 21140 14288 21146 14300
rect 21513 14297 21525 14300
rect 21559 14297 21571 14331
rect 21726 14328 21732 14340
rect 21687 14300 21732 14328
rect 21513 14291 21571 14297
rect 21726 14288 21732 14300
rect 21784 14328 21790 14340
rect 23676 14328 23704 14359
rect 23934 14356 23940 14368
rect 23992 14356 23998 14408
rect 24578 14405 24584 14408
rect 24555 14399 24584 14405
rect 24555 14365 24567 14399
rect 24555 14359 24584 14365
rect 24578 14356 24584 14359
rect 24636 14356 24642 14408
rect 24854 14396 24860 14408
rect 24815 14368 24860 14396
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 27816 14405 27844 14560
rect 27890 14424 27896 14476
rect 27948 14464 27954 14476
rect 27985 14467 28043 14473
rect 27985 14464 27997 14467
rect 27948 14436 27997 14464
rect 27948 14424 27954 14436
rect 27985 14433 27997 14436
rect 28031 14464 28043 14467
rect 28629 14467 28687 14473
rect 28629 14464 28641 14467
rect 28031 14436 28641 14464
rect 28031 14433 28043 14436
rect 27985 14427 28043 14433
rect 28629 14433 28641 14436
rect 28675 14433 28687 14467
rect 28629 14427 28687 14433
rect 27801 14399 27859 14405
rect 27801 14365 27813 14399
rect 27847 14365 27859 14399
rect 27801 14359 27859 14365
rect 24302 14328 24308 14340
rect 21784 14300 22094 14328
rect 23676 14300 24308 14328
rect 21784 14288 21790 14300
rect 9582 14260 9588 14272
rect 9140 14232 9588 14260
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 10928 14232 11161 14260
rect 10928 14220 10934 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11149 14223 11207 14229
rect 11517 14263 11575 14269
rect 11517 14229 11529 14263
rect 11563 14260 11575 14263
rect 11606 14260 11612 14272
rect 11563 14232 11612 14260
rect 11563 14229 11575 14232
rect 11517 14223 11575 14229
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 12618 14220 12624 14272
rect 12676 14260 12682 14272
rect 20070 14260 20076 14272
rect 12676 14232 20076 14260
rect 12676 14220 12682 14232
rect 20070 14220 20076 14232
rect 20128 14220 20134 14272
rect 21174 14220 21180 14272
rect 21232 14260 21238 14272
rect 21361 14263 21419 14269
rect 21361 14260 21373 14263
rect 21232 14232 21373 14260
rect 21232 14220 21238 14232
rect 21361 14229 21373 14232
rect 21407 14229 21419 14263
rect 22066 14260 22094 14300
rect 24302 14288 24308 14300
rect 24360 14328 24366 14340
rect 24673 14331 24731 14337
rect 24673 14328 24685 14331
rect 24360 14300 24685 14328
rect 24360 14288 24366 14300
rect 24673 14297 24685 14300
rect 24719 14297 24731 14331
rect 24673 14291 24731 14297
rect 24765 14331 24823 14337
rect 24765 14297 24777 14331
rect 24811 14328 24823 14331
rect 25590 14328 25596 14340
rect 24811 14300 25596 14328
rect 24811 14297 24823 14300
rect 24765 14291 24823 14297
rect 25590 14288 25596 14300
rect 25648 14288 25654 14340
rect 26326 14288 26332 14340
rect 26384 14328 26390 14340
rect 26421 14331 26479 14337
rect 26421 14328 26433 14331
rect 26384 14300 26433 14328
rect 26384 14288 26390 14300
rect 26421 14297 26433 14300
rect 26467 14328 26479 14331
rect 27893 14331 27951 14337
rect 27893 14328 27905 14331
rect 26467 14300 27905 14328
rect 26467 14297 26479 14300
rect 26421 14291 26479 14297
rect 27893 14297 27905 14300
rect 27939 14297 27951 14331
rect 27893 14291 27951 14297
rect 22554 14260 22560 14272
rect 22066 14232 22560 14260
rect 21361 14223 21419 14229
rect 22554 14220 22560 14232
rect 22612 14260 22618 14272
rect 25314 14260 25320 14272
rect 22612 14232 25320 14260
rect 22612 14220 22618 14232
rect 25314 14220 25320 14232
rect 25372 14220 25378 14272
rect 27433 14263 27491 14269
rect 27433 14229 27445 14263
rect 27479 14260 27491 14263
rect 27614 14260 27620 14272
rect 27479 14232 27620 14260
rect 27479 14229 27491 14232
rect 27433 14223 27491 14229
rect 27614 14220 27620 14232
rect 27672 14220 27678 14272
rect 1104 14170 29600 14192
rect 1104 14118 8034 14170
rect 8086 14118 8098 14170
rect 8150 14118 8162 14170
rect 8214 14118 8226 14170
rect 8278 14118 8290 14170
rect 8342 14118 15118 14170
rect 15170 14118 15182 14170
rect 15234 14118 15246 14170
rect 15298 14118 15310 14170
rect 15362 14118 15374 14170
rect 15426 14118 22202 14170
rect 22254 14118 22266 14170
rect 22318 14118 22330 14170
rect 22382 14118 22394 14170
rect 22446 14118 22458 14170
rect 22510 14118 29286 14170
rect 29338 14118 29350 14170
rect 29402 14118 29414 14170
rect 29466 14118 29478 14170
rect 29530 14118 29542 14170
rect 29594 14118 29600 14170
rect 1104 14096 29600 14118
rect 4249 14059 4307 14065
rect 4249 14025 4261 14059
rect 4295 14056 4307 14059
rect 4614 14056 4620 14068
rect 4295 14028 4620 14056
rect 4295 14025 4307 14028
rect 4249 14019 4307 14025
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 4893 14059 4951 14065
rect 4893 14025 4905 14059
rect 4939 14056 4951 14059
rect 5258 14056 5264 14068
rect 4939 14028 5264 14056
rect 4939 14025 4951 14028
rect 4893 14019 4951 14025
rect 4522 13948 4528 14000
rect 4580 13988 4586 14000
rect 4908 13988 4936 14019
rect 5258 14016 5264 14028
rect 5316 14056 5322 14068
rect 5445 14059 5503 14065
rect 5445 14056 5457 14059
rect 5316 14028 5457 14056
rect 5316 14016 5322 14028
rect 5445 14025 5457 14028
rect 5491 14025 5503 14059
rect 5445 14019 5503 14025
rect 8849 14059 8907 14065
rect 8849 14025 8861 14059
rect 8895 14056 8907 14059
rect 9674 14056 9680 14068
rect 8895 14028 9680 14056
rect 8895 14025 8907 14028
rect 8849 14019 8907 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 10594 14056 10600 14068
rect 10555 14028 10600 14056
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 15378 14056 15384 14068
rect 11572 14028 15384 14056
rect 11572 14016 11578 14028
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 15562 14056 15568 14068
rect 15523 14028 15568 14056
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 20622 14056 20628 14068
rect 19843 14028 20628 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 20622 14016 20628 14028
rect 20680 14016 20686 14068
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 21082 14056 21088 14068
rect 20864 14028 21088 14056
rect 20864 14016 20870 14028
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 23566 14056 23572 14068
rect 22066 14028 23572 14056
rect 6914 13988 6920 14000
rect 4580 13960 4936 13988
rect 6827 13960 6920 13988
rect 4580 13948 4586 13960
rect 6914 13948 6920 13960
rect 6972 13988 6978 14000
rect 7558 13988 7564 14000
rect 6972 13960 7564 13988
rect 6972 13948 6978 13960
rect 7558 13948 7564 13960
rect 7616 13948 7622 14000
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 12621 13991 12679 13997
rect 12621 13988 12633 13991
rect 10192 13960 12633 13988
rect 10192 13948 10198 13960
rect 12621 13957 12633 13960
rect 12667 13957 12679 13991
rect 12621 13951 12679 13957
rect 13998 13948 14004 14000
rect 14056 13988 14062 14000
rect 22066 13988 22094 14028
rect 23566 14016 23572 14028
rect 23624 14016 23630 14068
rect 24302 14016 24308 14068
rect 24360 14056 24366 14068
rect 24360 14028 24624 14056
rect 24360 14016 24366 14028
rect 24026 13988 24032 14000
rect 14056 13960 22094 13988
rect 22940 13960 24032 13988
rect 14056 13948 14062 13960
rect 1946 13920 1952 13932
rect 1907 13892 1952 13920
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13920 3755 13923
rect 4157 13923 4215 13929
rect 4157 13920 4169 13923
rect 3743 13892 4169 13920
rect 3743 13889 3755 13892
rect 3697 13883 3755 13889
rect 4157 13889 4169 13892
rect 4203 13920 4215 13923
rect 5810 13920 5816 13932
rect 4203 13892 5816 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 5810 13880 5816 13892
rect 5868 13880 5874 13932
rect 6822 13920 6828 13932
rect 6783 13892 6828 13920
rect 6822 13880 6828 13892
rect 6880 13880 6886 13932
rect 9030 13920 9036 13932
rect 8991 13892 9036 13920
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13920 9275 13923
rect 9490 13920 9496 13932
rect 9263 13892 9496 13920
rect 9263 13889 9275 13892
rect 9217 13883 9275 13889
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 9646 13892 10241 13920
rect 1854 13852 1860 13864
rect 1815 13824 1860 13852
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 9306 13852 9312 13864
rect 8444 13824 9312 13852
rect 8444 13812 8450 13824
rect 9306 13812 9312 13824
rect 9364 13852 9370 13864
rect 9646 13852 9674 13892
rect 10229 13889 10241 13892
rect 10275 13920 10287 13923
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 10275 13892 12081 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 12069 13889 12081 13892
rect 12115 13920 12127 13923
rect 12115 13892 12434 13920
rect 12115 13889 12127 13892
rect 12069 13883 12127 13889
rect 9364 13824 9674 13852
rect 9364 13812 9370 13824
rect 9766 13812 9772 13864
rect 9824 13852 9830 13864
rect 9950 13852 9956 13864
rect 9824 13824 9956 13852
rect 9824 13812 9830 13824
rect 9950 13812 9956 13824
rect 10008 13852 10014 13864
rect 10134 13852 10140 13864
rect 10008 13824 10140 13852
rect 10008 13812 10014 13824
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13821 10379 13855
rect 10321 13815 10379 13821
rect 9582 13744 9588 13796
rect 9640 13784 9646 13796
rect 10336 13784 10364 13815
rect 10410 13812 10416 13864
rect 10468 13852 10474 13864
rect 12406 13852 12434 13892
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 15473 13923 15531 13929
rect 15473 13920 15485 13923
rect 14332 13892 15485 13920
rect 14332 13880 14338 13892
rect 15473 13889 15485 13892
rect 15519 13889 15531 13923
rect 15473 13883 15531 13889
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 15838 13920 15844 13932
rect 15703 13892 15844 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 19705 13923 19763 13929
rect 19705 13920 19717 13923
rect 19352 13892 19717 13920
rect 19352 13864 19380 13892
rect 19705 13889 19717 13892
rect 19751 13889 19763 13923
rect 19705 13883 19763 13889
rect 19886 13880 19892 13932
rect 19944 13920 19950 13932
rect 20438 13920 20444 13932
rect 19944 13892 20444 13920
rect 19944 13880 19950 13892
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 20717 13923 20775 13929
rect 20717 13920 20729 13923
rect 20548 13892 20729 13920
rect 12618 13852 12624 13864
rect 10468 13824 10513 13852
rect 12406 13824 12624 13852
rect 10468 13812 10474 13824
rect 12618 13812 12624 13824
rect 12676 13812 12682 13864
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 19153 13855 19211 13861
rect 19153 13852 19165 13855
rect 12860 13824 19165 13852
rect 12860 13812 12866 13824
rect 19153 13821 19165 13824
rect 19199 13852 19211 13855
rect 19334 13852 19340 13864
rect 19199 13824 19340 13852
rect 19199 13821 19211 13824
rect 19153 13815 19211 13821
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 20548 13852 20576 13892
rect 20717 13889 20729 13892
rect 20763 13920 20775 13923
rect 21266 13920 21272 13932
rect 20763 13892 21272 13920
rect 20763 13889 20775 13892
rect 20717 13883 20775 13889
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 22940 13929 22968 13960
rect 24026 13948 24032 13960
rect 24084 13948 24090 14000
rect 24486 13988 24492 14000
rect 24447 13960 24492 13988
rect 24486 13948 24492 13960
rect 24544 13948 24550 14000
rect 24596 13997 24624 14028
rect 24762 14016 24768 14068
rect 24820 14056 24826 14068
rect 28626 14056 28632 14068
rect 24820 14028 24900 14056
rect 28587 14028 28632 14056
rect 24820 14016 24826 14028
rect 24581 13991 24639 13997
rect 24581 13957 24593 13991
rect 24627 13957 24639 13991
rect 24581 13951 24639 13957
rect 22925 13923 22983 13929
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 22925 13883 22983 13889
rect 23109 13923 23167 13929
rect 23109 13889 23121 13923
rect 23155 13889 23167 13923
rect 23109 13883 23167 13889
rect 24397 13923 24455 13929
rect 24397 13889 24409 13923
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 20806 13852 20812 13864
rect 20312 13824 20576 13852
rect 20767 13824 20812 13852
rect 20312 13812 20318 13824
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 11514 13784 11520 13796
rect 9640 13756 11520 13784
rect 9640 13744 9646 13756
rect 11514 13744 11520 13756
rect 11572 13744 11578 13796
rect 21266 13744 21272 13796
rect 21324 13784 21330 13796
rect 21818 13784 21824 13796
rect 21324 13756 21824 13784
rect 21324 13744 21330 13756
rect 21818 13744 21824 13756
rect 21876 13744 21882 13796
rect 23124 13784 23152 13883
rect 24412 13852 24440 13883
rect 24670 13880 24676 13932
rect 24728 13929 24734 13932
rect 24872 13929 24900 14028
rect 28626 14016 28632 14028
rect 28684 14016 28690 14068
rect 27430 13988 27436 14000
rect 27391 13960 27436 13988
rect 27430 13948 27436 13960
rect 27488 13948 27494 14000
rect 24728 13923 24757 13929
rect 24745 13889 24757 13923
rect 24728 13883 24757 13889
rect 24857 13923 24915 13929
rect 24857 13889 24869 13923
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 24728 13880 24734 13883
rect 27338 13880 27344 13932
rect 27396 13920 27402 13932
rect 27709 13923 27767 13929
rect 27709 13920 27721 13923
rect 27396 13892 27721 13920
rect 27396 13880 27402 13892
rect 27709 13889 27721 13892
rect 27755 13920 27767 13923
rect 28258 13920 28264 13932
rect 27755 13892 28264 13920
rect 27755 13889 27767 13892
rect 27709 13883 27767 13889
rect 28258 13880 28264 13892
rect 28316 13880 28322 13932
rect 28442 13920 28448 13932
rect 28403 13892 28448 13920
rect 28442 13880 28448 13892
rect 28500 13880 28506 13932
rect 26510 13852 26516 13864
rect 24412 13824 26516 13852
rect 26510 13812 26516 13824
rect 26568 13812 26574 13864
rect 27433 13855 27491 13861
rect 27433 13821 27445 13855
rect 27479 13852 27491 13855
rect 28074 13852 28080 13864
rect 27479 13824 28080 13852
rect 27479 13821 27491 13824
rect 27433 13815 27491 13821
rect 28074 13812 28080 13824
rect 28132 13812 28138 13864
rect 24578 13784 24584 13796
rect 23124 13756 24584 13784
rect 24578 13744 24584 13756
rect 24636 13744 24642 13796
rect 27614 13784 27620 13796
rect 27575 13756 27620 13784
rect 27614 13744 27620 13756
rect 27672 13744 27678 13796
rect 2130 13676 2136 13728
rect 2188 13716 2194 13728
rect 2225 13719 2283 13725
rect 2225 13716 2237 13719
rect 2188 13688 2237 13716
rect 2188 13676 2194 13688
rect 2225 13685 2237 13688
rect 2271 13685 2283 13719
rect 2225 13679 2283 13685
rect 10594 13676 10600 13728
rect 10652 13716 10658 13728
rect 11606 13716 11612 13728
rect 10652 13688 11612 13716
rect 10652 13676 10658 13688
rect 11606 13676 11612 13688
rect 11664 13716 11670 13728
rect 14734 13716 14740 13728
rect 11664 13688 14740 13716
rect 11664 13676 11670 13688
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 20438 13716 20444 13728
rect 20399 13688 20444 13716
rect 20438 13676 20444 13688
rect 20496 13676 20502 13728
rect 23014 13716 23020 13728
rect 22975 13688 23020 13716
rect 23014 13676 23020 13688
rect 23072 13676 23078 13728
rect 24210 13716 24216 13728
rect 24171 13688 24216 13716
rect 24210 13676 24216 13688
rect 24268 13676 24274 13728
rect 1104 13626 29440 13648
rect 1104 13574 4492 13626
rect 4544 13574 4556 13626
rect 4608 13574 4620 13626
rect 4672 13574 4684 13626
rect 4736 13574 4748 13626
rect 4800 13574 11576 13626
rect 11628 13574 11640 13626
rect 11692 13574 11704 13626
rect 11756 13574 11768 13626
rect 11820 13574 11832 13626
rect 11884 13574 18660 13626
rect 18712 13574 18724 13626
rect 18776 13574 18788 13626
rect 18840 13574 18852 13626
rect 18904 13574 18916 13626
rect 18968 13574 25744 13626
rect 25796 13574 25808 13626
rect 25860 13574 25872 13626
rect 25924 13574 25936 13626
rect 25988 13574 26000 13626
rect 26052 13574 29440 13626
rect 1104 13552 29440 13574
rect 10321 13515 10379 13521
rect 10321 13481 10333 13515
rect 10367 13512 10379 13515
rect 10410 13512 10416 13524
rect 10367 13484 10416 13512
rect 10367 13481 10379 13484
rect 10321 13475 10379 13481
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 10502 13472 10508 13524
rect 10560 13512 10566 13524
rect 10781 13515 10839 13521
rect 10781 13512 10793 13515
rect 10560 13484 10793 13512
rect 10560 13472 10566 13484
rect 10781 13481 10793 13484
rect 10827 13512 10839 13515
rect 10962 13512 10968 13524
rect 10827 13484 10968 13512
rect 10827 13481 10839 13484
rect 10781 13475 10839 13481
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 14366 13472 14372 13524
rect 14424 13512 14430 13524
rect 24210 13512 24216 13524
rect 14424 13484 24216 13512
rect 14424 13472 14430 13484
rect 24210 13472 24216 13484
rect 24268 13472 24274 13524
rect 25590 13472 25596 13524
rect 25648 13512 25654 13524
rect 25685 13515 25743 13521
rect 25685 13512 25697 13515
rect 25648 13484 25697 13512
rect 25648 13472 25654 13484
rect 25685 13481 25697 13484
rect 25731 13481 25743 13515
rect 26510 13512 26516 13524
rect 26471 13484 26516 13512
rect 25685 13475 25743 13481
rect 26510 13472 26516 13484
rect 26568 13472 26574 13524
rect 28353 13515 28411 13521
rect 28353 13481 28365 13515
rect 28399 13512 28411 13515
rect 28442 13512 28448 13524
rect 28399 13484 28448 13512
rect 28399 13481 28411 13484
rect 28353 13475 28411 13481
rect 28442 13472 28448 13484
rect 28500 13472 28506 13524
rect 12802 13404 12808 13456
rect 12860 13444 12866 13456
rect 13170 13444 13176 13456
rect 12860 13416 13176 13444
rect 12860 13404 12866 13416
rect 13170 13404 13176 13416
rect 13228 13404 13234 13456
rect 19334 13444 19340 13456
rect 19295 13416 19340 13444
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 20254 13444 20260 13456
rect 20215 13416 20260 13444
rect 20254 13404 20260 13416
rect 20312 13404 20318 13456
rect 22738 13444 22744 13456
rect 22699 13416 22744 13444
rect 22738 13404 22744 13416
rect 22796 13404 22802 13456
rect 23934 13404 23940 13456
rect 23992 13444 23998 13456
rect 24762 13444 24768 13456
rect 23992 13416 24768 13444
rect 23992 13404 23998 13416
rect 24762 13404 24768 13416
rect 24820 13444 24826 13456
rect 25041 13447 25099 13453
rect 25041 13444 25053 13447
rect 24820 13416 25053 13444
rect 24820 13404 24826 13416
rect 25041 13413 25053 13416
rect 25087 13413 25099 13447
rect 25041 13407 25099 13413
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 8570 13376 8576 13388
rect 7064 13348 8576 13376
rect 7064 13336 7070 13348
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 1719 13280 2268 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 2240 13181 2268 13280
rect 7466 13268 7472 13320
rect 7524 13308 7530 13320
rect 7944 13317 7972 13348
rect 8570 13336 8576 13348
rect 8628 13376 8634 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8628 13348 8953 13376
rect 8628 13336 8634 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 20438 13336 20444 13388
rect 20496 13376 20502 13388
rect 21453 13379 21511 13385
rect 21453 13376 21465 13379
rect 20496 13348 21465 13376
rect 20496 13336 20502 13348
rect 21453 13345 21465 13348
rect 21499 13345 21511 13379
rect 21453 13339 21511 13345
rect 25608 13348 26464 13376
rect 7745 13311 7803 13317
rect 7745 13308 7757 13311
rect 7524 13280 7757 13308
rect 7524 13268 7530 13280
rect 7745 13277 7757 13280
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13308 8355 13311
rect 10318 13308 10324 13320
rect 8343 13280 10324 13308
rect 8343 13277 8355 13280
rect 8297 13271 8355 13277
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 12621 13311 12679 13317
rect 12621 13277 12633 13311
rect 12667 13308 12679 13311
rect 12710 13308 12716 13320
rect 12667 13280 12716 13308
rect 12667 13277 12679 13280
rect 12621 13271 12679 13277
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 13354 13308 13360 13320
rect 12851 13280 13360 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 18138 13308 18144 13320
rect 13504 13280 18144 13308
rect 13504 13268 13510 13280
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 21174 13308 21180 13320
rect 21135 13280 21180 13308
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 21358 13308 21364 13320
rect 21319 13280 21364 13308
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 22554 13268 22560 13320
rect 22612 13308 22618 13320
rect 22925 13311 22983 13317
rect 22925 13308 22937 13311
rect 22612 13280 22937 13308
rect 22612 13268 22618 13280
rect 22925 13277 22937 13280
rect 22971 13277 22983 13311
rect 22925 13271 22983 13277
rect 23014 13268 23020 13320
rect 23072 13308 23078 13320
rect 23109 13311 23167 13317
rect 23109 13308 23121 13311
rect 23072 13280 23121 13308
rect 23072 13268 23078 13280
rect 23109 13277 23121 13280
rect 23155 13277 23167 13311
rect 24302 13308 24308 13320
rect 23109 13271 23167 13277
rect 23492 13280 24308 13308
rect 8662 13200 8668 13252
rect 8720 13240 8726 13252
rect 9582 13240 9588 13252
rect 8720 13212 9588 13240
rect 8720 13200 8726 13212
rect 9582 13200 9588 13212
rect 9640 13240 9646 13252
rect 9677 13243 9735 13249
rect 9677 13240 9689 13243
rect 9640 13212 9689 13240
rect 9640 13200 9646 13212
rect 9677 13209 9689 13212
rect 9723 13240 9735 13243
rect 11333 13243 11391 13249
rect 11333 13240 11345 13243
rect 9723 13212 11345 13240
rect 9723 13209 9735 13212
rect 9677 13203 9735 13209
rect 11333 13209 11345 13212
rect 11379 13209 11391 13243
rect 13464 13240 13492 13268
rect 23492 13252 23520 13280
rect 24302 13268 24308 13280
rect 24360 13308 24366 13320
rect 24397 13311 24455 13317
rect 24397 13308 24409 13311
rect 24360 13280 24409 13308
rect 24360 13268 24366 13280
rect 24397 13277 24409 13280
rect 24443 13277 24455 13311
rect 24397 13271 24455 13277
rect 25498 13268 25504 13320
rect 25556 13308 25562 13320
rect 25608 13317 25636 13348
rect 25593 13311 25651 13317
rect 25593 13308 25605 13311
rect 25556 13280 25605 13308
rect 25556 13268 25562 13280
rect 25593 13277 25605 13280
rect 25639 13277 25651 13311
rect 25593 13271 25651 13277
rect 25777 13311 25835 13317
rect 25777 13277 25789 13311
rect 25823 13308 25835 13311
rect 26234 13308 26240 13320
rect 25823 13280 26240 13308
rect 25823 13277 25835 13280
rect 25777 13271 25835 13277
rect 26234 13268 26240 13280
rect 26292 13268 26298 13320
rect 26436 13317 26464 13348
rect 26421 13311 26479 13317
rect 26421 13277 26433 13311
rect 26467 13277 26479 13311
rect 26602 13308 26608 13320
rect 26563 13280 26608 13308
rect 26421 13271 26479 13277
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 11333 13203 11391 13209
rect 12406 13212 13492 13240
rect 2225 13175 2283 13181
rect 2225 13141 2237 13175
rect 2271 13172 2283 13175
rect 2682 13172 2688 13184
rect 2271 13144 2688 13172
rect 2271 13141 2283 13144
rect 2225 13135 2283 13141
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 7929 13175 7987 13181
rect 7929 13172 7941 13175
rect 6880 13144 7941 13172
rect 6880 13132 6886 13144
rect 7929 13141 7941 13144
rect 7975 13141 7987 13175
rect 7929 13135 7987 13141
rect 8478 13132 8484 13184
rect 8536 13172 8542 13184
rect 12406 13172 12434 13212
rect 17310 13200 17316 13252
rect 17368 13240 17374 13252
rect 23474 13240 23480 13252
rect 17368 13212 23480 13240
rect 17368 13200 17374 13212
rect 23474 13200 23480 13212
rect 23532 13200 23538 13252
rect 8536 13144 12434 13172
rect 8536 13132 8542 13144
rect 12618 13132 12624 13184
rect 12676 13172 12682 13184
rect 12713 13175 12771 13181
rect 12713 13172 12725 13175
rect 12676 13144 12725 13172
rect 12676 13132 12682 13144
rect 12713 13141 12725 13144
rect 12759 13141 12771 13175
rect 15838 13172 15844 13184
rect 15799 13144 15844 13172
rect 12713 13135 12771 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 20530 13132 20536 13184
rect 20588 13172 20594 13184
rect 20993 13175 21051 13181
rect 20993 13172 21005 13175
rect 20588 13144 21005 13172
rect 20588 13132 20594 13144
rect 20993 13141 21005 13144
rect 21039 13141 21051 13175
rect 20993 13135 21051 13141
rect 23014 13132 23020 13184
rect 23072 13172 23078 13184
rect 23072 13144 23117 13172
rect 23072 13132 23078 13144
rect 23198 13132 23204 13184
rect 23256 13172 23262 13184
rect 23293 13175 23351 13181
rect 23293 13172 23305 13175
rect 23256 13144 23305 13172
rect 23256 13132 23262 13144
rect 23293 13141 23305 13144
rect 23339 13141 23351 13175
rect 23293 13135 23351 13141
rect 24489 13175 24547 13181
rect 24489 13141 24501 13175
rect 24535 13172 24547 13175
rect 24578 13172 24584 13184
rect 24535 13144 24584 13172
rect 24535 13141 24547 13144
rect 24489 13135 24547 13141
rect 24578 13132 24584 13144
rect 24636 13132 24642 13184
rect 27801 13175 27859 13181
rect 27801 13141 27813 13175
rect 27847 13172 27859 13175
rect 28166 13172 28172 13184
rect 27847 13144 28172 13172
rect 27847 13141 27859 13144
rect 27801 13135 27859 13141
rect 28166 13132 28172 13144
rect 28224 13132 28230 13184
rect 1104 13082 29600 13104
rect 1104 13030 8034 13082
rect 8086 13030 8098 13082
rect 8150 13030 8162 13082
rect 8214 13030 8226 13082
rect 8278 13030 8290 13082
rect 8342 13030 15118 13082
rect 15170 13030 15182 13082
rect 15234 13030 15246 13082
rect 15298 13030 15310 13082
rect 15362 13030 15374 13082
rect 15426 13030 22202 13082
rect 22254 13030 22266 13082
rect 22318 13030 22330 13082
rect 22382 13030 22394 13082
rect 22446 13030 22458 13082
rect 22510 13030 29286 13082
rect 29338 13030 29350 13082
rect 29402 13030 29414 13082
rect 29466 13030 29478 13082
rect 29530 13030 29542 13082
rect 29594 13030 29600 13082
rect 1104 13008 29600 13030
rect 7466 12968 7472 12980
rect 7427 12940 7472 12968
rect 7466 12928 7472 12940
rect 7524 12928 7530 12980
rect 10318 12968 10324 12980
rect 7576 12940 9168 12968
rect 10279 12940 10324 12968
rect 5994 12860 6000 12912
rect 6052 12900 6058 12912
rect 7576 12900 7604 12940
rect 8386 12900 8392 12912
rect 6052 12872 7604 12900
rect 8299 12872 8392 12900
rect 6052 12860 6058 12872
rect 8386 12860 8392 12872
rect 8444 12900 8450 12912
rect 8444 12872 9076 12900
rect 8444 12860 8450 12872
rect 9048 12844 9076 12872
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 5859 12804 6377 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6365 12801 6377 12804
rect 6411 12832 6423 12835
rect 6914 12832 6920 12844
rect 6411 12804 6920 12832
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7101 12835 7159 12841
rect 7101 12832 7113 12835
rect 7024 12804 7113 12832
rect 7024 12708 7052 12804
rect 7101 12801 7113 12804
rect 7147 12801 7159 12835
rect 7101 12795 7159 12801
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 8021 12835 8079 12841
rect 8021 12832 8033 12835
rect 7340 12804 8033 12832
rect 7340 12792 7346 12804
rect 8021 12801 8033 12804
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12832 8355 12835
rect 8478 12832 8484 12844
rect 8343 12804 8484 12832
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12733 7251 12767
rect 8036 12764 8064 12795
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 9030 12832 9036 12844
rect 8904 12804 8949 12832
rect 8991 12804 9036 12832
rect 8904 12792 8910 12804
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 8662 12764 8668 12776
rect 8036 12736 8668 12764
rect 7193 12727 7251 12733
rect 7006 12656 7012 12708
rect 7064 12656 7070 12708
rect 5721 12631 5779 12637
rect 5721 12597 5733 12631
rect 5767 12628 5779 12631
rect 5902 12628 5908 12640
rect 5767 12600 5908 12628
rect 5767 12597 5779 12600
rect 5721 12591 5779 12597
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 7208 12628 7236 12727
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 9140 12764 9168 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 14366 12968 14372 12980
rect 10520 12940 14372 12968
rect 10520 12863 10548 12940
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 14458 12928 14464 12980
rect 14516 12968 14522 12980
rect 14642 12968 14648 12980
rect 14516 12940 14648 12968
rect 14516 12928 14522 12940
rect 14642 12928 14648 12940
rect 14700 12928 14706 12980
rect 14734 12928 14740 12980
rect 14792 12968 14798 12980
rect 17034 12968 17040 12980
rect 14792 12940 17040 12968
rect 14792 12928 14798 12940
rect 17034 12928 17040 12940
rect 17092 12928 17098 12980
rect 17497 12971 17555 12977
rect 17497 12937 17509 12971
rect 17543 12968 17555 12971
rect 19058 12968 19064 12980
rect 17543 12940 19064 12968
rect 17543 12937 17555 12940
rect 17497 12931 17555 12937
rect 11974 12900 11980 12912
rect 10796 12872 11836 12900
rect 11935 12872 11980 12900
rect 10497 12857 10555 12863
rect 10497 12823 10509 12857
rect 10543 12823 10555 12857
rect 10497 12817 10555 12823
rect 10594 12792 10600 12844
rect 10652 12832 10658 12844
rect 10796 12841 10824 12872
rect 10781 12835 10839 12841
rect 10652 12804 10697 12832
rect 10652 12792 10658 12804
rect 10781 12801 10793 12835
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12801 10931 12835
rect 11808 12832 11836 12872
rect 11974 12860 11980 12872
rect 12032 12860 12038 12912
rect 14568 12872 16712 12900
rect 12066 12832 12072 12844
rect 11808 12804 12072 12832
rect 10873 12795 10931 12801
rect 9140 12736 9674 12764
rect 7834 12656 7840 12708
rect 7892 12696 7898 12708
rect 8846 12696 8852 12708
rect 7892 12668 8852 12696
rect 7892 12656 7898 12668
rect 8846 12656 8852 12668
rect 8904 12656 8910 12708
rect 9646 12696 9674 12736
rect 10888 12696 10916 12795
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 13446 12832 13452 12844
rect 13035 12804 13452 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 14568 12841 14596 12872
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12832 13691 12835
rect 14553 12835 14611 12841
rect 14553 12832 14565 12835
rect 13679 12804 14565 12832
rect 13679 12801 13691 12804
rect 13633 12795 13691 12801
rect 14553 12801 14565 12804
rect 14599 12801 14611 12835
rect 14734 12832 14740 12844
rect 14695 12804 14740 12832
rect 14553 12795 14611 12801
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 16482 12832 16488 12844
rect 15335 12804 16488 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 12802 12724 12808 12776
rect 12860 12764 12866 12776
rect 15378 12764 15384 12776
rect 12860 12736 15384 12764
rect 12860 12724 12866 12736
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 16684 12773 16712 12872
rect 16945 12835 17003 12841
rect 16945 12801 16957 12835
rect 16991 12832 17003 12835
rect 17512 12832 17540 12931
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 20165 12971 20223 12977
rect 20165 12937 20177 12971
rect 20211 12968 20223 12971
rect 20254 12968 20260 12980
rect 20211 12940 20260 12968
rect 20211 12937 20223 12940
rect 20165 12931 20223 12937
rect 18049 12903 18107 12909
rect 18049 12869 18061 12903
rect 18095 12900 18107 12903
rect 18322 12900 18328 12912
rect 18095 12872 18328 12900
rect 18095 12869 18107 12872
rect 18049 12863 18107 12869
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 20180 12900 20208 12931
rect 20254 12928 20260 12940
rect 20312 12928 20318 12980
rect 20717 12971 20775 12977
rect 20717 12937 20729 12971
rect 20763 12968 20775 12971
rect 20806 12968 20812 12980
rect 20763 12940 20812 12968
rect 20763 12937 20775 12940
rect 20717 12931 20775 12937
rect 20806 12928 20812 12940
rect 20864 12928 20870 12980
rect 23014 12928 23020 12980
rect 23072 12968 23078 12980
rect 23937 12971 23995 12977
rect 23937 12968 23949 12971
rect 23072 12940 23949 12968
rect 23072 12928 23078 12940
rect 23937 12937 23949 12940
rect 23983 12937 23995 12971
rect 23937 12931 23995 12937
rect 24762 12928 24768 12980
rect 24820 12968 24826 12980
rect 25317 12971 25375 12977
rect 25317 12968 25329 12971
rect 24820 12940 25329 12968
rect 24820 12928 24826 12940
rect 25317 12937 25329 12940
rect 25363 12937 25375 12971
rect 25317 12931 25375 12937
rect 26602 12928 26608 12980
rect 26660 12968 26666 12980
rect 26878 12968 26884 12980
rect 26660 12940 26884 12968
rect 26660 12928 26666 12940
rect 26878 12928 26884 12940
rect 26936 12968 26942 12980
rect 27249 12971 27307 12977
rect 27249 12968 27261 12971
rect 26936 12940 27261 12968
rect 26936 12928 26942 12940
rect 27249 12937 27261 12940
rect 27295 12937 27307 12971
rect 27249 12931 27307 12937
rect 27617 12971 27675 12977
rect 27617 12937 27629 12971
rect 27663 12968 27675 12971
rect 27706 12968 27712 12980
rect 27663 12940 27712 12968
rect 27663 12937 27675 12940
rect 27617 12931 27675 12937
rect 27706 12928 27712 12940
rect 27764 12928 27770 12980
rect 20898 12900 20904 12912
rect 19352 12872 20208 12900
rect 20859 12872 20904 12900
rect 16991 12804 17540 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 19061 12835 19119 12841
rect 19061 12832 19073 12835
rect 18564 12804 19073 12832
rect 18564 12792 18570 12804
rect 19061 12801 19073 12804
rect 19107 12801 19119 12835
rect 19061 12795 19119 12801
rect 19153 12835 19211 12841
rect 19153 12801 19165 12835
rect 19199 12832 19211 12835
rect 19242 12832 19248 12844
rect 19199 12804 19248 12832
rect 19199 12801 19211 12804
rect 19153 12795 19211 12801
rect 19242 12792 19248 12804
rect 19300 12792 19306 12844
rect 19352 12841 19380 12872
rect 20898 12860 20904 12872
rect 20956 12900 20962 12912
rect 22738 12900 22744 12912
rect 20956 12872 22744 12900
rect 20956 12860 20962 12872
rect 22738 12860 22744 12872
rect 22796 12860 22802 12912
rect 23474 12900 23480 12912
rect 23216 12872 23480 12900
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12801 19395 12835
rect 19337 12795 19395 12801
rect 19429 12835 19487 12841
rect 19429 12801 19441 12835
rect 19475 12832 19487 12835
rect 21082 12832 21088 12844
rect 19475 12804 21088 12832
rect 19475 12801 19487 12804
rect 19429 12795 19487 12801
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 23216 12841 23244 12872
rect 23474 12860 23480 12872
rect 23532 12900 23538 12912
rect 23658 12900 23664 12912
rect 23532 12872 23664 12900
rect 23532 12860 23538 12872
rect 23658 12860 23664 12872
rect 23716 12900 23722 12912
rect 23716 12872 23980 12900
rect 23716 12860 23722 12872
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 23293 12835 23351 12841
rect 23293 12801 23305 12835
rect 23339 12832 23351 12835
rect 23566 12832 23572 12844
rect 23339 12804 23572 12832
rect 23339 12801 23351 12804
rect 23293 12795 23351 12801
rect 23566 12792 23572 12804
rect 23624 12792 23630 12844
rect 23952 12841 23980 12872
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12832 24179 12835
rect 24949 12835 25007 12841
rect 24949 12832 24961 12835
rect 24167 12804 24961 12832
rect 24167 12801 24179 12804
rect 24121 12795 24179 12801
rect 24949 12801 24961 12804
rect 24995 12801 25007 12835
rect 25130 12832 25136 12844
rect 25091 12804 25136 12832
rect 24949 12795 25007 12801
rect 25130 12792 25136 12804
rect 25188 12792 25194 12844
rect 25409 12835 25467 12841
rect 25409 12801 25421 12835
rect 25455 12832 25467 12835
rect 26234 12832 26240 12844
rect 25455 12804 26240 12832
rect 25455 12801 25467 12804
rect 25409 12795 25467 12801
rect 26234 12792 26240 12804
rect 26292 12832 26298 12844
rect 27246 12832 27252 12844
rect 26292 12804 27252 12832
rect 26292 12792 26298 12804
rect 27246 12792 27252 12804
rect 27304 12792 27310 12844
rect 27522 12792 27528 12844
rect 27580 12832 27586 12844
rect 27580 12804 27844 12832
rect 27580 12792 27586 12804
rect 16669 12767 16727 12773
rect 16669 12733 16681 12767
rect 16715 12764 16727 12767
rect 23474 12764 23480 12776
rect 16715 12736 21036 12764
rect 23435 12736 23480 12764
rect 16715 12733 16727 12736
rect 16669 12727 16727 12733
rect 9646 12668 10916 12696
rect 15010 12656 15016 12708
rect 15068 12696 15074 12708
rect 16761 12699 16819 12705
rect 16761 12696 16773 12699
rect 15068 12668 16773 12696
rect 15068 12656 15074 12668
rect 16761 12665 16773 12668
rect 16807 12665 16819 12699
rect 16761 12659 16819 12665
rect 16853 12699 16911 12705
rect 16853 12665 16865 12699
rect 16899 12696 16911 12699
rect 18322 12696 18328 12708
rect 16899 12668 18328 12696
rect 16899 12665 16911 12668
rect 16853 12659 16911 12665
rect 18322 12656 18328 12668
rect 18380 12656 18386 12708
rect 19613 12699 19671 12705
rect 19613 12665 19625 12699
rect 19659 12696 19671 12699
rect 20898 12696 20904 12708
rect 19659 12668 20904 12696
rect 19659 12665 19671 12668
rect 19613 12659 19671 12665
rect 20898 12656 20904 12668
rect 20956 12656 20962 12708
rect 8941 12631 8999 12637
rect 8941 12628 8953 12631
rect 7208 12600 8953 12628
rect 8941 12597 8953 12600
rect 8987 12597 8999 12631
rect 8941 12591 8999 12597
rect 9769 12631 9827 12637
rect 9769 12597 9781 12631
rect 9815 12628 9827 12631
rect 9950 12628 9956 12640
rect 9815 12600 9956 12628
rect 9815 12597 9827 12600
rect 9769 12591 9827 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 13538 12628 13544 12640
rect 13499 12600 13544 12628
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 15102 12588 15108 12640
rect 15160 12628 15166 12640
rect 15289 12631 15347 12637
rect 15289 12628 15301 12631
rect 15160 12600 15301 12628
rect 15160 12588 15166 12600
rect 15289 12597 15301 12600
rect 15335 12597 15347 12631
rect 15289 12591 15347 12597
rect 15657 12631 15715 12637
rect 15657 12597 15669 12631
rect 15703 12628 15715 12631
rect 16022 12628 16028 12640
rect 15703 12600 16028 12628
rect 15703 12597 15715 12600
rect 15657 12591 15715 12597
rect 16022 12588 16028 12600
rect 16080 12588 16086 12640
rect 18506 12628 18512 12640
rect 18467 12600 18512 12628
rect 18506 12588 18512 12600
rect 18564 12588 18570 12640
rect 20070 12588 20076 12640
rect 20128 12628 20134 12640
rect 20254 12628 20260 12640
rect 20128 12600 20260 12628
rect 20128 12588 20134 12600
rect 20254 12588 20260 12600
rect 20312 12588 20318 12640
rect 21008 12628 21036 12736
rect 23474 12724 23480 12736
rect 23532 12724 23538 12776
rect 27706 12764 27712 12776
rect 27667 12736 27712 12764
rect 27706 12724 27712 12736
rect 27764 12724 27770 12776
rect 27816 12773 27844 12804
rect 27890 12792 27896 12844
rect 27948 12832 27954 12844
rect 28166 12832 28172 12844
rect 27948 12804 28172 12832
rect 27948 12792 27954 12804
rect 28166 12792 28172 12804
rect 28224 12832 28230 12844
rect 28445 12835 28503 12841
rect 28445 12832 28457 12835
rect 28224 12804 28457 12832
rect 28224 12792 28230 12804
rect 28445 12801 28457 12804
rect 28491 12801 28503 12835
rect 28445 12795 28503 12801
rect 27801 12767 27859 12773
rect 27801 12733 27813 12767
rect 27847 12764 27859 12767
rect 28258 12764 28264 12776
rect 27847 12736 28264 12764
rect 27847 12733 27859 12736
rect 27801 12727 27859 12733
rect 28258 12724 28264 12736
rect 28316 12724 28322 12776
rect 21358 12656 21364 12708
rect 21416 12696 21422 12708
rect 23385 12699 23443 12705
rect 23385 12696 23397 12699
rect 21416 12668 23397 12696
rect 21416 12656 21422 12668
rect 23385 12665 23397 12668
rect 23431 12665 23443 12699
rect 23385 12659 23443 12665
rect 24578 12628 24584 12640
rect 21008 12600 24584 12628
rect 24578 12588 24584 12600
rect 24636 12588 24642 12640
rect 28626 12628 28632 12640
rect 28587 12600 28632 12628
rect 28626 12588 28632 12600
rect 28684 12588 28690 12640
rect 1104 12538 29440 12560
rect 1104 12486 4492 12538
rect 4544 12486 4556 12538
rect 4608 12486 4620 12538
rect 4672 12486 4684 12538
rect 4736 12486 4748 12538
rect 4800 12486 11576 12538
rect 11628 12486 11640 12538
rect 11692 12486 11704 12538
rect 11756 12486 11768 12538
rect 11820 12486 11832 12538
rect 11884 12486 18660 12538
rect 18712 12486 18724 12538
rect 18776 12486 18788 12538
rect 18840 12486 18852 12538
rect 18904 12486 18916 12538
rect 18968 12486 25744 12538
rect 25796 12486 25808 12538
rect 25860 12486 25872 12538
rect 25924 12486 25936 12538
rect 25988 12486 26000 12538
rect 26052 12486 29440 12538
rect 1104 12464 29440 12486
rect 7466 12424 7472 12436
rect 7379 12396 7472 12424
rect 7466 12384 7472 12396
rect 7524 12424 7530 12436
rect 11698 12424 11704 12436
rect 7524 12396 11704 12424
rect 7524 12384 7530 12396
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12066 12424 12072 12436
rect 12027 12396 12072 12424
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 14458 12424 14464 12436
rect 14200 12396 14464 12424
rect 4706 12356 4712 12368
rect 4356 12328 4712 12356
rect 1762 12248 1768 12300
rect 1820 12288 1826 12300
rect 2041 12291 2099 12297
rect 2041 12288 2053 12291
rect 1820 12260 2053 12288
rect 1820 12248 1826 12260
rect 2041 12257 2053 12260
rect 2087 12257 2099 12291
rect 2041 12251 2099 12257
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 4356 12229 4384 12328
rect 4706 12316 4712 12328
rect 4764 12356 4770 12368
rect 5077 12359 5135 12365
rect 5077 12356 5089 12359
rect 4764 12328 5089 12356
rect 4764 12316 4770 12328
rect 5077 12325 5089 12328
rect 5123 12325 5135 12359
rect 5077 12319 5135 12325
rect 5813 12359 5871 12365
rect 5813 12325 5825 12359
rect 5859 12325 5871 12359
rect 9950 12356 9956 12368
rect 5813 12319 5871 12325
rect 8128 12328 9956 12356
rect 4982 12288 4988 12300
rect 4632 12260 4988 12288
rect 4632 12229 4660 12260
rect 4982 12248 4988 12260
rect 5040 12288 5046 12300
rect 5828 12288 5856 12319
rect 5040 12260 5856 12288
rect 5040 12248 5046 12260
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12189 4399 12223
rect 4341 12183 4399 12189
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12189 4675 12223
rect 5258 12220 5264 12232
rect 5219 12192 5264 12220
rect 4617 12183 4675 12189
rect 5258 12180 5264 12192
rect 5316 12180 5322 12232
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 5810 12220 5816 12232
rect 5399 12192 5488 12220
rect 5771 12192 5816 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 4246 12112 4252 12164
rect 4304 12152 4310 12164
rect 4525 12155 4583 12161
rect 4525 12152 4537 12155
rect 4304 12124 4537 12152
rect 4304 12112 4310 12124
rect 4525 12121 4537 12124
rect 4571 12121 4583 12155
rect 4525 12115 4583 12121
rect 5077 12155 5135 12161
rect 5077 12121 5089 12155
rect 5123 12121 5135 12155
rect 5460 12152 5488 12192
rect 5810 12180 5816 12192
rect 5868 12180 5874 12232
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 7101 12223 7159 12229
rect 5960 12192 6005 12220
rect 5960 12180 5966 12192
rect 7101 12189 7113 12223
rect 7147 12220 7159 12223
rect 7374 12220 7380 12232
rect 7147 12192 7380 12220
rect 7147 12189 7159 12192
rect 7101 12183 7159 12189
rect 7374 12180 7380 12192
rect 7432 12220 7438 12232
rect 8128 12229 8156 12328
rect 9950 12316 9956 12328
rect 10008 12316 10014 12368
rect 14200 12365 14228 12396
rect 14458 12384 14464 12396
rect 14516 12424 14522 12436
rect 14516 12396 15332 12424
rect 14516 12384 14522 12396
rect 10505 12359 10563 12365
rect 10505 12325 10517 12359
rect 10551 12325 10563 12359
rect 10505 12319 10563 12325
rect 11057 12359 11115 12365
rect 11057 12325 11069 12359
rect 11103 12356 11115 12359
rect 14185 12359 14243 12365
rect 11103 12328 12572 12356
rect 11103 12325 11115 12328
rect 11057 12319 11115 12325
rect 9401 12291 9459 12297
rect 9401 12257 9413 12291
rect 9447 12288 9459 12291
rect 10520 12288 10548 12319
rect 9447 12260 10456 12288
rect 10520 12260 12296 12288
rect 9447 12257 9459 12260
rect 9401 12251 9459 12257
rect 7929 12223 7987 12229
rect 7929 12220 7941 12223
rect 7432 12192 7941 12220
rect 7432 12180 7438 12192
rect 7929 12189 7941 12192
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 5920 12152 5948 12180
rect 5460 12124 5948 12152
rect 6089 12155 6147 12161
rect 5077 12115 5135 12121
rect 6089 12121 6101 12155
rect 6135 12152 6147 12155
rect 7006 12152 7012 12164
rect 6135 12124 7012 12152
rect 6135 12121 6147 12124
rect 6089 12115 6147 12121
rect 2501 12087 2559 12093
rect 2501 12053 2513 12087
rect 2547 12084 2559 12087
rect 2590 12084 2596 12096
rect 2547 12056 2596 12084
rect 2547 12053 2559 12056
rect 2501 12047 2559 12053
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 4157 12087 4215 12093
rect 4157 12053 4169 12087
rect 4203 12084 4215 12087
rect 4338 12084 4344 12096
rect 4203 12056 4344 12084
rect 4203 12053 4215 12056
rect 4157 12047 4215 12053
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 5092 12084 5120 12115
rect 6104 12084 6132 12115
rect 7006 12112 7012 12124
rect 7064 12112 7070 12164
rect 7285 12155 7343 12161
rect 7285 12121 7297 12155
rect 7331 12152 7343 12155
rect 8128 12152 8156 12183
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9824 12192 9873 12220
rect 9824 12180 9830 12192
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 9954 12223 10012 12229
rect 9954 12189 9966 12223
rect 10000 12189 10012 12223
rect 9954 12183 10012 12189
rect 7331 12124 8156 12152
rect 8297 12155 8355 12161
rect 7331 12121 7343 12124
rect 7285 12115 7343 12121
rect 8297 12121 8309 12155
rect 8343 12152 8355 12155
rect 9968 12152 9996 12183
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 10428 12230 10456 12260
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 10100 12192 10241 12220
rect 10100 12180 10106 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10326 12223 10384 12229
rect 10326 12189 10338 12223
rect 10372 12220 10384 12223
rect 10428 12220 10548 12230
rect 10686 12220 10692 12232
rect 10372 12202 10692 12220
rect 10372 12192 10456 12202
rect 10520 12192 10692 12202
rect 10372 12189 10384 12192
rect 10326 12183 10384 12189
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 10962 12220 10968 12232
rect 10836 12192 10968 12220
rect 10836 12180 10842 12192
rect 10962 12180 10968 12192
rect 11020 12220 11026 12232
rect 11241 12223 11299 12229
rect 11241 12220 11253 12223
rect 11020 12192 11253 12220
rect 11020 12180 11026 12192
rect 11241 12189 11253 12192
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 11514 12220 11520 12232
rect 11388 12192 11433 12220
rect 11475 12192 11520 12220
rect 11388 12180 11394 12192
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 11609 12201 11667 12207
rect 11609 12167 11621 12201
rect 11655 12167 11667 12201
rect 11698 12180 11704 12232
rect 11756 12220 11762 12232
rect 12268 12229 12296 12260
rect 12544 12229 12572 12328
rect 14185 12325 14197 12359
rect 14231 12325 14243 12359
rect 15102 12356 15108 12368
rect 14185 12319 14243 12325
rect 14292 12328 15108 12356
rect 14292 12288 14320 12328
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 15304 12356 15332 12396
rect 15838 12384 15844 12436
rect 15896 12424 15902 12436
rect 16482 12424 16488 12436
rect 15896 12396 16488 12424
rect 15896 12384 15902 12396
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 18506 12384 18512 12436
rect 18564 12424 18570 12436
rect 19518 12424 19524 12436
rect 18564 12396 19524 12424
rect 18564 12384 18570 12396
rect 19518 12384 19524 12396
rect 19576 12384 19582 12436
rect 19613 12427 19671 12433
rect 19613 12393 19625 12427
rect 19659 12424 19671 12427
rect 20070 12424 20076 12436
rect 19659 12396 20076 12424
rect 19659 12393 19671 12396
rect 19613 12387 19671 12393
rect 20070 12384 20076 12396
rect 20128 12424 20134 12436
rect 20254 12424 20260 12436
rect 20128 12396 20260 12424
rect 20128 12384 20134 12396
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 26142 12424 26148 12436
rect 26103 12396 26148 12424
rect 26142 12384 26148 12396
rect 26200 12384 26206 12436
rect 15304 12328 16344 12356
rect 13372 12260 14320 12288
rect 14369 12291 14427 12297
rect 13372 12232 13400 12260
rect 14369 12257 14381 12291
rect 14415 12288 14427 12291
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 14415 12260 14841 12288
rect 14415 12257 14427 12260
rect 14369 12251 14427 12257
rect 14829 12257 14841 12260
rect 14875 12257 14887 12291
rect 15378 12288 15384 12300
rect 14829 12251 14887 12257
rect 15028 12260 15384 12288
rect 12253 12223 12311 12229
rect 11756 12192 12112 12220
rect 11756 12180 11762 12192
rect 10134 12152 10140 12164
rect 8343 12124 9996 12152
rect 10095 12124 10140 12152
rect 8343 12121 8355 12124
rect 8297 12115 8355 12121
rect 5092 12056 6132 12084
rect 6641 12087 6699 12093
rect 6641 12053 6653 12087
rect 6687 12084 6699 12087
rect 6730 12084 6736 12096
rect 6687 12056 6736 12084
rect 6687 12053 6699 12056
rect 6641 12047 6699 12053
rect 6730 12044 6736 12056
rect 6788 12084 6794 12096
rect 7300 12084 7328 12115
rect 6788 12056 7328 12084
rect 6788 12044 6794 12056
rect 7926 12044 7932 12096
rect 7984 12084 7990 12096
rect 8312 12084 8340 12115
rect 10134 12112 10140 12124
rect 10192 12112 10198 12164
rect 11609 12161 11667 12167
rect 7984 12056 8340 12084
rect 7984 12044 7990 12056
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10152 12084 10180 12112
rect 9732 12056 10180 12084
rect 9732 12044 9738 12056
rect 11514 12044 11520 12096
rect 11572 12084 11578 12096
rect 11624 12084 11652 12161
rect 12084 12152 12112 12192
rect 12253 12189 12265 12223
rect 12299 12189 12311 12223
rect 12253 12183 12311 12189
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 12360 12152 12388 12183
rect 12618 12180 12624 12232
rect 12676 12220 12682 12232
rect 12676 12192 12721 12220
rect 12676 12180 12682 12192
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 13354 12220 13360 12232
rect 13044 12192 13360 12220
rect 13044 12180 13050 12192
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 13814 12220 13820 12232
rect 13587 12192 13820 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 15028 12229 15056 12260
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 15013 12223 15071 12229
rect 15013 12189 15025 12223
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 15197 12223 15255 12229
rect 15197 12189 15209 12223
rect 15243 12189 15255 12223
rect 15197 12183 15255 12189
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 15562 12220 15568 12232
rect 15335 12192 15568 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 12084 12124 12388 12152
rect 14108 12152 14136 12183
rect 14550 12152 14556 12164
rect 14108 12124 14556 12152
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 15212 12152 15240 12183
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 16022 12220 16028 12232
rect 15983 12192 16028 12220
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 16316 12229 16344 12328
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 22094 12356 22100 12368
rect 16448 12328 22100 12356
rect 16448 12316 16454 12328
rect 22094 12316 22100 12328
rect 22152 12316 22158 12368
rect 26881 12359 26939 12365
rect 23952 12328 26832 12356
rect 16408 12229 16436 12316
rect 20073 12291 20131 12297
rect 20073 12288 20085 12291
rect 19444 12260 20085 12288
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12189 16359 12223
rect 16301 12183 16359 12189
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 15378 12152 15384 12164
rect 15212 12124 15384 12152
rect 15378 12112 15384 12124
rect 15436 12112 15442 12164
rect 16224 12152 16252 12183
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 16540 12192 19288 12220
rect 16540 12180 16546 12192
rect 17862 12152 17868 12164
rect 16224 12124 17868 12152
rect 17862 12112 17868 12124
rect 17920 12112 17926 12164
rect 19260 12152 19288 12192
rect 19334 12180 19340 12232
rect 19392 12220 19398 12232
rect 19444 12229 19472 12260
rect 20073 12257 20085 12260
rect 20119 12257 20131 12291
rect 20073 12251 20131 12257
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 19392 12192 19441 12220
rect 19392 12180 19398 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19518 12180 19524 12232
rect 19576 12220 19582 12232
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 19576 12192 19625 12220
rect 19576 12180 19582 12192
rect 19613 12189 19625 12192
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 20806 12152 20812 12164
rect 19260 12124 20812 12152
rect 20806 12112 20812 12124
rect 20864 12152 20870 12164
rect 21177 12155 21235 12161
rect 21177 12152 21189 12155
rect 20864 12124 21189 12152
rect 20864 12112 20870 12124
rect 21177 12121 21189 12124
rect 21223 12121 21235 12155
rect 21177 12115 21235 12121
rect 22094 12112 22100 12164
rect 22152 12152 22158 12164
rect 22830 12152 22836 12164
rect 22152 12124 22836 12152
rect 22152 12112 22158 12124
rect 22830 12112 22836 12124
rect 22888 12112 22894 12164
rect 11572 12056 11652 12084
rect 13449 12087 13507 12093
rect 11572 12044 11578 12056
rect 13449 12053 13461 12087
rect 13495 12084 13507 12087
rect 13630 12084 13636 12096
rect 13495 12056 13636 12084
rect 13495 12053 13507 12056
rect 13449 12047 13507 12053
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 14369 12087 14427 12093
rect 14369 12053 14381 12087
rect 14415 12084 14427 12087
rect 14734 12084 14740 12096
rect 14415 12056 14740 12084
rect 14415 12053 14427 12056
rect 14369 12047 14427 12053
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 16666 12084 16672 12096
rect 16627 12056 16672 12084
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 17770 12084 17776 12096
rect 17731 12056 17776 12084
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 18506 12044 18512 12096
rect 18564 12084 18570 12096
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 18564 12056 18613 12084
rect 18564 12044 18570 12056
rect 18601 12053 18613 12056
rect 18647 12053 18659 12087
rect 19242 12084 19248 12096
rect 19203 12056 19248 12084
rect 18601 12047 18659 12053
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 23952 12084 23980 12328
rect 24854 12248 24860 12300
rect 24912 12288 24918 12300
rect 25498 12288 25504 12300
rect 24912 12260 25504 12288
rect 24912 12248 24918 12260
rect 25498 12248 25504 12260
rect 25556 12248 25562 12300
rect 26804 12288 26832 12328
rect 26881 12325 26893 12359
rect 26927 12356 26939 12359
rect 28166 12356 28172 12368
rect 26927 12328 28172 12356
rect 26927 12325 26939 12328
rect 26881 12319 26939 12325
rect 28166 12316 28172 12328
rect 28224 12316 28230 12368
rect 27985 12291 28043 12297
rect 26804 12260 27936 12288
rect 25222 12220 25228 12232
rect 25183 12192 25228 12220
rect 25222 12180 25228 12192
rect 25280 12180 25286 12232
rect 26142 12180 26148 12232
rect 26200 12220 26206 12232
rect 27801 12223 27859 12229
rect 27801 12220 27813 12223
rect 26200 12192 27813 12220
rect 26200 12180 26206 12192
rect 27801 12189 27813 12192
rect 27847 12189 27859 12223
rect 27801 12183 27859 12189
rect 24670 12112 24676 12164
rect 24728 12152 24734 12164
rect 26694 12152 26700 12164
rect 24728 12124 25360 12152
rect 26655 12124 26700 12152
rect 24728 12112 24734 12124
rect 19392 12056 23980 12084
rect 19392 12044 19398 12056
rect 24026 12044 24032 12096
rect 24084 12084 24090 12096
rect 25332 12093 25360 12124
rect 26694 12112 26700 12124
rect 26752 12112 26758 12164
rect 27709 12155 27767 12161
rect 27709 12121 27721 12155
rect 27755 12152 27767 12155
rect 27908 12152 27936 12260
rect 27985 12257 27997 12291
rect 28031 12288 28043 12291
rect 28074 12288 28080 12300
rect 28031 12260 28080 12288
rect 28031 12257 28043 12260
rect 27985 12251 28043 12257
rect 28074 12248 28080 12260
rect 28132 12248 28138 12300
rect 28350 12152 28356 12164
rect 27755 12124 28356 12152
rect 27755 12121 27767 12124
rect 27709 12115 27767 12121
rect 28350 12112 28356 12124
rect 28408 12152 28414 12164
rect 28537 12155 28595 12161
rect 28537 12152 28549 12155
rect 28408 12124 28549 12152
rect 28408 12112 28414 12124
rect 28537 12121 28549 12124
rect 28583 12121 28595 12155
rect 28537 12115 28595 12121
rect 24857 12087 24915 12093
rect 24857 12084 24869 12087
rect 24084 12056 24869 12084
rect 24084 12044 24090 12056
rect 24857 12053 24869 12056
rect 24903 12053 24915 12087
rect 24857 12047 24915 12053
rect 25317 12087 25375 12093
rect 25317 12053 25329 12087
rect 25363 12084 25375 12087
rect 26142 12084 26148 12096
rect 25363 12056 26148 12084
rect 25363 12053 25375 12056
rect 25317 12047 25375 12053
rect 26142 12044 26148 12056
rect 26200 12044 26206 12096
rect 27341 12087 27399 12093
rect 27341 12053 27353 12087
rect 27387 12084 27399 12087
rect 27614 12084 27620 12096
rect 27387 12056 27620 12084
rect 27387 12053 27399 12056
rect 27341 12047 27399 12053
rect 27614 12044 27620 12056
rect 27672 12044 27678 12096
rect 1104 11994 29600 12016
rect 1104 11942 8034 11994
rect 8086 11942 8098 11994
rect 8150 11942 8162 11994
rect 8214 11942 8226 11994
rect 8278 11942 8290 11994
rect 8342 11942 15118 11994
rect 15170 11942 15182 11994
rect 15234 11942 15246 11994
rect 15298 11942 15310 11994
rect 15362 11942 15374 11994
rect 15426 11942 22202 11994
rect 22254 11942 22266 11994
rect 22318 11942 22330 11994
rect 22382 11942 22394 11994
rect 22446 11942 22458 11994
rect 22510 11942 29286 11994
rect 29338 11942 29350 11994
rect 29402 11942 29414 11994
rect 29466 11942 29478 11994
rect 29530 11942 29542 11994
rect 29594 11942 29600 11994
rect 1104 11920 29600 11942
rect 3050 11840 3056 11892
rect 3108 11880 3114 11892
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 3108 11852 3157 11880
rect 3108 11840 3114 11852
rect 3145 11849 3157 11852
rect 3191 11849 3203 11883
rect 3145 11843 3203 11849
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 5316 11852 5457 11880
rect 5316 11840 5322 11852
rect 5445 11849 5457 11852
rect 5491 11880 5503 11883
rect 5810 11880 5816 11892
rect 5491 11852 5816 11880
rect 5491 11849 5503 11852
rect 5445 11843 5503 11849
rect 5810 11840 5816 11852
rect 5868 11880 5874 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 5868 11852 6377 11880
rect 5868 11840 5874 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6380 11812 6408 11843
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 7285 11883 7343 11889
rect 7285 11880 7297 11883
rect 7064 11852 7297 11880
rect 7064 11840 7070 11852
rect 7285 11849 7297 11852
rect 7331 11849 7343 11883
rect 7285 11843 7343 11849
rect 8754 11840 8760 11892
rect 8812 11880 8818 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 8812 11852 9229 11880
rect 8812 11840 8818 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 9217 11843 9275 11849
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 10318 11880 10324 11892
rect 9824 11852 10324 11880
rect 9824 11840 9830 11852
rect 10318 11840 10324 11852
rect 10376 11880 10382 11892
rect 10873 11883 10931 11889
rect 10873 11880 10885 11883
rect 10376 11852 10885 11880
rect 10376 11840 10382 11852
rect 10873 11849 10885 11852
rect 10919 11849 10931 11883
rect 11514 11880 11520 11892
rect 11475 11852 11520 11880
rect 10873 11843 10931 11849
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 14550 11880 14556 11892
rect 14511 11852 14556 11880
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 18414 11840 18420 11892
rect 18472 11880 18478 11892
rect 19334 11880 19340 11892
rect 18472 11852 19340 11880
rect 18472 11840 18478 11852
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 20714 11880 20720 11892
rect 20548 11852 20720 11880
rect 8478 11812 8484 11824
rect 6380 11784 8484 11812
rect 8478 11772 8484 11784
rect 8536 11812 8542 11824
rect 8665 11815 8723 11821
rect 8665 11812 8677 11815
rect 8536 11784 8677 11812
rect 8536 11772 8542 11784
rect 8665 11781 8677 11784
rect 8711 11781 8723 11815
rect 10410 11812 10416 11824
rect 10371 11784 10416 11812
rect 8665 11775 8723 11781
rect 10410 11772 10416 11784
rect 10468 11812 10474 11824
rect 11054 11812 11060 11824
rect 10468 11784 11060 11812
rect 10468 11772 10474 11784
rect 11054 11772 11060 11784
rect 11112 11812 11118 11824
rect 11669 11815 11727 11821
rect 11669 11812 11681 11815
rect 11112 11784 11681 11812
rect 11112 11772 11118 11784
rect 11669 11781 11681 11784
rect 11715 11781 11727 11815
rect 11669 11775 11727 11781
rect 11885 11815 11943 11821
rect 11885 11781 11897 11815
rect 11931 11812 11943 11815
rect 18506 11812 18512 11824
rect 11931 11784 18512 11812
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 2314 11744 2320 11756
rect 2275 11716 2320 11744
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 2590 11744 2596 11756
rect 2551 11716 2596 11744
rect 2590 11704 2596 11716
rect 2648 11704 2654 11756
rect 4982 11744 4988 11756
rect 4943 11716 4988 11744
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11713 7343 11747
rect 7466 11744 7472 11756
rect 7427 11716 7472 11744
rect 7285 11707 7343 11713
rect 7300 11676 7328 11707
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10870 11744 10876 11756
rect 10100 11716 10876 11744
rect 10100 11704 10106 11716
rect 10870 11704 10876 11716
rect 10928 11744 10934 11756
rect 11900 11744 11928 11775
rect 18506 11772 18512 11784
rect 18564 11772 18570 11824
rect 12802 11744 12808 11756
rect 10928 11716 11928 11744
rect 12763 11716 12808 11744
rect 10928 11704 10934 11716
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 12986 11744 12992 11756
rect 12947 11716 12992 11744
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13170 11744 13176 11756
rect 13127 11716 13176 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11744 13323 11747
rect 13722 11744 13728 11756
rect 13311 11716 13728 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 17034 11744 17040 11756
rect 16995 11716 17040 11744
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 17310 11744 17316 11756
rect 17271 11716 17316 11744
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 18414 11744 18420 11756
rect 18375 11716 18420 11744
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 19242 11744 19248 11756
rect 19203 11716 19248 11744
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 20548 11753 20576 11852
rect 20714 11840 20720 11852
rect 20772 11840 20778 11892
rect 20806 11840 20812 11892
rect 20864 11880 20870 11892
rect 20864 11852 22692 11880
rect 20864 11840 20870 11852
rect 22296 11821 22324 11852
rect 22097 11815 22155 11821
rect 22097 11812 22109 11815
rect 20640 11784 22109 11812
rect 20640 11753 20668 11784
rect 22097 11781 22109 11784
rect 22143 11781 22155 11815
rect 22097 11775 22155 11781
rect 22281 11815 22339 11821
rect 22281 11781 22293 11815
rect 22327 11812 22339 11815
rect 22664 11812 22692 11852
rect 22830 11840 22836 11892
rect 22888 11880 22894 11892
rect 23290 11880 23296 11892
rect 22888 11852 23296 11880
rect 22888 11840 22894 11852
rect 23290 11840 23296 11852
rect 23348 11840 23354 11892
rect 23474 11840 23480 11892
rect 23532 11880 23538 11892
rect 24489 11883 24547 11889
rect 24489 11880 24501 11883
rect 23532 11852 24501 11880
rect 23532 11840 23538 11852
rect 24489 11849 24501 11852
rect 24535 11849 24547 11883
rect 27246 11880 27252 11892
rect 27207 11852 27252 11880
rect 24489 11843 24547 11849
rect 27246 11840 27252 11852
rect 27304 11840 27310 11892
rect 27617 11883 27675 11889
rect 27617 11849 27629 11883
rect 27663 11880 27675 11883
rect 27706 11880 27712 11892
rect 27663 11852 27712 11880
rect 27663 11849 27675 11852
rect 27617 11843 27675 11849
rect 27706 11840 27712 11852
rect 27764 11840 27770 11892
rect 28074 11840 28080 11892
rect 28132 11880 28138 11892
rect 28445 11883 28503 11889
rect 28445 11880 28457 11883
rect 28132 11852 28457 11880
rect 28132 11840 28138 11852
rect 28445 11849 28457 11852
rect 28491 11849 28503 11883
rect 28445 11843 28503 11849
rect 23750 11812 23756 11824
rect 22327 11784 22361 11812
rect 22664 11784 23756 11812
rect 22327 11781 22339 11784
rect 22281 11775 22339 11781
rect 23750 11772 23756 11784
rect 23808 11772 23814 11824
rect 24578 11772 24584 11824
rect 24636 11812 24642 11824
rect 24636 11784 25084 11812
rect 24636 11772 24642 11784
rect 20533 11747 20591 11753
rect 20533 11744 20545 11747
rect 20496 11716 20545 11744
rect 20496 11704 20502 11716
rect 20533 11713 20545 11716
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11713 20683 11747
rect 20806 11744 20812 11756
rect 20767 11716 20812 11744
rect 20625 11707 20683 11713
rect 7926 11676 7932 11688
rect 7300 11648 7932 11676
rect 7926 11636 7932 11648
rect 7984 11636 7990 11688
rect 19150 11676 19156 11688
rect 19111 11648 19156 11676
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 19886 11636 19892 11688
rect 19944 11676 19950 11688
rect 20640 11676 20668 11707
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 20898 11704 20904 11756
rect 20956 11744 20962 11756
rect 23014 11744 23020 11756
rect 20956 11716 21001 11744
rect 22066 11716 23020 11744
rect 20956 11704 20962 11716
rect 19944 11648 20668 11676
rect 21085 11679 21143 11685
rect 19944 11636 19950 11648
rect 21085 11645 21097 11679
rect 21131 11676 21143 11679
rect 22066 11676 22094 11716
rect 23014 11704 23020 11716
rect 23072 11704 23078 11756
rect 23201 11747 23259 11753
rect 23201 11713 23213 11747
rect 23247 11713 23259 11747
rect 23201 11707 23259 11713
rect 21131 11648 22094 11676
rect 22465 11679 22523 11685
rect 21131 11645 21143 11648
rect 21085 11639 21143 11645
rect 22465 11645 22477 11679
rect 22511 11676 22523 11679
rect 23216 11676 23244 11707
rect 23658 11704 23664 11756
rect 23716 11744 23722 11756
rect 23842 11744 23848 11756
rect 23716 11716 23848 11744
rect 23716 11704 23722 11716
rect 23842 11704 23848 11716
rect 23900 11704 23906 11756
rect 24026 11744 24032 11756
rect 23987 11716 24032 11744
rect 24026 11704 24032 11716
rect 24084 11704 24090 11756
rect 24670 11744 24676 11756
rect 24631 11716 24676 11744
rect 24670 11704 24676 11716
rect 24728 11704 24734 11756
rect 24762 11704 24768 11756
rect 24820 11744 24826 11756
rect 24946 11744 24952 11756
rect 24820 11716 24865 11744
rect 24907 11716 24952 11744
rect 24820 11704 24826 11716
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 25056 11753 25084 11784
rect 25041 11747 25099 11753
rect 25041 11713 25053 11747
rect 25087 11713 25099 11747
rect 25041 11707 25099 11713
rect 23290 11676 23296 11688
rect 22511 11648 23296 11676
rect 22511 11645 22523 11648
rect 22465 11639 22523 11645
rect 23290 11636 23296 11648
rect 23348 11636 23354 11688
rect 23385 11679 23443 11685
rect 23385 11645 23397 11679
rect 23431 11676 23443 11679
rect 26694 11676 26700 11688
rect 23431 11648 26700 11676
rect 23431 11645 23443 11648
rect 23385 11639 23443 11645
rect 26694 11636 26700 11648
rect 26752 11636 26758 11688
rect 27706 11676 27712 11688
rect 27667 11648 27712 11676
rect 27706 11636 27712 11648
rect 27764 11636 27770 11688
rect 27893 11679 27951 11685
rect 27893 11645 27905 11679
rect 27939 11676 27951 11679
rect 28258 11676 28264 11688
rect 27939 11648 28264 11676
rect 27939 11645 27951 11648
rect 27893 11639 27951 11645
rect 28258 11636 28264 11648
rect 28316 11636 28322 11688
rect 12897 11611 12955 11617
rect 12897 11577 12909 11611
rect 12943 11608 12955 11611
rect 13906 11608 13912 11620
rect 12943 11580 13912 11608
rect 12943 11577 12955 11580
rect 12897 11571 12955 11577
rect 13906 11568 13912 11580
rect 13964 11568 13970 11620
rect 17497 11611 17555 11617
rect 17497 11577 17509 11611
rect 17543 11608 17555 11611
rect 17586 11608 17592 11620
rect 17543 11580 17592 11608
rect 17543 11577 17555 11580
rect 17497 11571 17555 11577
rect 17586 11568 17592 11580
rect 17644 11568 17650 11620
rect 19242 11608 19248 11620
rect 19203 11580 19248 11608
rect 19242 11568 19248 11580
rect 19300 11568 19306 11620
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4525 11543 4583 11549
rect 4525 11540 4537 11543
rect 4304 11512 4537 11540
rect 4304 11500 4310 11512
rect 4525 11509 4537 11512
rect 4571 11509 4583 11543
rect 4706 11540 4712 11552
rect 4667 11512 4712 11540
rect 4525 11503 4583 11509
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 7929 11543 7987 11549
rect 7929 11540 7941 11543
rect 6788 11512 7941 11540
rect 6788 11500 6794 11512
rect 7929 11509 7941 11512
rect 7975 11509 7987 11543
rect 7929 11503 7987 11509
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 10134 11540 10140 11552
rect 9907 11512 10140 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 10134 11500 10140 11512
rect 10192 11540 10198 11552
rect 10962 11540 10968 11552
rect 10192 11512 10968 11540
rect 10192 11500 10198 11512
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 11388 11512 11713 11540
rect 11388 11500 11394 11512
rect 11701 11509 11713 11512
rect 11747 11509 11759 11543
rect 11701 11503 11759 11509
rect 12621 11543 12679 11549
rect 12621 11509 12633 11543
rect 12667 11540 12679 11543
rect 12802 11540 12808 11552
rect 12667 11512 12808 11540
rect 12667 11509 12679 11512
rect 12621 11503 12679 11509
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 13722 11540 13728 11552
rect 13683 11512 13728 11540
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 20070 11540 20076 11552
rect 20031 11512 20076 11540
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 23934 11540 23940 11552
rect 23895 11512 23940 11540
rect 23934 11500 23940 11512
rect 23992 11500 23998 11552
rect 1104 11450 29440 11472
rect 1104 11398 4492 11450
rect 4544 11398 4556 11450
rect 4608 11398 4620 11450
rect 4672 11398 4684 11450
rect 4736 11398 4748 11450
rect 4800 11398 11576 11450
rect 11628 11398 11640 11450
rect 11692 11398 11704 11450
rect 11756 11398 11768 11450
rect 11820 11398 11832 11450
rect 11884 11398 18660 11450
rect 18712 11398 18724 11450
rect 18776 11398 18788 11450
rect 18840 11398 18852 11450
rect 18904 11398 18916 11450
rect 18968 11398 25744 11450
rect 25796 11398 25808 11450
rect 25860 11398 25872 11450
rect 25924 11398 25936 11450
rect 25988 11398 26000 11450
rect 26052 11398 29440 11450
rect 1104 11376 29440 11398
rect 1762 11336 1768 11348
rect 1723 11308 1768 11336
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 17218 11336 17224 11348
rect 17179 11308 17224 11336
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 17770 11336 17776 11348
rect 17328 11308 17776 11336
rect 4525 11271 4583 11277
rect 4525 11237 4537 11271
rect 4571 11268 4583 11271
rect 5626 11268 5632 11280
rect 4571 11240 5632 11268
rect 4571 11237 4583 11240
rect 4525 11231 4583 11237
rect 5626 11228 5632 11240
rect 5684 11228 5690 11280
rect 9858 11228 9864 11280
rect 9916 11268 9922 11280
rect 17328 11268 17356 11308
rect 17770 11296 17776 11308
rect 17828 11336 17834 11348
rect 18325 11339 18383 11345
rect 18325 11336 18337 11339
rect 17828 11308 18337 11336
rect 17828 11296 17834 11308
rect 18325 11305 18337 11308
rect 18371 11305 18383 11339
rect 18325 11299 18383 11305
rect 18506 11296 18512 11348
rect 18564 11336 18570 11348
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 18564 11308 19257 11336
rect 18564 11296 18570 11308
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 19245 11299 19303 11305
rect 19705 11339 19763 11345
rect 19705 11305 19717 11339
rect 19751 11336 19763 11339
rect 19886 11336 19892 11348
rect 19751 11308 19892 11336
rect 19751 11305 19763 11308
rect 19705 11299 19763 11305
rect 9916 11240 17356 11268
rect 18141 11271 18199 11277
rect 9916 11228 9922 11240
rect 18141 11237 18153 11271
rect 18187 11268 18199 11271
rect 19150 11268 19156 11280
rect 18187 11240 19156 11268
rect 18187 11237 18199 11240
rect 18141 11231 18199 11237
rect 19150 11228 19156 11240
rect 19208 11228 19214 11280
rect 19260 11268 19288 11299
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 20070 11296 20076 11348
rect 20128 11336 20134 11348
rect 21269 11339 21327 11345
rect 21269 11336 21281 11339
rect 20128 11308 21281 11336
rect 20128 11296 20134 11308
rect 21269 11305 21281 11308
rect 21315 11305 21327 11339
rect 21269 11299 21327 11305
rect 22649 11339 22707 11345
rect 22649 11305 22661 11339
rect 22695 11336 22707 11339
rect 23750 11336 23756 11348
rect 22695 11308 23756 11336
rect 22695 11305 22707 11308
rect 22649 11299 22707 11305
rect 23750 11296 23756 11308
rect 23808 11296 23814 11348
rect 24489 11339 24547 11345
rect 24489 11305 24501 11339
rect 24535 11336 24547 11339
rect 24762 11336 24768 11348
rect 24535 11308 24768 11336
rect 24535 11305 24547 11308
rect 24489 11299 24547 11305
rect 24762 11296 24768 11308
rect 24820 11296 24826 11348
rect 27614 11336 27620 11348
rect 27575 11308 27620 11336
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 27709 11339 27767 11345
rect 27709 11305 27721 11339
rect 27755 11336 27767 11339
rect 27798 11336 27804 11348
rect 27755 11308 27804 11336
rect 27755 11305 27767 11308
rect 27709 11299 27767 11305
rect 27798 11296 27804 11308
rect 27856 11296 27862 11348
rect 20717 11271 20775 11277
rect 20717 11268 20729 11271
rect 19260 11240 20729 11268
rect 20717 11237 20729 11240
rect 20763 11237 20775 11271
rect 20717 11231 20775 11237
rect 23201 11271 23259 11277
rect 23201 11237 23213 11271
rect 23247 11268 23259 11271
rect 23382 11268 23388 11280
rect 23247 11240 23388 11268
rect 23247 11237 23259 11240
rect 23201 11231 23259 11237
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11200 2283 11203
rect 4617 11203 4675 11209
rect 2271 11172 2774 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 2130 11132 2136 11144
rect 2091 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 2746 11064 2774 11172
rect 4617 11169 4629 11203
rect 4663 11200 4675 11203
rect 4890 11200 4896 11212
rect 4663 11172 4896 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 8021 11203 8079 11209
rect 8021 11200 8033 11203
rect 7892 11172 8033 11200
rect 7892 11160 7898 11172
rect 8021 11169 8033 11172
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11200 8263 11203
rect 9030 11200 9036 11212
rect 8251 11172 9036 11200
rect 8251 11169 8263 11172
rect 8205 11163 8263 11169
rect 9030 11160 9036 11172
rect 9088 11160 9094 11212
rect 10413 11203 10471 11209
rect 10413 11200 10425 11203
rect 9646 11172 10425 11200
rect 4246 11132 4252 11144
rect 4207 11104 4252 11132
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11132 4399 11135
rect 4798 11132 4804 11144
rect 4387 11104 4804 11132
rect 4387 11101 4399 11104
rect 4341 11095 4399 11101
rect 4798 11092 4804 11104
rect 4856 11132 4862 11144
rect 5166 11132 5172 11144
rect 4856 11104 5172 11132
rect 4856 11092 4862 11104
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 7926 11132 7932 11144
rect 7887 11104 7932 11132
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8386 11132 8392 11144
rect 8159 11104 8392 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8386 11092 8392 11104
rect 8444 11132 8450 11144
rect 8662 11132 8668 11144
rect 8444 11104 8668 11132
rect 8444 11092 8450 11104
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8772 11104 8953 11132
rect 2869 11067 2927 11073
rect 2869 11064 2881 11067
rect 2746 11036 2881 11064
rect 2869 11033 2881 11036
rect 2915 11064 2927 11067
rect 3326 11064 3332 11076
rect 2915 11036 3332 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 3326 11024 3332 11036
rect 3384 11024 3390 11076
rect 4706 11064 4712 11076
rect 4448 11036 4712 11064
rect 4448 11005 4476 11036
rect 4706 11024 4712 11036
rect 4764 11064 4770 11076
rect 5074 11064 5080 11076
rect 4764 11036 5080 11064
rect 4764 11024 4770 11036
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 6730 11024 6736 11076
rect 6788 11064 6794 11076
rect 7193 11067 7251 11073
rect 7193 11064 7205 11067
rect 6788 11036 7205 11064
rect 6788 11024 6794 11036
rect 7193 11033 7205 11036
rect 7239 11064 7251 11067
rect 8772 11064 8800 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9646 11132 9674 11172
rect 10413 11169 10425 11172
rect 10459 11200 10471 11203
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 10459 11172 10977 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10965 11169 10977 11172
rect 11011 11200 11023 11203
rect 11330 11200 11336 11212
rect 11011 11172 11336 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 12894 11200 12900 11212
rect 12855 11172 12900 11200
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11200 13047 11203
rect 13538 11200 13544 11212
rect 13035 11172 13544 11200
rect 13035 11169 13047 11172
rect 12989 11163 13047 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11200 14519 11203
rect 15010 11200 15016 11212
rect 14507 11172 15016 11200
rect 14507 11169 14519 11172
rect 14461 11163 14519 11169
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 18506 11160 18512 11212
rect 18564 11200 18570 11212
rect 19337 11203 19395 11209
rect 19337 11200 19349 11203
rect 18564 11172 19349 11200
rect 18564 11160 18570 11172
rect 19337 11169 19349 11172
rect 19383 11169 19395 11203
rect 19337 11163 19395 11169
rect 21266 11160 21272 11212
rect 21324 11200 21330 11212
rect 21821 11203 21879 11209
rect 21821 11200 21833 11203
rect 21324 11172 21833 11200
rect 21324 11160 21330 11172
rect 21821 11169 21833 11172
rect 21867 11169 21879 11203
rect 21821 11163 21879 11169
rect 27154 11160 27160 11212
rect 27212 11200 27218 11212
rect 27801 11203 27859 11209
rect 27801 11200 27813 11203
rect 27212 11172 27813 11200
rect 27212 11160 27218 11172
rect 27801 11169 27813 11172
rect 27847 11200 27859 11203
rect 28166 11200 28172 11212
rect 27847 11172 28172 11200
rect 27847 11169 27859 11172
rect 27801 11163 27859 11169
rect 28166 11160 28172 11172
rect 28224 11160 28230 11212
rect 9180 11104 9273 11132
rect 9600 11104 9674 11132
rect 9180 11092 9186 11104
rect 7239 11036 8800 11064
rect 7239 11033 7251 11036
rect 7193 11027 7251 11033
rect 8846 11024 8852 11076
rect 8904 11064 8910 11076
rect 9140 11064 9168 11092
rect 9600 11073 9628 11104
rect 10686 11092 10692 11144
rect 10744 11132 10750 11144
rect 13081 11135 13139 11141
rect 10744 11104 12940 11132
rect 10744 11092 10750 11104
rect 12912 11076 12940 11104
rect 13081 11101 13093 11135
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 9585 11067 9643 11073
rect 9585 11064 9597 11067
rect 8904 11036 9597 11064
rect 8904 11024 8910 11036
rect 9585 11033 9597 11036
rect 9631 11033 9643 11067
rect 9585 11027 9643 11033
rect 9766 11024 9772 11076
rect 9824 11064 9830 11076
rect 10778 11064 10784 11076
rect 9824 11036 10784 11064
rect 9824 11024 9830 11036
rect 10778 11024 10784 11036
rect 10836 11064 10842 11076
rect 11701 11067 11759 11073
rect 11701 11064 11713 11067
rect 10836 11036 11713 11064
rect 10836 11024 10842 11036
rect 11701 11033 11713 11036
rect 11747 11064 11759 11067
rect 11747 11036 12848 11064
rect 11747 11033 11759 11036
rect 11701 11027 11759 11033
rect 4433 10999 4491 11005
rect 4433 10965 4445 10999
rect 4479 10965 4491 10999
rect 4433 10959 4491 10965
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 7745 10999 7803 11005
rect 7745 10996 7757 10999
rect 7708 10968 7757 10996
rect 7708 10956 7714 10968
rect 7745 10965 7757 10968
rect 7791 10965 7803 10999
rect 12710 10996 12716 11008
rect 12671 10968 12716 10996
rect 7745 10959 7803 10965
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 12820 10996 12848 11036
rect 12894 11024 12900 11076
rect 12952 11024 12958 11076
rect 13096 11064 13124 11095
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 14182 11132 14188 11144
rect 13228 11104 13273 11132
rect 14143 11104 14188 11132
rect 13228 11092 13234 11104
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 14292 11064 14320 11095
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 14424 11104 14469 11132
rect 14424 11092 14430 11104
rect 14642 11092 14648 11144
rect 14700 11092 14706 11144
rect 17126 11132 17132 11144
rect 17087 11104 17132 11132
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11101 18383 11135
rect 18325 11095 18383 11101
rect 18417 11135 18475 11141
rect 18417 11101 18429 11135
rect 18463 11132 18475 11135
rect 18463 11104 19104 11132
rect 18463 11101 18475 11104
rect 18417 11095 18475 11101
rect 14660 11064 14688 11092
rect 16574 11064 16580 11076
rect 13096 11036 14688 11064
rect 16535 11036 16580 11064
rect 16574 11024 16580 11036
rect 16632 11064 16638 11076
rect 18340 11064 18368 11095
rect 16632 11036 18368 11064
rect 18601 11067 18659 11073
rect 16632 11024 16638 11036
rect 18601 11033 18613 11067
rect 18647 11064 18659 11067
rect 19076 11064 19104 11104
rect 19150 11092 19156 11144
rect 19208 11132 19214 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 19208 11104 19257 11132
rect 19208 11092 19214 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11132 19579 11135
rect 20070 11132 20076 11144
rect 19567 11104 20076 11132
rect 19567 11101 19579 11104
rect 19521 11095 19579 11101
rect 20070 11092 20076 11104
rect 20128 11092 20134 11144
rect 25498 11092 25504 11144
rect 25556 11132 25562 11144
rect 27338 11132 27344 11144
rect 25556 11104 27344 11132
rect 25556 11092 25562 11104
rect 27338 11092 27344 11104
rect 27396 11132 27402 11144
rect 27525 11135 27583 11141
rect 27525 11132 27537 11135
rect 27396 11104 27537 11132
rect 27396 11092 27402 11104
rect 27525 11101 27537 11104
rect 27571 11101 27583 11135
rect 27525 11095 27583 11101
rect 19886 11064 19892 11076
rect 18647 11036 19012 11064
rect 19076 11036 19892 11064
rect 18647 11033 18659 11036
rect 18601 11027 18659 11033
rect 12986 10996 12992 11008
rect 12820 10968 12992 10996
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 14642 10996 14648 11008
rect 14603 10968 14648 10996
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 18984 10996 19012 11036
rect 19886 11024 19892 11036
rect 19944 11064 19950 11076
rect 20165 11067 20223 11073
rect 20165 11064 20177 11067
rect 19944 11036 20177 11064
rect 19944 11024 19950 11036
rect 20165 11033 20177 11036
rect 20211 11033 20223 11067
rect 27540 11064 27568 11095
rect 27798 11064 27804 11076
rect 27540 11036 27804 11064
rect 20165 11027 20223 11033
rect 27798 11024 27804 11036
rect 27856 11024 27862 11076
rect 19334 10996 19340 11008
rect 18984 10968 19340 10996
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 1104 10906 29600 10928
rect 1104 10854 8034 10906
rect 8086 10854 8098 10906
rect 8150 10854 8162 10906
rect 8214 10854 8226 10906
rect 8278 10854 8290 10906
rect 8342 10854 15118 10906
rect 15170 10854 15182 10906
rect 15234 10854 15246 10906
rect 15298 10854 15310 10906
rect 15362 10854 15374 10906
rect 15426 10854 22202 10906
rect 22254 10854 22266 10906
rect 22318 10854 22330 10906
rect 22382 10854 22394 10906
rect 22446 10854 22458 10906
rect 22510 10854 29286 10906
rect 29338 10854 29350 10906
rect 29402 10854 29414 10906
rect 29466 10854 29478 10906
rect 29530 10854 29542 10906
rect 29594 10854 29600 10906
rect 1104 10832 29600 10854
rect 1486 10792 1492 10804
rect 1447 10764 1492 10792
rect 1486 10752 1492 10764
rect 1544 10752 1550 10804
rect 5626 10752 5632 10804
rect 5684 10801 5690 10804
rect 5684 10795 5703 10801
rect 5691 10761 5703 10795
rect 5684 10755 5703 10761
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 5994 10792 6000 10804
rect 5859 10764 6000 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 5684 10752 5690 10755
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 10928 10764 11529 10792
rect 10928 10752 10934 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 14001 10795 14059 10801
rect 14001 10761 14013 10795
rect 14047 10792 14059 10795
rect 14182 10792 14188 10804
rect 14047 10764 14188 10792
rect 14047 10761 14059 10764
rect 14001 10755 14059 10761
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 17313 10795 17371 10801
rect 17313 10761 17325 10795
rect 17359 10792 17371 10795
rect 17402 10792 17408 10804
rect 17359 10764 17408 10792
rect 17359 10761 17371 10764
rect 17313 10755 17371 10761
rect 17402 10752 17408 10764
rect 17460 10752 17466 10804
rect 18230 10792 18236 10804
rect 18191 10764 18236 10792
rect 18230 10752 18236 10764
rect 18288 10752 18294 10804
rect 20622 10792 20628 10804
rect 20583 10764 20628 10792
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 20806 10752 20812 10804
rect 20864 10792 20870 10804
rect 21542 10792 21548 10804
rect 20864 10764 21548 10792
rect 20864 10752 20870 10764
rect 21542 10752 21548 10764
rect 21600 10752 21606 10804
rect 23382 10752 23388 10804
rect 23440 10792 23446 10804
rect 23440 10764 23612 10792
rect 23440 10752 23446 10764
rect 5442 10724 5448 10736
rect 5403 10696 5448 10724
rect 5442 10684 5448 10696
rect 5500 10684 5506 10736
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 7892 10696 8340 10724
rect 7892 10684 7898 10696
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2222 10656 2228 10668
rect 1719 10628 2228 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10656 4675 10659
rect 4890 10656 4896 10668
rect 4663 10628 4896 10656
rect 4663 10625 4675 10628
rect 4617 10619 4675 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5460 10656 5488 10684
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5460 10628 6377 10656
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 7926 10656 7932 10668
rect 7887 10628 7932 10656
rect 6365 10619 6423 10625
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8312 10665 8340 10696
rect 13464 10696 14596 10724
rect 13464 10668 13492 10696
rect 14568 10668 14596 10696
rect 17126 10684 17132 10736
rect 17184 10724 17190 10736
rect 19242 10724 19248 10736
rect 17184 10696 19248 10724
rect 17184 10684 17190 10696
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 8662 10656 8668 10668
rect 8623 10628 8668 10656
rect 8297 10619 8355 10625
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 9030 10656 9036 10668
rect 8991 10628 9036 10656
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 9490 10656 9496 10668
rect 9451 10628 9496 10656
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 12894 10616 12900 10668
rect 12952 10656 12958 10668
rect 13265 10659 13323 10665
rect 13265 10656 13277 10659
rect 12952 10628 13277 10656
rect 12952 10616 12958 10628
rect 13265 10625 13277 10628
rect 13311 10625 13323 10659
rect 13446 10656 13452 10668
rect 13359 10628 13452 10656
rect 13265 10619 13323 10625
rect 13446 10616 13452 10628
rect 13504 10616 13510 10668
rect 13630 10656 13636 10668
rect 13591 10628 13636 10656
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 14550 10656 14556 10668
rect 14511 10628 14556 10656
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 17236 10665 17264 10696
rect 17221 10659 17279 10665
rect 17221 10625 17233 10659
rect 17267 10625 17279 10659
rect 17402 10656 17408 10668
rect 17363 10628 17408 10656
rect 17221 10619 17279 10625
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 18248 10665 18276 10696
rect 19242 10684 19248 10696
rect 19300 10724 19306 10736
rect 23014 10724 23020 10736
rect 19300 10696 21496 10724
rect 19300 10684 19306 10696
rect 21468 10668 21496 10696
rect 22572 10696 23020 10724
rect 18233 10659 18291 10665
rect 18233 10625 18245 10659
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 18417 10659 18475 10665
rect 18417 10625 18429 10659
rect 18463 10656 18475 10659
rect 18463 10628 19380 10656
rect 18463 10625 18475 10628
rect 18417 10619 18475 10625
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 4525 10591 4583 10597
rect 4525 10588 4537 10591
rect 4304 10560 4537 10588
rect 4304 10548 4310 10560
rect 4525 10557 4537 10560
rect 4571 10557 4583 10591
rect 4706 10588 4712 10600
rect 4667 10560 4712 10588
rect 4525 10551 4583 10557
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 4798 10548 4804 10600
rect 4856 10588 4862 10600
rect 5350 10588 5356 10600
rect 4856 10560 5356 10588
rect 4856 10548 4862 10560
rect 5350 10548 5356 10560
rect 5408 10548 5414 10600
rect 9398 10520 9404 10532
rect 9359 10492 9404 10520
rect 9398 10480 9404 10492
rect 9456 10480 9462 10532
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 19352 10529 19380 10628
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19705 10659 19763 10665
rect 19705 10656 19717 10659
rect 19484 10628 19717 10656
rect 19484 10616 19490 10628
rect 19705 10625 19717 10628
rect 19751 10625 19763 10659
rect 21085 10659 21143 10665
rect 21085 10656 21097 10659
rect 19705 10619 19763 10625
rect 19996 10628 21097 10656
rect 19996 10600 20024 10628
rect 21085 10625 21097 10628
rect 21131 10656 21143 10659
rect 21266 10656 21272 10668
rect 21131 10628 21272 10656
rect 21131 10625 21143 10628
rect 21085 10619 21143 10625
rect 21266 10616 21272 10628
rect 21324 10616 21330 10668
rect 21450 10616 21456 10668
rect 21508 10656 21514 10668
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 21508 10628 21833 10656
rect 21508 10616 21514 10628
rect 21821 10625 21833 10628
rect 21867 10625 21879 10659
rect 21821 10619 21879 10625
rect 21910 10616 21916 10668
rect 21968 10656 21974 10668
rect 22097 10659 22155 10665
rect 21968 10628 22013 10656
rect 21968 10616 21974 10628
rect 22097 10625 22109 10659
rect 22143 10656 22155 10659
rect 22278 10656 22284 10668
rect 22143 10628 22284 10656
rect 22143 10625 22155 10628
rect 22097 10619 22155 10625
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 22572 10665 22600 10696
rect 23014 10684 23020 10696
rect 23072 10724 23078 10736
rect 23072 10696 23428 10724
rect 23072 10684 23078 10696
rect 23400 10668 23428 10696
rect 22557 10659 22615 10665
rect 22557 10625 22569 10659
rect 22603 10625 22615 10659
rect 22738 10656 22744 10668
rect 22699 10628 22744 10656
rect 22557 10619 22615 10625
rect 22738 10616 22744 10628
rect 22796 10616 22802 10668
rect 23290 10656 23296 10668
rect 23251 10628 23296 10656
rect 23290 10616 23296 10628
rect 23348 10616 23354 10668
rect 23382 10616 23388 10668
rect 23440 10656 23446 10668
rect 23477 10659 23535 10665
rect 23477 10656 23489 10659
rect 23440 10628 23489 10656
rect 23440 10616 23446 10628
rect 23477 10625 23489 10628
rect 23523 10625 23535 10659
rect 23477 10619 23535 10625
rect 19797 10591 19855 10597
rect 19797 10557 19809 10591
rect 19843 10557 19855 10591
rect 19797 10551 19855 10557
rect 19337 10523 19395 10529
rect 12032 10492 13584 10520
rect 12032 10480 12038 10492
rect 13556 10464 13584 10492
rect 19337 10489 19349 10523
rect 19383 10489 19395 10523
rect 19337 10483 19395 10489
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 2501 10455 2559 10461
rect 2501 10452 2513 10455
rect 2188 10424 2513 10452
rect 2188 10412 2194 10424
rect 2501 10421 2513 10424
rect 2547 10452 2559 10455
rect 3142 10452 3148 10464
rect 2547 10424 3148 10452
rect 2547 10421 2559 10424
rect 2501 10415 2559 10421
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 4985 10455 5043 10461
rect 4985 10452 4997 10455
rect 4948 10424 4997 10452
rect 4948 10412 4954 10424
rect 4985 10421 4997 10424
rect 5031 10452 5043 10455
rect 5629 10455 5687 10461
rect 5629 10452 5641 10455
rect 5031 10424 5641 10452
rect 5031 10421 5043 10424
rect 4985 10415 5043 10421
rect 5629 10421 5641 10424
rect 5675 10421 5687 10455
rect 5629 10415 5687 10421
rect 12805 10455 12863 10461
rect 12805 10421 12817 10455
rect 12851 10452 12863 10455
rect 12894 10452 12900 10464
rect 12851 10424 12900 10452
rect 12851 10421 12863 10424
rect 12805 10415 12863 10421
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 13538 10452 13544 10464
rect 13499 10424 13544 10452
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 13722 10452 13728 10464
rect 13683 10424 13728 10452
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 19812 10452 19840 10551
rect 19978 10548 19984 10600
rect 20036 10588 20042 10600
rect 20714 10588 20720 10600
rect 20036 10560 20129 10588
rect 20675 10560 20720 10588
rect 20036 10548 20042 10560
rect 20714 10548 20720 10560
rect 20772 10548 20778 10600
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10588 20867 10591
rect 21468 10588 21496 10616
rect 20855 10560 21496 10588
rect 23201 10591 23259 10597
rect 20855 10557 20867 10560
rect 20809 10551 20867 10557
rect 23201 10557 23213 10591
rect 23247 10588 23259 10591
rect 23584 10588 23612 10764
rect 25130 10752 25136 10804
rect 25188 10792 25194 10804
rect 25593 10795 25651 10801
rect 25593 10792 25605 10795
rect 25188 10764 25605 10792
rect 25188 10752 25194 10764
rect 25593 10761 25605 10764
rect 25639 10761 25651 10795
rect 25593 10755 25651 10761
rect 27617 10795 27675 10801
rect 27617 10761 27629 10795
rect 27663 10792 27675 10795
rect 27706 10792 27712 10804
rect 27663 10764 27712 10792
rect 27663 10761 27675 10764
rect 27617 10755 27675 10761
rect 27706 10752 27712 10764
rect 27764 10752 27770 10804
rect 23661 10727 23719 10733
rect 23661 10693 23673 10727
rect 23707 10724 23719 10727
rect 28258 10724 28264 10736
rect 23707 10696 25084 10724
rect 23707 10693 23719 10696
rect 23661 10687 23719 10693
rect 23842 10616 23848 10668
rect 23900 10656 23906 10668
rect 24121 10659 24179 10665
rect 24121 10656 24133 10659
rect 23900 10628 24133 10656
rect 23900 10616 23906 10628
rect 24121 10625 24133 10628
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 24305 10659 24363 10665
rect 24305 10625 24317 10659
rect 24351 10625 24363 10659
rect 24854 10656 24860 10668
rect 24815 10628 24860 10656
rect 24305 10619 24363 10625
rect 23247 10560 23612 10588
rect 23247 10557 23259 10560
rect 23201 10551 23259 10557
rect 23308 10532 23336 10560
rect 20346 10480 20352 10532
rect 20404 10520 20410 10532
rect 21821 10523 21879 10529
rect 21821 10520 21833 10523
rect 20404 10492 21833 10520
rect 20404 10480 20410 10492
rect 21821 10489 21833 10492
rect 21867 10489 21879 10523
rect 21821 10483 21879 10489
rect 23290 10480 23296 10532
rect 23348 10480 23354 10532
rect 24210 10520 24216 10532
rect 24171 10492 24216 10520
rect 24210 10480 24216 10492
rect 24268 10480 24274 10532
rect 24320 10520 24348 10619
rect 24854 10616 24860 10628
rect 24912 10616 24918 10668
rect 25056 10665 25084 10696
rect 25424 10696 28264 10724
rect 25041 10659 25099 10665
rect 25041 10625 25053 10659
rect 25087 10625 25099 10659
rect 25041 10619 25099 10625
rect 25314 10616 25320 10668
rect 25372 10656 25378 10668
rect 25424 10665 25452 10696
rect 28258 10684 28264 10696
rect 28316 10684 28322 10736
rect 25409 10659 25467 10665
rect 25409 10656 25421 10659
rect 25372 10628 25421 10656
rect 25372 10616 25378 10628
rect 25409 10625 25421 10628
rect 25455 10625 25467 10659
rect 25409 10619 25467 10625
rect 25682 10616 25688 10668
rect 25740 10656 25746 10668
rect 26973 10659 27031 10665
rect 26973 10656 26985 10659
rect 25740 10628 26985 10656
rect 25740 10616 25746 10628
rect 26973 10625 26985 10628
rect 27019 10625 27031 10659
rect 27154 10656 27160 10668
rect 27115 10628 27160 10656
rect 26973 10619 27031 10625
rect 27154 10616 27160 10628
rect 27212 10656 27218 10668
rect 27212 10628 27660 10656
rect 27212 10616 27218 10628
rect 24872 10588 24900 10616
rect 25130 10588 25136 10600
rect 24872 10560 24992 10588
rect 25091 10560 25136 10588
rect 24854 10520 24860 10532
rect 24320 10492 24860 10520
rect 24854 10480 24860 10492
rect 24912 10480 24918 10532
rect 24964 10520 24992 10560
rect 25130 10548 25136 10560
rect 25188 10548 25194 10600
rect 27632 10597 27660 10628
rect 27798 10616 27804 10668
rect 27856 10656 27862 10668
rect 27893 10659 27951 10665
rect 27893 10656 27905 10659
rect 27856 10628 27905 10656
rect 27856 10616 27862 10628
rect 27893 10625 27905 10628
rect 27939 10625 27951 10659
rect 27893 10619 27951 10625
rect 25225 10591 25283 10597
rect 25225 10557 25237 10591
rect 25271 10588 25283 10591
rect 27617 10591 27675 10597
rect 25271 10560 25728 10588
rect 25271 10557 25283 10560
rect 25225 10551 25283 10557
rect 25590 10520 25596 10532
rect 24964 10492 25596 10520
rect 25590 10480 25596 10492
rect 25648 10480 25654 10532
rect 25700 10520 25728 10560
rect 27617 10557 27629 10591
rect 27663 10557 27675 10591
rect 27617 10551 27675 10557
rect 27065 10523 27123 10529
rect 27065 10520 27077 10523
rect 25700 10492 27077 10520
rect 27065 10489 27077 10492
rect 27111 10520 27123 10523
rect 28166 10520 28172 10532
rect 27111 10492 28172 10520
rect 27111 10489 27123 10492
rect 27065 10483 27123 10489
rect 28166 10480 28172 10492
rect 28224 10480 28230 10532
rect 20806 10452 20812 10464
rect 19812 10424 20812 10452
rect 20806 10412 20812 10424
rect 20864 10412 20870 10464
rect 20898 10412 20904 10464
rect 20956 10452 20962 10464
rect 20993 10455 21051 10461
rect 20993 10452 21005 10455
rect 20956 10424 21005 10452
rect 20956 10412 20962 10424
rect 20993 10421 21005 10424
rect 21039 10421 21051 10455
rect 22554 10452 22560 10464
rect 22515 10424 22560 10452
rect 20993 10415 21051 10421
rect 22554 10412 22560 10424
rect 22612 10412 22618 10464
rect 22738 10412 22744 10464
rect 22796 10452 22802 10464
rect 25682 10452 25688 10464
rect 22796 10424 25688 10452
rect 22796 10412 22802 10424
rect 25682 10412 25688 10424
rect 25740 10412 25746 10464
rect 27798 10412 27804 10464
rect 27856 10452 27862 10464
rect 27856 10424 27901 10452
rect 27856 10412 27862 10424
rect 1104 10362 29440 10384
rect 1104 10310 4492 10362
rect 4544 10310 4556 10362
rect 4608 10310 4620 10362
rect 4672 10310 4684 10362
rect 4736 10310 4748 10362
rect 4800 10310 11576 10362
rect 11628 10310 11640 10362
rect 11692 10310 11704 10362
rect 11756 10310 11768 10362
rect 11820 10310 11832 10362
rect 11884 10310 18660 10362
rect 18712 10310 18724 10362
rect 18776 10310 18788 10362
rect 18840 10310 18852 10362
rect 18904 10310 18916 10362
rect 18968 10310 25744 10362
rect 25796 10310 25808 10362
rect 25860 10310 25872 10362
rect 25924 10310 25936 10362
rect 25988 10310 26000 10362
rect 26052 10310 29440 10362
rect 1104 10288 29440 10310
rect 9033 10251 9091 10257
rect 9033 10217 9045 10251
rect 9079 10248 9091 10251
rect 9490 10248 9496 10260
rect 9079 10220 9496 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 12710 10248 12716 10260
rect 9600 10220 12716 10248
rect 9600 10180 9628 10220
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 12989 10251 13047 10257
rect 12989 10217 13001 10251
rect 13035 10248 13047 10251
rect 13170 10248 13176 10260
rect 13035 10220 13176 10248
rect 13035 10217 13047 10220
rect 12989 10211 13047 10217
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 17310 10208 17316 10260
rect 17368 10248 17374 10260
rect 17405 10251 17463 10257
rect 17405 10248 17417 10251
rect 17368 10220 17417 10248
rect 17368 10208 17374 10220
rect 17405 10217 17417 10220
rect 17451 10217 17463 10251
rect 19978 10248 19984 10260
rect 19939 10220 19984 10248
rect 17405 10211 17463 10217
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 20714 10208 20720 10260
rect 20772 10248 20778 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20772 10220 20913 10248
rect 20772 10208 20778 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 4816 10152 9628 10180
rect 10965 10183 11023 10189
rect 4816 10121 4844 10152
rect 10965 10149 10977 10183
rect 11011 10180 11023 10183
rect 13722 10180 13728 10192
rect 11011 10152 13728 10180
rect 11011 10149 11023 10152
rect 10965 10143 11023 10149
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 17880 10152 20852 10180
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10081 4859 10115
rect 7650 10112 7656 10124
rect 7611 10084 7656 10112
rect 4801 10075 4859 10081
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 10336 10084 11437 10112
rect 10336 10056 10364 10084
rect 11425 10081 11437 10084
rect 11471 10112 11483 10115
rect 13814 10112 13820 10124
rect 11471 10084 13820 10112
rect 11471 10081 11483 10084
rect 11425 10075 11483 10081
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4212 10016 4537 10044
rect 4212 10004 4218 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10044 7619 10047
rect 8386 10044 8392 10056
rect 7607 10016 8392 10044
rect 7607 10013 7619 10016
rect 7561 10007 7619 10013
rect 8386 10004 8392 10016
rect 8444 10044 8450 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8444 10016 8953 10044
rect 8444 10004 8450 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 8941 10007 8999 10013
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10502 10044 10508 10056
rect 10463 10016 10508 10044
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 10778 10044 10784 10056
rect 10739 10016 10784 10044
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 12342 10044 12348 10056
rect 12303 10016 12348 10044
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12810 10047 12868 10053
rect 12492 10016 12537 10044
rect 12492 10004 12498 10016
rect 12810 10013 12822 10047
rect 12856 10044 12868 10047
rect 12986 10044 12992 10056
rect 12856 10016 12992 10044
rect 12856 10013 12868 10016
rect 12810 10007 12868 10013
rect 12986 10004 12992 10016
rect 13044 10044 13050 10056
rect 14645 10047 14703 10053
rect 14645 10044 14657 10047
rect 13044 10016 14657 10044
rect 13044 10004 13050 10016
rect 14645 10013 14657 10016
rect 14691 10044 14703 10047
rect 15746 10044 15752 10056
rect 14691 10016 15752 10044
rect 14691 10013 14703 10016
rect 14645 10007 14703 10013
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 16758 10004 16764 10056
rect 16816 10044 16822 10056
rect 17880 10053 17908 10152
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10112 18107 10115
rect 18095 10084 18736 10112
rect 18095 10081 18107 10084
rect 18049 10075 18107 10081
rect 17865 10047 17923 10053
rect 17865 10044 17877 10047
rect 16816 10016 17877 10044
rect 16816 10004 16822 10016
rect 17865 10013 17877 10016
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 12250 9936 12256 9988
rect 12308 9976 12314 9988
rect 12621 9979 12679 9985
rect 12621 9976 12633 9979
rect 12308 9948 12633 9976
rect 12308 9936 12314 9948
rect 12621 9945 12633 9948
rect 12667 9945 12679 9979
rect 12621 9939 12679 9945
rect 12713 9979 12771 9985
rect 12713 9945 12725 9979
rect 12759 9945 12771 9979
rect 12713 9939 12771 9945
rect 2406 9868 2412 9920
rect 2464 9908 2470 9920
rect 2593 9911 2651 9917
rect 2593 9908 2605 9911
rect 2464 9880 2605 9908
rect 2464 9868 2470 9880
rect 2593 9877 2605 9880
rect 2639 9877 2651 9911
rect 7926 9908 7932 9920
rect 7887 9880 7932 9908
rect 2593 9871 2651 9877
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 12728 9908 12756 9939
rect 13078 9936 13084 9988
rect 13136 9976 13142 9988
rect 13538 9976 13544 9988
rect 13136 9948 13544 9976
rect 13136 9936 13142 9948
rect 13538 9936 13544 9948
rect 13596 9976 13602 9988
rect 14093 9979 14151 9985
rect 14093 9976 14105 9979
rect 13596 9948 14105 9976
rect 13596 9936 13602 9948
rect 14093 9945 14105 9948
rect 14139 9945 14151 9979
rect 14093 9939 14151 9945
rect 16393 9979 16451 9985
rect 16393 9945 16405 9979
rect 16439 9976 16451 9979
rect 16439 9948 17816 9976
rect 16439 9945 16451 9948
rect 16393 9939 16451 9945
rect 17788 9920 17816 9948
rect 18708 9920 18736 10084
rect 19334 10044 19340 10056
rect 19295 10016 19340 10044
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10044 20591 10047
rect 20622 10044 20628 10056
rect 20579 10016 20628 10044
rect 20579 10013 20591 10016
rect 20533 10007 20591 10013
rect 20622 10004 20628 10016
rect 20680 10004 20686 10056
rect 20714 9976 20720 9988
rect 20675 9948 20720 9976
rect 20714 9936 20720 9948
rect 20772 9936 20778 9988
rect 20824 9976 20852 10152
rect 20916 10044 20944 10211
rect 21910 10208 21916 10260
rect 21968 10248 21974 10260
rect 22278 10248 22284 10260
rect 21968 10220 22094 10248
rect 22239 10220 22284 10248
rect 21968 10208 21974 10220
rect 22066 10180 22094 10220
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 23382 10208 23388 10260
rect 23440 10248 23446 10260
rect 24397 10251 24455 10257
rect 24397 10248 24409 10251
rect 23440 10220 24409 10248
rect 23440 10208 23446 10220
rect 24397 10217 24409 10220
rect 24443 10217 24455 10251
rect 24397 10211 24455 10217
rect 25130 10208 25136 10260
rect 25188 10248 25194 10260
rect 25317 10251 25375 10257
rect 25317 10248 25329 10251
rect 25188 10220 25329 10248
rect 25188 10208 25194 10220
rect 25317 10217 25329 10220
rect 25363 10217 25375 10251
rect 25317 10211 25375 10217
rect 23201 10183 23259 10189
rect 23201 10180 23213 10183
rect 22066 10152 23213 10180
rect 23201 10149 23213 10152
rect 23247 10180 23259 10183
rect 25409 10183 25467 10189
rect 25409 10180 25421 10183
rect 23247 10152 25421 10180
rect 23247 10149 23259 10152
rect 23201 10143 23259 10149
rect 25409 10149 25421 10152
rect 25455 10149 25467 10183
rect 25409 10143 25467 10149
rect 21821 10115 21879 10121
rect 21821 10081 21833 10115
rect 21867 10112 21879 10115
rect 22738 10112 22744 10124
rect 21867 10084 22744 10112
rect 21867 10081 21879 10084
rect 21821 10075 21879 10081
rect 22738 10072 22744 10084
rect 22796 10072 22802 10124
rect 23106 10072 23112 10124
rect 23164 10112 23170 10124
rect 25225 10115 25283 10121
rect 23164 10084 24440 10112
rect 23164 10072 23170 10084
rect 21361 10047 21419 10053
rect 21361 10044 21373 10047
rect 20916 10016 21373 10044
rect 21361 10013 21373 10016
rect 21407 10013 21419 10047
rect 21634 10044 21640 10056
rect 21595 10016 21640 10044
rect 21361 10007 21419 10013
rect 21634 10004 21640 10016
rect 21692 10004 21698 10056
rect 24412 10053 24440 10084
rect 25225 10081 25237 10115
rect 25271 10112 25283 10115
rect 25314 10112 25320 10124
rect 25271 10084 25320 10112
rect 25271 10081 25283 10084
rect 25225 10075 25283 10081
rect 25314 10072 25320 10084
rect 25372 10072 25378 10124
rect 25590 10072 25596 10124
rect 25648 10112 25654 10124
rect 27065 10115 27123 10121
rect 27065 10112 27077 10115
rect 25648 10084 27077 10112
rect 25648 10072 25654 10084
rect 27065 10081 27077 10084
rect 27111 10081 27123 10115
rect 28166 10112 28172 10124
rect 28127 10084 28172 10112
rect 27065 10075 27123 10081
rect 28166 10072 28172 10084
rect 28224 10072 28230 10124
rect 28258 10072 28264 10124
rect 28316 10112 28322 10124
rect 28316 10084 28361 10112
rect 28316 10072 28322 10084
rect 23569 10047 23627 10053
rect 23569 10044 23581 10047
rect 22388 10016 23581 10044
rect 20898 9976 20904 9988
rect 20824 9948 20904 9976
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 21453 9979 21511 9985
rect 21453 9945 21465 9979
rect 21499 9976 21511 9979
rect 22186 9976 22192 9988
rect 21499 9948 22192 9976
rect 21499 9945 21511 9948
rect 21453 9939 21511 9945
rect 22186 9936 22192 9948
rect 22244 9936 22250 9988
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 12728 9880 13461 9908
rect 13449 9877 13461 9880
rect 13495 9908 13507 9911
rect 13906 9908 13912 9920
rect 13495 9880 13912 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 16853 9911 16911 9917
rect 16853 9908 16865 9911
rect 16816 9880 16865 9908
rect 16816 9868 16822 9880
rect 16853 9877 16865 9880
rect 16899 9877 16911 9911
rect 17770 9908 17776 9920
rect 17731 9880 17776 9908
rect 16853 9871 16911 9877
rect 17770 9868 17776 9880
rect 17828 9868 17834 9920
rect 18690 9908 18696 9920
rect 18651 9880 18696 9908
rect 18690 9868 18696 9880
rect 18748 9868 18754 9920
rect 19426 9868 19432 9920
rect 19484 9908 19490 9920
rect 22388 9908 22416 10016
rect 23569 10013 23581 10016
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 24397 10047 24455 10053
rect 24397 10013 24409 10047
rect 24443 10013 24455 10047
rect 24397 10007 24455 10013
rect 24489 10047 24547 10053
rect 24489 10013 24501 10047
rect 24535 10013 24547 10047
rect 25498 10044 25504 10056
rect 25459 10016 25504 10044
rect 24489 10007 24547 10013
rect 22465 9979 22523 9985
rect 22465 9945 22477 9979
rect 22511 9945 22523 9979
rect 22465 9939 22523 9945
rect 22649 9979 22707 9985
rect 22649 9945 22661 9979
rect 22695 9976 22707 9979
rect 22738 9976 22744 9988
rect 22695 9948 22744 9976
rect 22695 9945 22707 9948
rect 22649 9939 22707 9945
rect 19484 9880 22416 9908
rect 22480 9908 22508 9939
rect 22738 9936 22744 9948
rect 22796 9936 22802 9988
rect 23290 9936 23296 9988
rect 23348 9976 23354 9988
rect 23385 9979 23443 9985
rect 23385 9976 23397 9979
rect 23348 9948 23397 9976
rect 23348 9936 23354 9948
rect 23385 9945 23397 9948
rect 23431 9976 23443 9979
rect 24504 9976 24532 10007
rect 25498 10004 25504 10016
rect 25556 10004 25562 10056
rect 26878 10044 26884 10056
rect 26839 10016 26884 10044
rect 26878 10004 26884 10016
rect 26936 10004 26942 10056
rect 27706 10004 27712 10056
rect 27764 10044 27770 10056
rect 28077 10047 28135 10053
rect 28077 10044 28089 10047
rect 27764 10016 28089 10044
rect 27764 10004 27770 10016
rect 28077 10013 28089 10016
rect 28123 10013 28135 10047
rect 28077 10007 28135 10013
rect 25961 9979 26019 9985
rect 25961 9976 25973 9979
rect 23431 9948 25973 9976
rect 23431 9945 23443 9948
rect 23385 9939 23443 9945
rect 25961 9945 25973 9948
rect 26007 9945 26019 9979
rect 25961 9939 26019 9945
rect 27614 9936 27620 9988
rect 27672 9976 27678 9988
rect 28276 9976 28304 10072
rect 27672 9948 28304 9976
rect 27672 9936 27678 9948
rect 22922 9908 22928 9920
rect 22480 9880 22928 9908
rect 19484 9868 19490 9880
rect 22922 9868 22928 9880
rect 22980 9868 22986 9920
rect 24765 9911 24823 9917
rect 24765 9877 24777 9911
rect 24811 9908 24823 9911
rect 25406 9908 25412 9920
rect 24811 9880 25412 9908
rect 24811 9877 24823 9880
rect 24765 9871 24823 9877
rect 25406 9868 25412 9880
rect 25464 9868 25470 9920
rect 26510 9908 26516 9920
rect 26471 9880 26516 9908
rect 26510 9868 26516 9880
rect 26568 9868 26574 9920
rect 26973 9911 27031 9917
rect 26973 9877 26985 9911
rect 27019 9908 27031 9911
rect 27709 9911 27767 9917
rect 27709 9908 27721 9911
rect 27019 9880 27721 9908
rect 27019 9877 27031 9880
rect 26973 9871 27031 9877
rect 27709 9877 27721 9880
rect 27755 9877 27767 9911
rect 27709 9871 27767 9877
rect 1104 9818 29600 9840
rect 1104 9766 8034 9818
rect 8086 9766 8098 9818
rect 8150 9766 8162 9818
rect 8214 9766 8226 9818
rect 8278 9766 8290 9818
rect 8342 9766 15118 9818
rect 15170 9766 15182 9818
rect 15234 9766 15246 9818
rect 15298 9766 15310 9818
rect 15362 9766 15374 9818
rect 15426 9766 22202 9818
rect 22254 9766 22266 9818
rect 22318 9766 22330 9818
rect 22382 9766 22394 9818
rect 22446 9766 22458 9818
rect 22510 9766 29286 9818
rect 29338 9766 29350 9818
rect 29402 9766 29414 9818
rect 29466 9766 29478 9818
rect 29530 9766 29542 9818
rect 29594 9766 29600 9818
rect 1104 9744 29600 9766
rect 9232 9676 9812 9704
rect 9232 9648 9260 9676
rect 2133 9639 2191 9645
rect 2133 9605 2145 9639
rect 2179 9636 2191 9639
rect 2222 9636 2228 9648
rect 2179 9608 2228 9636
rect 2179 9605 2191 9608
rect 2133 9599 2191 9605
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 3142 9636 3148 9648
rect 3055 9608 3148 9636
rect 3142 9596 3148 9608
rect 3200 9636 3206 9648
rect 3878 9636 3884 9648
rect 3200 9608 3884 9636
rect 3200 9596 3206 9608
rect 3878 9596 3884 9608
rect 3936 9636 3942 9648
rect 7282 9636 7288 9648
rect 3936 9608 7288 9636
rect 3936 9596 3942 9608
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 8021 9639 8079 9645
rect 8021 9605 8033 9639
rect 8067 9636 8079 9639
rect 8294 9636 8300 9648
rect 8067 9608 8300 9636
rect 8067 9605 8079 9608
rect 8021 9599 8079 9605
rect 8294 9596 8300 9608
rect 8352 9636 8358 9648
rect 8570 9636 8576 9648
rect 8352 9608 8576 9636
rect 8352 9596 8358 9608
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 9214 9636 9220 9648
rect 9127 9608 9220 9636
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9568 2375 9571
rect 2406 9568 2412 9580
rect 2363 9540 2412 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 2406 9528 2412 9540
rect 2464 9528 2470 9580
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 4338 9568 4344 9580
rect 3384 9540 3924 9568
rect 4299 9540 4344 9568
rect 3384 9528 3390 9540
rect 3896 9441 3924 9540
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 7064 9540 7113 9568
rect 7064 9528 7070 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7926 9568 7932 9580
rect 7887 9540 7932 9568
rect 7101 9531 7159 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 8220 9500 8248 9531
rect 8386 9528 8392 9580
rect 8444 9568 8450 9580
rect 9140 9577 9168 9608
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 9674 9636 9680 9648
rect 9324 9608 9680 9636
rect 9324 9577 9352 9608
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 9784 9636 9812 9676
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 10965 9707 11023 9713
rect 10965 9704 10977 9707
rect 10560 9676 10977 9704
rect 10560 9664 10566 9676
rect 10965 9673 10977 9676
rect 11011 9673 11023 9707
rect 12342 9704 12348 9716
rect 12303 9676 12348 9704
rect 10965 9667 11023 9673
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 17402 9704 17408 9716
rect 17363 9676 17408 9704
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 21821 9707 21879 9713
rect 21821 9704 21833 9707
rect 20772 9676 21833 9704
rect 20772 9664 20778 9676
rect 21821 9673 21833 9676
rect 21867 9704 21879 9707
rect 22462 9704 22468 9716
rect 21867 9676 22468 9704
rect 21867 9673 21879 9676
rect 21821 9667 21879 9673
rect 22462 9664 22468 9676
rect 22520 9664 22526 9716
rect 22922 9704 22928 9716
rect 22883 9676 22928 9704
rect 22922 9664 22928 9676
rect 22980 9664 22986 9716
rect 27798 9704 27804 9716
rect 27759 9676 27804 9704
rect 27798 9664 27804 9676
rect 27856 9664 27862 9716
rect 13722 9636 13728 9648
rect 9784 9608 10364 9636
rect 9033 9571 9091 9577
rect 9033 9568 9045 9571
rect 8444 9540 9045 9568
rect 8444 9528 8450 9540
rect 9033 9537 9045 9540
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 10336 9509 10364 9608
rect 12406 9608 13728 9636
rect 10597 9571 10655 9577
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 10962 9568 10968 9580
rect 10643 9540 10968 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 10962 9528 10968 9540
rect 11020 9568 11026 9580
rect 12406 9568 12434 9608
rect 13722 9596 13728 9608
rect 13780 9636 13786 9648
rect 14369 9639 14427 9645
rect 14369 9636 14381 9639
rect 13780 9608 14381 9636
rect 13780 9596 13786 9608
rect 14369 9605 14381 9608
rect 14415 9605 14427 9639
rect 15841 9639 15899 9645
rect 15841 9636 15853 9639
rect 14369 9599 14427 9605
rect 15120 9608 15853 9636
rect 11020 9540 12434 9568
rect 11020 9528 11026 9540
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12860 9540 12909 9568
rect 12860 9528 12866 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 14918 9568 14924 9580
rect 14148 9540 14924 9568
rect 14148 9528 14154 9540
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 15120 9577 15148 9608
rect 15841 9605 15853 9608
rect 15887 9636 15899 9639
rect 17586 9636 17592 9648
rect 15887 9608 17592 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 17586 9596 17592 9608
rect 17644 9596 17650 9648
rect 17865 9639 17923 9645
rect 17865 9636 17877 9639
rect 17696 9608 17877 9636
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9537 15163 9571
rect 15286 9568 15292 9580
rect 15247 9540 15292 9568
rect 15105 9531 15163 9537
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 17034 9528 17040 9580
rect 17092 9568 17098 9580
rect 17696 9568 17724 9608
rect 17865 9605 17877 9608
rect 17911 9605 17923 9639
rect 18690 9636 18696 9648
rect 17865 9599 17923 9605
rect 18064 9608 18696 9636
rect 17092 9540 17724 9568
rect 17773 9571 17831 9577
rect 17092 9528 17098 9540
rect 17773 9537 17785 9571
rect 17819 9537 17831 9571
rect 17773 9531 17831 9537
rect 10321 9503 10379 9509
rect 8220 9472 10272 9500
rect 3881 9435 3939 9441
rect 3881 9401 3893 9435
rect 3927 9432 3939 9435
rect 7926 9432 7932 9444
rect 3927 9404 7932 9432
rect 3927 9401 3939 9404
rect 3881 9395 3939 9401
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 10244 9432 10272 9472
rect 10321 9469 10333 9503
rect 10367 9469 10379 9503
rect 10321 9463 10379 9469
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9500 10563 9503
rect 11054 9500 11060 9512
rect 10551 9472 11060 9500
rect 10551 9469 10563 9472
rect 10505 9463 10563 9469
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 12250 9460 12256 9512
rect 12308 9500 12314 9512
rect 12526 9500 12532 9512
rect 12308 9472 12532 9500
rect 12308 9460 12314 9472
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9500 12679 9503
rect 13078 9500 13084 9512
rect 12667 9472 13084 9500
rect 12667 9469 12679 9472
rect 12621 9463 12679 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14550 9500 14556 9512
rect 13964 9472 14556 9500
rect 13964 9460 13970 9472
rect 14550 9460 14556 9472
rect 14608 9500 14614 9512
rect 17788 9500 17816 9531
rect 18064 9509 18092 9608
rect 18690 9596 18696 9608
rect 18748 9636 18754 9648
rect 19610 9636 19616 9648
rect 18748 9608 19616 9636
rect 18748 9596 18754 9608
rect 19610 9596 19616 9608
rect 19668 9636 19674 9648
rect 22940 9636 22968 9664
rect 19668 9608 22968 9636
rect 19668 9596 19674 9608
rect 23290 9596 23296 9648
rect 23348 9636 23354 9648
rect 23661 9639 23719 9645
rect 23661 9636 23673 9639
rect 23348 9608 23673 9636
rect 23348 9596 23354 9608
rect 23661 9605 23673 9608
rect 23707 9636 23719 9639
rect 24305 9639 24363 9645
rect 24305 9636 24317 9639
rect 23707 9608 24317 9636
rect 23707 9605 23719 9608
rect 23661 9599 23719 9605
rect 24305 9605 24317 9608
rect 24351 9605 24363 9639
rect 24946 9636 24952 9648
rect 24907 9608 24952 9636
rect 24305 9599 24363 9605
rect 24946 9596 24952 9608
rect 25004 9596 25010 9648
rect 25130 9596 25136 9648
rect 25188 9636 25194 9648
rect 25188 9608 25360 9636
rect 25188 9596 25194 9608
rect 20441 9571 20499 9577
rect 20441 9537 20453 9571
rect 20487 9568 20499 9571
rect 20806 9568 20812 9580
rect 20487 9540 20812 9568
rect 20487 9537 20499 9540
rect 20441 9531 20499 9537
rect 20806 9528 20812 9540
rect 20864 9528 20870 9580
rect 20898 9528 20904 9580
rect 20956 9568 20962 9580
rect 20956 9540 21001 9568
rect 20956 9528 20962 9540
rect 22462 9528 22468 9580
rect 22520 9568 22526 9580
rect 23308 9568 23336 9596
rect 23842 9568 23848 9580
rect 22520 9540 23336 9568
rect 23803 9540 23848 9568
rect 22520 9528 22526 9540
rect 23842 9528 23848 9540
rect 23900 9528 23906 9580
rect 25222 9568 25228 9580
rect 25183 9540 25228 9568
rect 25222 9528 25228 9540
rect 25280 9528 25286 9580
rect 25332 9577 25360 9608
rect 25317 9571 25375 9577
rect 25317 9537 25329 9571
rect 25363 9537 25375 9571
rect 25317 9531 25375 9537
rect 25406 9528 25412 9580
rect 25464 9568 25470 9580
rect 25590 9568 25596 9580
rect 25464 9540 25509 9568
rect 25551 9540 25596 9568
rect 25464 9528 25470 9540
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 27617 9571 27675 9577
rect 27617 9568 27629 9571
rect 25700 9540 27629 9568
rect 14608 9472 17816 9500
rect 14608 9460 14614 9472
rect 14642 9432 14648 9444
rect 10244 9404 14648 9432
rect 14642 9392 14648 9404
rect 14700 9392 14706 9444
rect 2498 9364 2504 9376
rect 2459 9336 2504 9364
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 2958 9364 2964 9376
rect 2919 9336 2964 9364
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 4338 9324 4344 9376
rect 4396 9364 4402 9376
rect 4433 9367 4491 9373
rect 4433 9364 4445 9367
rect 4396 9336 4445 9364
rect 4396 9324 4402 9336
rect 4433 9333 4445 9336
rect 4479 9333 4491 9367
rect 4433 9327 4491 9333
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 7616 9336 8401 9364
rect 7616 9324 7622 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 8389 9327 8447 9333
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 11020 9336 11529 9364
rect 11020 9324 11026 9336
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 12526 9364 12532 9376
rect 12487 9336 12532 9364
rect 11517 9327 11575 9333
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 12618 9324 12624 9376
rect 12676 9364 12682 9376
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 12676 9336 13461 9364
rect 12676 9324 12682 9336
rect 13449 9333 13461 9336
rect 13495 9364 13507 9367
rect 14182 9364 14188 9376
rect 13495 9336 14188 9364
rect 13495 9333 13507 9336
rect 13449 9327 13507 9333
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 14918 9324 14924 9376
rect 14976 9364 14982 9376
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 14976 9336 15301 9364
rect 14976 9324 14982 9336
rect 15289 9333 15301 9336
rect 15335 9333 15347 9367
rect 15289 9327 15347 9333
rect 16945 9367 17003 9373
rect 16945 9333 16957 9367
rect 16991 9364 17003 9367
rect 17034 9364 17040 9376
rect 16991 9336 17040 9364
rect 16991 9333 17003 9336
rect 16945 9327 17003 9333
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 17788 9364 17816 9472
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9469 18107 9503
rect 23474 9500 23480 9512
rect 23387 9472 23480 9500
rect 18049 9463 18107 9469
rect 23474 9460 23480 9472
rect 23532 9500 23538 9512
rect 25700 9500 25728 9540
rect 27617 9537 27629 9540
rect 27663 9537 27675 9571
rect 28718 9568 28724 9580
rect 28679 9540 28724 9568
rect 27617 9531 27675 9537
rect 28718 9528 28724 9540
rect 28776 9528 28782 9580
rect 23532 9472 25728 9500
rect 27341 9503 27399 9509
rect 23532 9460 23538 9472
rect 27341 9469 27353 9503
rect 27387 9500 27399 9503
rect 28074 9500 28080 9512
rect 27387 9472 28080 9500
rect 27387 9469 27399 9472
rect 27341 9463 27399 9469
rect 28074 9460 28080 9472
rect 28132 9460 28138 9512
rect 27433 9435 27491 9441
rect 27433 9432 27445 9435
rect 22066 9404 27445 9432
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 17788 9336 19257 9364
rect 19245 9333 19257 9336
rect 19291 9364 19303 9367
rect 20622 9364 20628 9376
rect 19291 9336 20628 9364
rect 19291 9333 19303 9336
rect 19245 9327 19303 9333
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 20898 9324 20904 9376
rect 20956 9364 20962 9376
rect 22066 9364 22094 9404
rect 27433 9401 27445 9404
rect 27479 9432 27491 9435
rect 27614 9432 27620 9444
rect 27479 9404 27620 9432
rect 27479 9401 27491 9404
rect 27433 9395 27491 9401
rect 27614 9392 27620 9404
rect 27672 9392 27678 9444
rect 28810 9432 28816 9444
rect 27724 9404 28816 9432
rect 20956 9336 22094 9364
rect 22465 9367 22523 9373
rect 20956 9324 20962 9336
rect 22465 9333 22477 9367
rect 22511 9364 22523 9367
rect 22738 9364 22744 9376
rect 22511 9336 22744 9364
rect 22511 9333 22523 9336
rect 22465 9327 22523 9333
rect 22738 9324 22744 9336
rect 22796 9364 22802 9376
rect 22922 9364 22928 9376
rect 22796 9336 22928 9364
rect 22796 9324 22802 9336
rect 22922 9324 22928 9336
rect 22980 9324 22986 9376
rect 23658 9324 23664 9376
rect 23716 9364 23722 9376
rect 27724 9364 27752 9404
rect 28810 9392 28816 9404
rect 28868 9392 28874 9444
rect 28534 9364 28540 9376
rect 23716 9336 27752 9364
rect 28495 9336 28540 9364
rect 23716 9324 23722 9336
rect 28534 9324 28540 9336
rect 28592 9324 28598 9376
rect 1104 9274 29440 9296
rect 1104 9222 4492 9274
rect 4544 9222 4556 9274
rect 4608 9222 4620 9274
rect 4672 9222 4684 9274
rect 4736 9222 4748 9274
rect 4800 9222 11576 9274
rect 11628 9222 11640 9274
rect 11692 9222 11704 9274
rect 11756 9222 11768 9274
rect 11820 9222 11832 9274
rect 11884 9222 18660 9274
rect 18712 9222 18724 9274
rect 18776 9222 18788 9274
rect 18840 9222 18852 9274
rect 18904 9222 18916 9274
rect 18968 9222 25744 9274
rect 25796 9222 25808 9274
rect 25860 9222 25872 9274
rect 25924 9222 25936 9274
rect 25988 9222 26000 9274
rect 26052 9222 29440 9274
rect 1104 9200 29440 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2314 9160 2320 9172
rect 1995 9132 2320 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 3878 9160 3884 9172
rect 3839 9132 3884 9160
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 4801 9163 4859 9169
rect 4801 9129 4813 9163
rect 4847 9160 4859 9163
rect 5074 9160 5080 9172
rect 4847 9132 5080 9160
rect 4847 9129 4859 9132
rect 4801 9123 4859 9129
rect 5074 9120 5080 9132
rect 5132 9160 5138 9172
rect 5537 9163 5595 9169
rect 5537 9160 5549 9163
rect 5132 9132 5549 9160
rect 5132 9120 5138 9132
rect 5537 9129 5549 9132
rect 5583 9129 5595 9163
rect 7006 9160 7012 9172
rect 6967 9132 7012 9160
rect 5537 9123 5595 9129
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 8294 9160 8300 9172
rect 8255 9132 8300 9160
rect 8294 9120 8300 9132
rect 8352 9160 8358 9172
rect 8754 9160 8760 9172
rect 8352 9132 8760 9160
rect 8352 9120 8358 9132
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 9674 9160 9680 9172
rect 9587 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9160 9738 9172
rect 10778 9160 10784 9172
rect 9732 9132 10784 9160
rect 9732 9120 9738 9132
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 11054 9160 11060 9172
rect 11015 9132 11060 9160
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 14384 9132 15669 9160
rect 8570 9092 8576 9104
rect 2746 9064 8576 9092
rect 2746 9036 2774 9064
rect 8570 9052 8576 9064
rect 8628 9052 8634 9104
rect 12989 9095 13047 9101
rect 12989 9061 13001 9095
rect 13035 9092 13047 9095
rect 14090 9092 14096 9104
rect 13035 9064 14096 9092
rect 13035 9061 13047 9064
rect 12989 9055 13047 9061
rect 14090 9052 14096 9064
rect 14148 9052 14154 9104
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 9024 2467 9027
rect 2746 9024 2780 9036
rect 2455 8996 2780 9024
rect 2455 8993 2467 8996
rect 2409 8987 2467 8993
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 4890 9024 4896 9036
rect 4851 8996 4896 9024
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 9024 6607 9027
rect 8294 9024 8300 9036
rect 6595 8996 8300 9024
rect 6595 8993 6607 8996
rect 6549 8987 6607 8993
rect 2314 8956 2320 8968
rect 2275 8928 2320 8956
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 4338 8916 4344 8968
rect 4396 8956 4402 8968
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 4396 8928 4537 8956
rect 4396 8916 4402 8928
rect 4525 8925 4537 8928
rect 4571 8956 4583 8959
rect 4798 8956 4804 8968
rect 4571 8928 4804 8956
rect 4571 8925 4583 8928
rect 4525 8919 4583 8925
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 5626 8956 5632 8968
rect 5000 8928 5632 8956
rect 5000 8888 5028 8928
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 7190 8956 7196 8968
rect 7151 8928 7196 8956
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 7300 8965 7328 8996
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 9508 8996 10241 9024
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 4724 8860 5028 8888
rect 5353 8891 5411 8897
rect 4614 8820 4620 8832
rect 4575 8792 4620 8820
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 4724 8829 4752 8860
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 5442 8888 5448 8900
rect 5399 8860 5448 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 7484 8888 7512 8919
rect 7558 8916 7564 8968
rect 7616 8956 7622 8968
rect 7616 8928 7661 8956
rect 7616 8916 7622 8928
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9508 8965 9536 8996
rect 10229 8993 10241 8996
rect 10275 9024 10287 9027
rect 13446 9024 13452 9036
rect 10275 8996 13452 9024
rect 10275 8993 10287 8996
rect 10229 8987 10287 8993
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 14384 9024 14412 9132
rect 15657 9129 15669 9132
rect 15703 9129 15715 9163
rect 15657 9123 15715 9129
rect 23109 9163 23167 9169
rect 23109 9129 23121 9163
rect 23155 9160 23167 9163
rect 23290 9160 23296 9172
rect 23155 9132 23296 9160
rect 23155 9129 23167 9132
rect 23109 9123 23167 9129
rect 23290 9120 23296 9132
rect 23348 9120 23354 9172
rect 24854 9120 24860 9172
rect 24912 9160 24918 9172
rect 24949 9163 25007 9169
rect 24949 9160 24961 9163
rect 24912 9132 24961 9160
rect 24912 9120 24918 9132
rect 24949 9129 24961 9132
rect 24995 9129 25007 9163
rect 24949 9123 25007 9129
rect 27249 9163 27307 9169
rect 27249 9129 27261 9163
rect 27295 9160 27307 9163
rect 27614 9160 27620 9172
rect 27295 9132 27620 9160
rect 27295 9129 27307 9132
rect 27249 9123 27307 9129
rect 27614 9120 27620 9132
rect 27672 9120 27678 9172
rect 27985 9163 28043 9169
rect 27985 9129 27997 9163
rect 28031 9160 28043 9163
rect 28074 9160 28080 9172
rect 28031 9132 28080 9160
rect 28031 9129 28043 9132
rect 27985 9123 28043 9129
rect 28074 9120 28080 9132
rect 28132 9160 28138 9172
rect 28350 9160 28356 9172
rect 28132 9132 28356 9160
rect 28132 9120 28138 9132
rect 28350 9120 28356 9132
rect 28408 9120 28414 9172
rect 28718 9160 28724 9172
rect 28679 9132 28724 9160
rect 28718 9120 28724 9132
rect 28776 9120 28782 9172
rect 14458 9052 14464 9104
rect 14516 9092 14522 9104
rect 14516 9064 17816 9092
rect 14516 9052 14522 9064
rect 17788 9036 17816 9064
rect 20622 9052 20628 9104
rect 20680 9092 20686 9104
rect 21269 9095 21327 9101
rect 21269 9092 21281 9095
rect 20680 9064 21281 9092
rect 20680 9052 20686 9064
rect 21269 9061 21281 9064
rect 21315 9092 21327 9095
rect 28166 9092 28172 9104
rect 21315 9064 28172 9092
rect 21315 9061 21327 9064
rect 21269 9055 21327 9061
rect 28166 9052 28172 9064
rect 28224 9092 28230 9104
rect 28534 9092 28540 9104
rect 28224 9064 28540 9092
rect 28224 9052 28230 9064
rect 28534 9052 28540 9064
rect 28592 9052 28598 9104
rect 13872 8996 14596 9024
rect 13872 8984 13878 8996
rect 9493 8959 9551 8965
rect 9493 8956 9505 8959
rect 9088 8928 9505 8956
rect 9088 8916 9094 8928
rect 9493 8925 9505 8928
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 9582 8916 9588 8968
rect 9640 8956 9646 8968
rect 9677 8959 9735 8965
rect 9677 8956 9689 8959
rect 9640 8928 9689 8956
rect 9640 8916 9646 8928
rect 9677 8925 9689 8928
rect 9723 8956 9735 8959
rect 14458 8956 14464 8968
rect 9723 8928 14464 8956
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 14568 8965 14596 8996
rect 14826 8984 14832 9036
rect 14884 8984 14890 9036
rect 15102 9024 15108 9036
rect 14936 8996 15108 9024
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 14701 8959 14759 8965
rect 14701 8925 14713 8959
rect 14747 8956 14759 8959
rect 14844 8956 14872 8984
rect 14747 8928 14872 8956
rect 14747 8925 14759 8928
rect 14701 8919 14759 8925
rect 13630 8888 13636 8900
rect 5736 8860 7512 8888
rect 7576 8860 13636 8888
rect 4709 8823 4767 8829
rect 4709 8789 4721 8823
rect 4755 8789 4767 8823
rect 4709 8783 4767 8789
rect 4982 8780 4988 8832
rect 5040 8820 5046 8832
rect 5736 8829 5764 8860
rect 5553 8823 5611 8829
rect 5553 8820 5565 8823
rect 5040 8792 5565 8820
rect 5040 8780 5046 8792
rect 5553 8789 5565 8792
rect 5599 8789 5611 8823
rect 5553 8783 5611 8789
rect 5721 8823 5779 8829
rect 5721 8789 5733 8823
rect 5767 8789 5779 8823
rect 5721 8783 5779 8789
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 7576 8820 7604 8860
rect 13630 8848 13636 8860
rect 13688 8848 13694 8900
rect 13722 8848 13728 8900
rect 13780 8888 13786 8900
rect 14936 8897 14964 8996
rect 15102 8984 15108 8996
rect 15160 8984 15166 9036
rect 17770 8984 17776 9036
rect 17828 9024 17834 9036
rect 23842 9024 23848 9036
rect 17828 8996 23848 9024
rect 17828 8984 17834 8996
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 25590 9024 25596 9036
rect 25551 8996 25596 9024
rect 25590 8984 25596 8996
rect 25648 8984 25654 9036
rect 15018 8959 15076 8965
rect 15018 8925 15030 8959
rect 15064 8956 15076 8959
rect 16022 8956 16028 8968
rect 15064 8928 16028 8956
rect 15064 8925 15076 8928
rect 15018 8919 15076 8925
rect 14829 8891 14887 8897
rect 14829 8888 14841 8891
rect 13780 8860 14841 8888
rect 13780 8848 13786 8860
rect 14829 8857 14841 8860
rect 14875 8857 14887 8891
rect 14829 8851 14887 8857
rect 14921 8891 14979 8897
rect 14921 8857 14933 8891
rect 14967 8857 14979 8891
rect 14921 8851 14979 8857
rect 6604 8792 7604 8820
rect 6604 8780 6610 8792
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 8478 8820 8484 8832
rect 8352 8792 8484 8820
rect 8352 8780 8358 8792
rect 8478 8780 8484 8792
rect 8536 8820 8542 8832
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 8536 8792 9045 8820
rect 8536 8780 8542 8792
rect 9033 8789 9045 8792
rect 9079 8820 9091 8823
rect 9582 8820 9588 8832
rect 9079 8792 9588 8820
rect 9079 8789 9091 8792
rect 9033 8783 9091 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 12894 8820 12900 8832
rect 12676 8792 12900 8820
rect 12676 8780 12682 8792
rect 12894 8780 12900 8792
rect 12952 8820 12958 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 12952 8792 13553 8820
rect 12952 8780 12958 8792
rect 13541 8789 13553 8792
rect 13587 8820 13599 8823
rect 15120 8820 15148 8928
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 17037 8959 17095 8965
rect 17037 8925 17049 8959
rect 17083 8956 17095 8959
rect 17586 8956 17592 8968
rect 17083 8928 17592 8956
rect 17083 8925 17095 8928
rect 17037 8919 17095 8925
rect 17586 8916 17592 8928
rect 17644 8956 17650 8968
rect 17681 8959 17739 8965
rect 17681 8956 17693 8959
rect 17644 8928 17693 8956
rect 17644 8916 17650 8928
rect 17681 8925 17693 8928
rect 17727 8925 17739 8959
rect 17681 8919 17739 8925
rect 25317 8959 25375 8965
rect 25317 8925 25329 8959
rect 25363 8956 25375 8959
rect 26418 8956 26424 8968
rect 25363 8928 26424 8956
rect 25363 8925 25375 8928
rect 25317 8919 25375 8925
rect 26418 8916 26424 8928
rect 26476 8916 26482 8968
rect 17865 8891 17923 8897
rect 17865 8857 17877 8891
rect 17911 8888 17923 8891
rect 25222 8888 25228 8900
rect 17911 8860 25228 8888
rect 17911 8857 17923 8860
rect 17865 8851 17923 8857
rect 25222 8848 25228 8860
rect 25280 8848 25286 8900
rect 13587 8792 15148 8820
rect 15197 8823 15255 8829
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 15197 8789 15209 8823
rect 15243 8820 15255 8823
rect 15470 8820 15476 8832
rect 15243 8792 15476 8820
rect 15243 8789 15255 8792
rect 15197 8783 15255 8789
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 17497 8823 17555 8829
rect 17497 8789 17509 8823
rect 17543 8820 17555 8823
rect 17586 8820 17592 8832
rect 17543 8792 17592 8820
rect 17543 8789 17555 8792
rect 17497 8783 17555 8789
rect 17586 8780 17592 8792
rect 17644 8780 17650 8832
rect 23661 8823 23719 8829
rect 23661 8789 23673 8823
rect 23707 8820 23719 8823
rect 23842 8820 23848 8832
rect 23707 8792 23848 8820
rect 23707 8789 23719 8792
rect 23661 8783 23719 8789
rect 23842 8780 23848 8792
rect 23900 8820 23906 8832
rect 24210 8820 24216 8832
rect 23900 8792 24216 8820
rect 23900 8780 23906 8792
rect 24210 8780 24216 8792
rect 24268 8780 24274 8832
rect 25406 8780 25412 8832
rect 25464 8820 25470 8832
rect 25464 8792 25509 8820
rect 25464 8780 25470 8792
rect 1104 8730 29600 8752
rect 1104 8678 8034 8730
rect 8086 8678 8098 8730
rect 8150 8678 8162 8730
rect 8214 8678 8226 8730
rect 8278 8678 8290 8730
rect 8342 8678 15118 8730
rect 15170 8678 15182 8730
rect 15234 8678 15246 8730
rect 15298 8678 15310 8730
rect 15362 8678 15374 8730
rect 15426 8678 22202 8730
rect 22254 8678 22266 8730
rect 22318 8678 22330 8730
rect 22382 8678 22394 8730
rect 22446 8678 22458 8730
rect 22510 8678 29286 8730
rect 29338 8678 29350 8730
rect 29402 8678 29414 8730
rect 29466 8678 29478 8730
rect 29530 8678 29542 8730
rect 29594 8678 29600 8730
rect 1104 8656 29600 8678
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 4982 8616 4988 8628
rect 4663 8588 4988 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 5442 8576 5448 8628
rect 5500 8616 5506 8628
rect 6365 8619 6423 8625
rect 6365 8616 6377 8619
rect 5500 8588 6377 8616
rect 5500 8576 5506 8588
rect 6365 8585 6377 8588
rect 6411 8585 6423 8619
rect 6365 8579 6423 8585
rect 7190 8576 7196 8628
rect 7248 8616 7254 8628
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 7248 8588 7481 8616
rect 7248 8576 7254 8588
rect 7469 8585 7481 8588
rect 7515 8616 7527 8619
rect 7515 8588 8708 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 1578 8548 1584 8560
rect 1539 8520 1584 8548
rect 1578 8508 1584 8520
rect 1636 8508 1642 8560
rect 4154 8548 4160 8560
rect 2746 8520 4160 8548
rect 2314 8440 2320 8492
rect 2372 8480 2378 8492
rect 2593 8483 2651 8489
rect 2593 8480 2605 8483
rect 2372 8452 2605 8480
rect 2372 8440 2378 8452
rect 2593 8449 2605 8452
rect 2639 8480 2651 8483
rect 2746 8480 2774 8520
rect 4154 8508 4160 8520
rect 4212 8508 4218 8560
rect 4890 8508 4896 8560
rect 4948 8508 4954 8560
rect 5718 8548 5724 8560
rect 5631 8520 5724 8548
rect 5718 8508 5724 8520
rect 5776 8548 5782 8560
rect 6546 8548 6552 8560
rect 5776 8520 6552 8548
rect 5776 8508 5782 8520
rect 6546 8508 6552 8520
rect 6604 8508 6610 8560
rect 7926 8508 7932 8560
rect 7984 8548 7990 8560
rect 8021 8551 8079 8557
rect 8021 8548 8033 8551
rect 7984 8520 8033 8548
rect 7984 8508 7990 8520
rect 8021 8517 8033 8520
rect 8067 8517 8079 8551
rect 8680 8548 8708 8588
rect 8754 8576 8760 8628
rect 8812 8616 8818 8628
rect 8812 8588 10180 8616
rect 8812 8576 8818 8588
rect 9766 8548 9772 8560
rect 8680 8520 9772 8548
rect 8021 8511 8079 8517
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 10152 8557 10180 8588
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 11112 8588 11529 8616
rect 11112 8576 11118 8588
rect 11517 8585 11529 8588
rect 11563 8585 11575 8619
rect 11517 8579 11575 8585
rect 14001 8619 14059 8625
rect 14001 8585 14013 8619
rect 14047 8616 14059 8619
rect 14826 8616 14832 8628
rect 14047 8588 14832 8616
rect 14047 8585 14059 8588
rect 14001 8579 14059 8585
rect 14826 8576 14832 8588
rect 14884 8576 14890 8628
rect 15470 8576 15476 8628
rect 15528 8576 15534 8628
rect 17218 8576 17224 8628
rect 17276 8616 17282 8628
rect 18049 8619 18107 8625
rect 18049 8616 18061 8619
rect 17276 8588 18061 8616
rect 17276 8576 17282 8588
rect 18049 8585 18061 8588
rect 18095 8585 18107 8619
rect 18049 8579 18107 8585
rect 21177 8619 21235 8625
rect 21177 8585 21189 8619
rect 21223 8616 21235 8619
rect 22094 8616 22100 8628
rect 21223 8588 22100 8616
rect 21223 8585 21235 8588
rect 21177 8579 21235 8585
rect 10137 8551 10195 8557
rect 10137 8517 10149 8551
rect 10183 8548 10195 8551
rect 12250 8548 12256 8560
rect 10183 8520 12256 8548
rect 10183 8517 10195 8520
rect 10137 8511 10195 8517
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 14918 8548 14924 8560
rect 14879 8520 14924 8548
rect 14918 8508 14924 8520
rect 14976 8508 14982 8560
rect 15488 8548 15516 8576
rect 15396 8520 15516 8548
rect 2639 8452 2774 8480
rect 2639 8449 2651 8452
rect 2593 8443 2651 8449
rect 2866 8440 2872 8492
rect 2924 8480 2930 8492
rect 4908 8480 4936 8508
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 2924 8452 2969 8480
rect 4908 8452 4997 8480
rect 2924 8440 2930 8452
rect 4985 8449 4997 8452
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8480 8263 8483
rect 8938 8480 8944 8492
rect 8251 8452 8944 8480
rect 8251 8449 8263 8452
rect 8205 8443 8263 8449
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8480 13875 8483
rect 13906 8480 13912 8492
rect 13863 8452 13912 8480
rect 13863 8449 13875 8452
rect 13817 8443 13875 8449
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8480 14059 8483
rect 14090 8480 14096 8492
rect 14047 8452 14096 8480
rect 14047 8449 14059 8452
rect 14001 8443 14059 8449
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 14642 8480 14648 8492
rect 14603 8452 14648 8480
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 14734 8440 14740 8492
rect 14792 8480 14798 8492
rect 15396 8489 15424 8520
rect 16666 8508 16672 8560
rect 16724 8548 16730 8560
rect 20070 8548 20076 8560
rect 16724 8520 17448 8548
rect 20031 8520 20076 8548
rect 16724 8508 16730 8520
rect 15381 8483 15439 8489
rect 14792 8452 14837 8480
rect 14792 8440 14798 8452
rect 15381 8449 15393 8483
rect 15427 8449 15439 8483
rect 15381 8443 15439 8449
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 15654 8480 15660 8492
rect 15528 8452 15573 8480
rect 15615 8452 15660 8480
rect 15528 8440 15534 8452
rect 15654 8440 15660 8452
rect 15712 8440 15718 8492
rect 17218 8480 17224 8492
rect 17179 8452 17224 8480
rect 17218 8440 17224 8452
rect 17276 8440 17282 8492
rect 17420 8489 17448 8520
rect 20070 8508 20076 8520
rect 20128 8508 20134 8560
rect 21192 8548 21220 8579
rect 22094 8576 22100 8588
rect 22152 8616 22158 8628
rect 22370 8616 22376 8628
rect 22152 8588 22376 8616
rect 22152 8576 22158 8588
rect 22370 8576 22376 8588
rect 22428 8576 22434 8628
rect 23014 8616 23020 8628
rect 22975 8588 23020 8616
rect 23014 8576 23020 8588
rect 23072 8576 23078 8628
rect 23658 8616 23664 8628
rect 23619 8588 23664 8616
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 25222 8616 25228 8628
rect 25183 8588 25228 8616
rect 25222 8576 25228 8588
rect 25280 8576 25286 8628
rect 25406 8576 25412 8628
rect 25464 8616 25470 8628
rect 25593 8619 25651 8625
rect 25593 8616 25605 8619
rect 25464 8588 25605 8616
rect 25464 8576 25470 8588
rect 25593 8585 25605 8588
rect 25639 8616 25651 8619
rect 26973 8619 27031 8625
rect 26973 8616 26985 8619
rect 25639 8588 26985 8616
rect 25639 8585 25651 8588
rect 25593 8579 25651 8585
rect 26973 8585 26985 8588
rect 27019 8585 27031 8619
rect 26973 8579 27031 8585
rect 27341 8619 27399 8625
rect 27341 8585 27353 8619
rect 27387 8616 27399 8619
rect 27430 8616 27436 8628
rect 27387 8588 27436 8616
rect 27387 8585 27399 8588
rect 27341 8579 27399 8585
rect 27430 8576 27436 8588
rect 27488 8576 27494 8628
rect 20364 8520 21220 8548
rect 21913 8551 21971 8557
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8449 17463 8483
rect 17586 8480 17592 8492
rect 17547 8452 17592 8480
rect 17405 8443 17463 8449
rect 1854 8372 1860 8424
rect 1912 8372 1918 8424
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8412 2835 8415
rect 4798 8412 4804 8424
rect 2823 8384 3464 8412
rect 4759 8384 4804 8412
rect 2823 8381 2835 8384
rect 2777 8375 2835 8381
rect 1872 8344 1900 8372
rect 2792 8344 2820 8375
rect 1872 8316 2820 8344
rect 3436 8288 3464 8384
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 5258 8412 5264 8424
rect 5123 8384 5264 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 4908 8344 4936 8375
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 5626 8372 5632 8424
rect 5684 8372 5690 8424
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 8628 8384 9321 8412
rect 8628 8372 8634 8384
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8412 9643 8415
rect 13078 8412 13084 8424
rect 9631 8384 12434 8412
rect 13039 8384 13084 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 5644 8344 5672 8372
rect 4908 8316 5672 8344
rect 12406 8344 12434 8384
rect 13078 8372 13084 8384
rect 13136 8372 13142 8424
rect 13630 8372 13636 8424
rect 13688 8412 13694 8424
rect 17236 8412 17264 8440
rect 13688 8384 17264 8412
rect 13688 8372 13694 8384
rect 17328 8356 17356 8443
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 20254 8480 20260 8492
rect 20215 8452 20260 8480
rect 20254 8440 20260 8452
rect 20312 8440 20318 8492
rect 20364 8489 20392 8520
rect 21913 8517 21925 8551
rect 21959 8548 21971 8551
rect 22646 8548 22652 8560
rect 21959 8520 22652 8548
rect 21959 8517 21971 8520
rect 21913 8511 21971 8517
rect 22646 8508 22652 8520
rect 22704 8508 22710 8560
rect 20349 8483 20407 8489
rect 20349 8449 20361 8483
rect 20395 8449 20407 8483
rect 20530 8480 20536 8492
rect 20491 8452 20536 8480
rect 20349 8443 20407 8449
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8480 20683 8483
rect 20990 8480 20996 8492
rect 20671 8452 20996 8480
rect 20671 8449 20683 8452
rect 20625 8443 20683 8449
rect 20990 8440 20996 8452
rect 21048 8440 21054 8492
rect 22094 8440 22100 8492
rect 22152 8480 22158 8492
rect 22373 8483 22431 8489
rect 22373 8480 22385 8483
rect 22152 8452 22385 8480
rect 22152 8440 22158 8452
rect 22373 8449 22385 8452
rect 22419 8480 22431 8483
rect 23032 8480 23060 8576
rect 22419 8452 23060 8480
rect 22419 8449 22431 8452
rect 22373 8443 22431 8449
rect 25590 8440 25596 8492
rect 25648 8480 25654 8492
rect 25648 8452 25820 8480
rect 25648 8440 25654 8452
rect 22281 8415 22339 8421
rect 22281 8381 22293 8415
rect 22327 8412 22339 8415
rect 22554 8412 22560 8424
rect 22327 8384 22560 8412
rect 22327 8381 22339 8384
rect 22281 8375 22339 8381
rect 22554 8372 22560 8384
rect 22612 8372 22618 8424
rect 25792 8421 25820 8452
rect 25685 8415 25743 8421
rect 25685 8381 25697 8415
rect 25731 8381 25743 8415
rect 25685 8375 25743 8381
rect 25777 8415 25835 8421
rect 25777 8381 25789 8415
rect 25823 8381 25835 8415
rect 27430 8412 27436 8424
rect 27391 8384 27436 8412
rect 25777 8375 25835 8381
rect 14461 8347 14519 8353
rect 14461 8344 14473 8347
rect 12406 8316 14473 8344
rect 14461 8313 14473 8316
rect 14507 8313 14519 8347
rect 14461 8307 14519 8313
rect 14844 8316 15148 8344
rect 1854 8276 1860 8288
rect 1815 8248 1860 8276
rect 1854 8236 1860 8248
rect 1912 8236 1918 8288
rect 1946 8236 1952 8288
rect 2004 8276 2010 8288
rect 2409 8279 2467 8285
rect 2409 8276 2421 8279
rect 2004 8248 2421 8276
rect 2004 8236 2010 8248
rect 2409 8245 2421 8248
rect 2455 8245 2467 8279
rect 2409 8239 2467 8245
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 3418 8276 3424 8288
rect 2832 8248 2877 8276
rect 3379 8248 3424 8276
rect 2832 8236 2838 8248
rect 3418 8236 3424 8248
rect 3476 8236 3482 8288
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 5258 8276 5264 8288
rect 4672 8248 5264 8276
rect 4672 8236 4678 8248
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 10686 8236 10692 8288
rect 10744 8276 10750 8288
rect 14844 8276 14872 8316
rect 10744 8248 14872 8276
rect 14921 8279 14979 8285
rect 10744 8236 10750 8248
rect 14921 8245 14933 8279
rect 14967 8276 14979 8279
rect 15010 8276 15016 8288
rect 14967 8248 15016 8276
rect 14967 8245 14979 8248
rect 14921 8239 14979 8245
rect 15010 8236 15016 8248
rect 15068 8236 15074 8288
rect 15120 8276 15148 8316
rect 15562 8304 15568 8356
rect 15620 8344 15626 8356
rect 15657 8347 15715 8353
rect 15657 8344 15669 8347
rect 15620 8316 15669 8344
rect 15620 8304 15626 8316
rect 15657 8313 15669 8316
rect 15703 8313 15715 8347
rect 15657 8307 15715 8313
rect 17310 8304 17316 8356
rect 17368 8304 17374 8356
rect 25590 8304 25596 8356
rect 25648 8344 25654 8356
rect 25700 8344 25728 8375
rect 27430 8372 27436 8384
rect 27488 8372 27494 8424
rect 27522 8372 27528 8424
rect 27580 8412 27586 8424
rect 27580 8384 27625 8412
rect 27580 8372 27586 8384
rect 25648 8316 25728 8344
rect 25648 8304 25654 8316
rect 16758 8276 16764 8288
rect 15120 8248 16764 8276
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 16942 8276 16948 8288
rect 16903 8248 16948 8276
rect 16942 8236 16948 8248
rect 17000 8236 17006 8288
rect 22373 8279 22431 8285
rect 22373 8245 22385 8279
rect 22419 8276 22431 8279
rect 22462 8276 22468 8288
rect 22419 8248 22468 8276
rect 22419 8245 22431 8248
rect 22373 8239 22431 8245
rect 22462 8236 22468 8248
rect 22520 8236 22526 8288
rect 22557 8279 22615 8285
rect 22557 8245 22569 8279
rect 22603 8276 22615 8279
rect 22830 8276 22836 8288
rect 22603 8248 22836 8276
rect 22603 8245 22615 8248
rect 22557 8239 22615 8245
rect 22830 8236 22836 8248
rect 22888 8236 22894 8288
rect 1104 8186 29440 8208
rect 1104 8134 4492 8186
rect 4544 8134 4556 8186
rect 4608 8134 4620 8186
rect 4672 8134 4684 8186
rect 4736 8134 4748 8186
rect 4800 8134 11576 8186
rect 11628 8134 11640 8186
rect 11692 8134 11704 8186
rect 11756 8134 11768 8186
rect 11820 8134 11832 8186
rect 11884 8134 18660 8186
rect 18712 8134 18724 8186
rect 18776 8134 18788 8186
rect 18840 8134 18852 8186
rect 18904 8134 18916 8186
rect 18968 8134 25744 8186
rect 25796 8134 25808 8186
rect 25860 8134 25872 8186
rect 25924 8134 25936 8186
rect 25988 8134 26000 8186
rect 26052 8134 29440 8186
rect 1104 8112 29440 8134
rect 1489 8075 1547 8081
rect 1489 8041 1501 8075
rect 1535 8072 1547 8075
rect 1578 8072 1584 8084
rect 1535 8044 1584 8072
rect 1535 8041 1547 8044
rect 1489 8035 1547 8041
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 2225 8075 2283 8081
rect 2225 8041 2237 8075
rect 2271 8072 2283 8075
rect 2958 8072 2964 8084
rect 2271 8044 2964 8072
rect 2271 8041 2283 8044
rect 2225 8035 2283 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 6178 8072 6184 8084
rect 4448 8044 6184 8072
rect 2133 8007 2191 8013
rect 2133 7973 2145 8007
rect 2179 8004 2191 8007
rect 4448 8004 4476 8044
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 8938 8072 8944 8084
rect 8899 8044 8944 8072
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 11241 8075 11299 8081
rect 11241 8041 11253 8075
rect 11287 8072 11299 8075
rect 12434 8072 12440 8084
rect 11287 8044 12440 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 13078 8032 13084 8084
rect 13136 8072 13142 8084
rect 15473 8075 15531 8081
rect 13136 8044 15148 8072
rect 13136 8032 13142 8044
rect 4982 8004 4988 8016
rect 2179 7976 4476 8004
rect 4724 7976 4988 8004
rect 2179 7973 2191 7976
rect 2133 7967 2191 7973
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7936 2375 7939
rect 2498 7936 2504 7948
rect 2363 7908 2504 7936
rect 2363 7905 2375 7908
rect 2317 7899 2375 7905
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 4724 7945 4752 7976
rect 4982 7964 4988 7976
rect 5040 8004 5046 8016
rect 5166 8004 5172 8016
rect 5040 7976 5172 8004
rect 5040 7964 5046 7976
rect 5166 7964 5172 7976
rect 5224 7964 5230 8016
rect 5350 7964 5356 8016
rect 5408 8004 5414 8016
rect 5997 8007 6055 8013
rect 5997 8004 6009 8007
rect 5408 7976 6009 8004
rect 5408 7964 5414 7976
rect 5997 7973 6009 7976
rect 6043 7973 6055 8007
rect 5997 7967 6055 7973
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 5718 7936 5724 7948
rect 5123 7908 5724 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 6181 7939 6239 7945
rect 6181 7905 6193 7939
rect 6227 7936 6239 7939
rect 6227 7908 9536 7936
rect 6227 7905 6239 7908
rect 6181 7899 6239 7905
rect 1946 7868 1952 7880
rect 1907 7840 1952 7868
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 4614 7868 4620 7880
rect 4575 7840 4620 7868
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 4982 7868 4988 7880
rect 4943 7840 4988 7868
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 9122 7868 9128 7880
rect 9083 7840 9128 7868
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9508 7877 9536 7908
rect 9858 7896 9864 7948
rect 9916 7936 9922 7948
rect 10781 7939 10839 7945
rect 10781 7936 10793 7939
rect 9916 7908 10793 7936
rect 9916 7896 9922 7908
rect 10781 7905 10793 7908
rect 10827 7905 10839 7939
rect 13096 7936 13124 8032
rect 14090 8004 14096 8016
rect 14051 7976 14096 8004
rect 14090 7964 14096 7976
rect 14148 8004 14154 8016
rect 14458 8004 14464 8016
rect 14148 7976 14464 8004
rect 14148 7964 14154 7976
rect 14458 7964 14464 7976
rect 14516 7964 14522 8016
rect 14826 7964 14832 8016
rect 14884 8004 14890 8016
rect 15120 8004 15148 8044
rect 15473 8041 15485 8075
rect 15519 8072 15531 8075
rect 15654 8072 15660 8084
rect 15519 8044 15660 8072
rect 15519 8041 15531 8044
rect 15473 8035 15531 8041
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 17129 8075 17187 8081
rect 17129 8072 17141 8075
rect 15804 8044 17141 8072
rect 15804 8032 15810 8044
rect 17129 8041 17141 8044
rect 17175 8072 17187 8075
rect 19610 8072 19616 8084
rect 17175 8044 19616 8072
rect 17175 8041 17187 8044
rect 17129 8035 17187 8041
rect 19610 8032 19616 8044
rect 19668 8072 19674 8084
rect 20990 8072 20996 8084
rect 19668 8044 20576 8072
rect 20951 8044 20996 8072
rect 19668 8032 19674 8044
rect 14884 7976 15056 8004
rect 15120 7976 16160 8004
rect 14884 7964 14890 7976
rect 15028 7945 15056 7976
rect 10781 7899 10839 7905
rect 12406 7908 13124 7936
rect 15013 7939 15071 7945
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7837 9551 7871
rect 10870 7868 10876 7880
rect 10831 7840 10876 7868
rect 9493 7831 9551 7837
rect 5261 7803 5319 7809
rect 5261 7769 5273 7803
rect 5307 7800 5319 7803
rect 5721 7803 5779 7809
rect 5721 7800 5733 7803
rect 5307 7772 5733 7800
rect 5307 7769 5319 7772
rect 5261 7763 5319 7769
rect 5721 7769 5733 7772
rect 5767 7769 5779 7803
rect 5721 7763 5779 7769
rect 7926 7760 7932 7812
rect 7984 7800 7990 7812
rect 9232 7800 9260 7831
rect 7984 7772 9260 7800
rect 9416 7800 9444 7831
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 11146 7800 11152 7812
rect 9416 7772 11152 7800
rect 7984 7760 7990 7772
rect 11146 7760 11152 7772
rect 11204 7760 11210 7812
rect 2038 7732 2044 7744
rect 1999 7704 2044 7732
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2958 7732 2964 7744
rect 2919 7704 2964 7732
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 4893 7735 4951 7741
rect 4893 7701 4905 7735
rect 4939 7732 4951 7735
rect 5074 7732 5080 7744
rect 4939 7704 5080 7732
rect 4939 7701 4951 7704
rect 4893 7695 4951 7701
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 10134 7732 10140 7744
rect 10095 7704 10140 7732
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 10318 7692 10324 7744
rect 10376 7732 10382 7744
rect 11701 7735 11759 7741
rect 11701 7732 11713 7735
rect 10376 7704 11713 7732
rect 10376 7692 10382 7704
rect 11701 7701 11713 7704
rect 11747 7732 11759 7735
rect 12406 7732 12434 7908
rect 15013 7905 15025 7939
rect 15059 7905 15071 7939
rect 15013 7899 15071 7905
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7868 14887 7871
rect 15470 7868 15476 7880
rect 14875 7840 15476 7868
rect 14875 7837 14887 7840
rect 14829 7831 14887 7837
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 15654 7877 15660 7880
rect 15652 7868 15660 7877
rect 15615 7840 15660 7868
rect 15652 7831 15660 7840
rect 15654 7828 15660 7831
rect 15712 7828 15718 7880
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 13541 7803 13599 7809
rect 13541 7769 13553 7803
rect 13587 7800 13599 7803
rect 13906 7800 13912 7812
rect 13587 7772 13912 7800
rect 13587 7769 13599 7772
rect 13541 7763 13599 7769
rect 13906 7760 13912 7772
rect 13964 7800 13970 7812
rect 15764 7800 15792 7831
rect 15930 7828 15936 7880
rect 15988 7877 15994 7880
rect 16132 7877 16160 7976
rect 19978 7936 19984 7948
rect 19260 7908 19984 7936
rect 19260 7877 19288 7908
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 20548 7945 20576 8044
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 22462 8072 22468 8084
rect 22423 8044 22468 8072
rect 22462 8032 22468 8044
rect 22520 8032 22526 8084
rect 25590 8032 25596 8084
rect 25648 8072 25654 8084
rect 25961 8075 26019 8081
rect 25961 8072 25973 8075
rect 25648 8044 25973 8072
rect 25648 8032 25654 8044
rect 25961 8041 25973 8044
rect 26007 8041 26019 8075
rect 25961 8035 26019 8041
rect 26142 8032 26148 8084
rect 26200 8072 26206 8084
rect 27157 8075 27215 8081
rect 27157 8072 27169 8075
rect 26200 8044 27169 8072
rect 26200 8032 26206 8044
rect 27157 8041 27169 8044
rect 27203 8041 27215 8075
rect 27157 8035 27215 8041
rect 27522 7964 27528 8016
rect 27580 7964 27586 8016
rect 20533 7939 20591 7945
rect 20533 7905 20545 7939
rect 20579 7936 20591 7939
rect 22005 7939 22063 7945
rect 22005 7936 22017 7939
rect 20579 7908 22017 7936
rect 20579 7905 20591 7908
rect 20533 7899 20591 7905
rect 15988 7871 16027 7877
rect 16015 7837 16027 7871
rect 15988 7831 16027 7837
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7837 16175 7871
rect 16117 7831 16175 7837
rect 19245 7871 19303 7877
rect 19245 7837 19257 7871
rect 19291 7837 19303 7871
rect 19426 7868 19432 7880
rect 19387 7840 19432 7868
rect 19245 7831 19303 7837
rect 15988 7828 15994 7831
rect 13964 7772 15792 7800
rect 13964 7760 13970 7772
rect 15764 7744 15792 7772
rect 15838 7760 15844 7812
rect 15896 7800 15902 7812
rect 16132 7800 16160 7831
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 21266 7868 21272 7880
rect 21227 7840 21272 7868
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 21928 7868 21956 7908
rect 22005 7905 22017 7908
rect 22051 7905 22063 7939
rect 22005 7899 22063 7905
rect 22097 7939 22155 7945
rect 22097 7905 22109 7939
rect 22143 7936 22155 7939
rect 23658 7936 23664 7948
rect 22143 7908 23664 7936
rect 22143 7905 22155 7908
rect 22097 7899 22155 7905
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 26605 7939 26663 7945
rect 26605 7905 26617 7939
rect 26651 7936 26663 7939
rect 27540 7936 27568 7964
rect 27709 7939 27767 7945
rect 27709 7936 27721 7939
rect 26651 7908 27721 7936
rect 26651 7905 26663 7908
rect 26605 7899 26663 7905
rect 27709 7905 27721 7908
rect 27755 7905 27767 7939
rect 27709 7899 27767 7905
rect 22189 7871 22247 7877
rect 21928 7840 22048 7868
rect 22189 7862 22201 7871
rect 16669 7803 16727 7809
rect 16669 7800 16681 7803
rect 15896 7772 15941 7800
rect 16132 7772 16681 7800
rect 15896 7760 15902 7772
rect 16669 7769 16681 7772
rect 16715 7800 16727 7803
rect 20346 7800 20352 7812
rect 16715 7772 20352 7800
rect 16715 7769 16727 7772
rect 16669 7763 16727 7769
rect 20346 7760 20352 7772
rect 20404 7760 20410 7812
rect 20993 7803 21051 7809
rect 20993 7769 21005 7803
rect 21039 7800 21051 7803
rect 21910 7800 21916 7812
rect 21039 7772 21916 7800
rect 21039 7769 21051 7772
rect 20993 7763 21051 7769
rect 21910 7760 21916 7772
rect 21968 7760 21974 7812
rect 12986 7732 12992 7744
rect 11747 7704 12434 7732
rect 12947 7704 12992 7732
rect 11747 7701 11759 7704
rect 11701 7695 11759 7701
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 14274 7692 14280 7744
rect 14332 7732 14338 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 14332 7704 14657 7732
rect 14332 7692 14338 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 14645 7695 14703 7701
rect 15746 7692 15752 7744
rect 15804 7692 15810 7744
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 17865 7735 17923 7741
rect 17865 7732 17877 7735
rect 16080 7704 17877 7732
rect 16080 7692 16086 7704
rect 17865 7701 17877 7704
rect 17911 7732 17923 7735
rect 18230 7732 18236 7744
rect 17911 7704 18236 7732
rect 17911 7701 17923 7704
rect 17865 7695 17923 7701
rect 18230 7692 18236 7704
rect 18288 7732 18294 7744
rect 18601 7735 18659 7741
rect 18601 7732 18613 7735
rect 18288 7704 18613 7732
rect 18288 7692 18294 7704
rect 18601 7701 18613 7704
rect 18647 7701 18659 7735
rect 18601 7695 18659 7701
rect 19337 7735 19395 7741
rect 19337 7701 19349 7735
rect 19383 7732 19395 7735
rect 19426 7732 19432 7744
rect 19383 7704 19432 7732
rect 19383 7701 19395 7704
rect 19337 7695 19395 7701
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 19978 7732 19984 7744
rect 19939 7704 19984 7732
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 21174 7732 21180 7744
rect 21135 7704 21180 7732
rect 21174 7692 21180 7704
rect 21232 7692 21238 7744
rect 22020 7732 22048 7840
rect 22112 7837 22201 7862
rect 22235 7837 22247 7871
rect 22112 7834 22247 7837
rect 22112 7800 22140 7834
rect 22189 7831 22247 7834
rect 22280 7871 22338 7877
rect 22280 7837 22292 7871
rect 22326 7862 22338 7871
rect 22646 7868 22652 7880
rect 22388 7862 22652 7868
rect 22326 7840 22652 7862
rect 22326 7837 22416 7840
rect 22280 7834 22416 7837
rect 22280 7831 22338 7834
rect 22646 7828 22652 7840
rect 22704 7868 22710 7880
rect 22925 7871 22983 7877
rect 22925 7868 22937 7871
rect 22704 7840 22937 7868
rect 22704 7828 22710 7840
rect 22925 7837 22937 7840
rect 22971 7837 22983 7871
rect 22925 7831 22983 7837
rect 23842 7828 23848 7880
rect 23900 7868 23906 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 23900 7840 24409 7868
rect 23900 7828 23906 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 27430 7828 27436 7880
rect 27488 7868 27494 7880
rect 27525 7871 27583 7877
rect 27525 7868 27537 7871
rect 27488 7840 27537 7868
rect 27488 7828 27494 7840
rect 27525 7837 27537 7840
rect 27571 7837 27583 7871
rect 27525 7831 27583 7837
rect 23860 7800 23888 7828
rect 22112 7772 23888 7800
rect 26329 7803 26387 7809
rect 26329 7769 26341 7803
rect 26375 7800 26387 7803
rect 27617 7803 27675 7809
rect 27617 7800 27629 7803
rect 26375 7772 27629 7800
rect 26375 7769 26387 7772
rect 26329 7763 26387 7769
rect 27617 7769 27629 7772
rect 27663 7800 27675 7803
rect 27706 7800 27712 7812
rect 27663 7772 27712 7800
rect 27663 7769 27675 7772
rect 27617 7763 27675 7769
rect 27706 7760 27712 7772
rect 27764 7760 27770 7812
rect 28442 7800 28448 7812
rect 28403 7772 28448 7800
rect 28442 7760 28448 7772
rect 28500 7760 28506 7812
rect 28629 7803 28687 7809
rect 28629 7769 28641 7803
rect 28675 7800 28687 7803
rect 28718 7800 28724 7812
rect 28675 7772 28724 7800
rect 28675 7769 28687 7772
rect 28629 7763 28687 7769
rect 28718 7760 28724 7772
rect 28776 7760 28782 7812
rect 22738 7732 22744 7744
rect 22020 7704 22744 7732
rect 22738 7692 22744 7704
rect 22796 7732 22802 7744
rect 23569 7735 23627 7741
rect 23569 7732 23581 7735
rect 22796 7704 23581 7732
rect 22796 7692 22802 7704
rect 23569 7701 23581 7704
rect 23615 7732 23627 7735
rect 23750 7732 23756 7744
rect 23615 7704 23756 7732
rect 23615 7701 23627 7704
rect 23569 7695 23627 7701
rect 23750 7692 23756 7704
rect 23808 7692 23814 7744
rect 25958 7692 25964 7744
rect 26016 7732 26022 7744
rect 26421 7735 26479 7741
rect 26421 7732 26433 7735
rect 26016 7704 26433 7732
rect 26016 7692 26022 7704
rect 26421 7701 26433 7704
rect 26467 7701 26479 7735
rect 26421 7695 26479 7701
rect 1104 7642 29600 7664
rect 1104 7590 8034 7642
rect 8086 7590 8098 7642
rect 8150 7590 8162 7642
rect 8214 7590 8226 7642
rect 8278 7590 8290 7642
rect 8342 7590 15118 7642
rect 15170 7590 15182 7642
rect 15234 7590 15246 7642
rect 15298 7590 15310 7642
rect 15362 7590 15374 7642
rect 15426 7590 22202 7642
rect 22254 7590 22266 7642
rect 22318 7590 22330 7642
rect 22382 7590 22394 7642
rect 22446 7590 22458 7642
rect 22510 7590 29286 7642
rect 29338 7590 29350 7642
rect 29402 7590 29414 7642
rect 29466 7590 29478 7642
rect 29530 7590 29542 7642
rect 29594 7590 29600 7642
rect 1104 7568 29600 7590
rect 5350 7528 5356 7540
rect 5311 7500 5356 7528
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 7926 7528 7932 7540
rect 7887 7500 7932 7528
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 8846 7528 8852 7540
rect 8128 7500 8852 7528
rect 8128 7460 8156 7500
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9217 7531 9275 7537
rect 9217 7528 9229 7531
rect 9180 7500 9229 7528
rect 9180 7488 9186 7500
rect 9217 7497 9229 7500
rect 9263 7497 9275 7531
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 9217 7491 9275 7497
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 11054 7528 11060 7540
rect 10428 7500 11060 7528
rect 7392 7432 8156 7460
rect 8220 7432 9076 7460
rect 4982 7392 4988 7404
rect 4895 7364 4988 7392
rect 4982 7352 4988 7364
rect 5040 7392 5046 7404
rect 6457 7395 6515 7401
rect 6457 7392 6469 7395
rect 5040 7364 6469 7392
rect 5040 7352 5046 7364
rect 6457 7361 6469 7364
rect 6503 7361 6515 7395
rect 6457 7355 6515 7361
rect 6546 7352 6552 7404
rect 6604 7392 6610 7404
rect 6604 7364 6649 7392
rect 6604 7352 6610 7364
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 4672 7296 4905 7324
rect 4672 7284 4678 7296
rect 4893 7293 4905 7296
rect 4939 7293 4951 7327
rect 5074 7324 5080 7336
rect 5035 7296 5080 7324
rect 4893 7287 4951 7293
rect 4908 7256 4936 7287
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 5166 7284 5172 7336
rect 5224 7324 5230 7336
rect 5224 7296 5269 7324
rect 5224 7284 5230 7296
rect 7190 7284 7196 7336
rect 7248 7324 7254 7336
rect 7392 7333 7420 7432
rect 8220 7401 8248 7432
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8754 7392 8760 7404
rect 8715 7364 8760 7392
rect 8205 7355 8263 7361
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 9048 7401 9076 7432
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9214 7392 9220 7404
rect 9079 7364 9220 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 10318 7392 10324 7404
rect 10279 7364 10324 7392
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 10428 7401 10456 7500
rect 11054 7488 11060 7500
rect 11112 7528 11118 7540
rect 11330 7528 11336 7540
rect 11112 7500 11336 7528
rect 11112 7488 11118 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12526 7528 12532 7540
rect 12299 7500 12532 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 14553 7531 14611 7537
rect 14292 7500 14504 7528
rect 10686 7420 10692 7472
rect 10744 7460 10750 7472
rect 12621 7463 12679 7469
rect 12621 7460 12633 7463
rect 10744 7432 10789 7460
rect 12176 7432 12633 7460
rect 10744 7420 10750 7432
rect 10414 7395 10472 7401
rect 10414 7361 10426 7395
rect 10460 7361 10472 7395
rect 10594 7392 10600 7404
rect 10555 7364 10600 7392
rect 10414 7355 10472 7361
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 10786 7395 10844 7401
rect 10786 7361 10798 7395
rect 10832 7361 10844 7395
rect 10786 7355 10844 7361
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 7248 7296 7389 7324
rect 7248 7284 7254 7296
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 7377 7287 7435 7293
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8941 7327 8999 7333
rect 8941 7324 8953 7327
rect 8159 7296 8953 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8941 7293 8953 7296
rect 8987 7324 8999 7327
rect 9398 7324 9404 7336
rect 8987 7296 9404 7324
rect 8987 7293 8999 7296
rect 8941 7287 8999 7293
rect 4982 7256 4988 7268
rect 4908 7228 4988 7256
rect 4982 7216 4988 7228
rect 5040 7216 5046 7268
rect 7944 7256 7972 7287
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 9766 7284 9772 7336
rect 9824 7324 9830 7336
rect 10796 7324 10824 7355
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 12176 7392 12204 7432
rect 12621 7429 12633 7432
rect 12667 7460 12679 7463
rect 12986 7460 12992 7472
rect 12667 7432 12992 7460
rect 12667 7429 12679 7432
rect 12621 7423 12679 7429
rect 12986 7420 12992 7432
rect 13044 7460 13050 7472
rect 13044 7432 14136 7460
rect 13044 7420 13050 7432
rect 11020 7364 12204 7392
rect 12391 7395 12449 7401
rect 11020 7352 11026 7364
rect 12391 7361 12403 7395
rect 12437 7361 12449 7395
rect 12391 7355 12449 7361
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7361 12587 7395
rect 12529 7355 12587 7361
rect 9824 7296 10824 7324
rect 9824 7284 9830 7296
rect 8849 7259 8907 7265
rect 8849 7256 8861 7259
rect 7944 7228 8861 7256
rect 8849 7225 8861 7228
rect 8895 7256 8907 7259
rect 9306 7256 9312 7268
rect 8895 7228 9312 7256
rect 8895 7225 8907 7228
rect 8849 7219 8907 7225
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 10870 7216 10876 7268
rect 10928 7256 10934 7268
rect 11701 7259 11759 7265
rect 11701 7256 11713 7259
rect 10928 7228 11713 7256
rect 10928 7216 10934 7228
rect 11701 7225 11713 7228
rect 11747 7256 11759 7259
rect 12406 7256 12434 7355
rect 12544 7324 12572 7355
rect 12710 7352 12716 7404
rect 12768 7401 12774 7404
rect 12768 7395 12807 7401
rect 12795 7361 12807 7395
rect 12768 7355 12807 7361
rect 12768 7352 12774 7355
rect 12894 7352 12900 7404
rect 12952 7392 12958 7404
rect 14108 7392 14136 7432
rect 14182 7420 14188 7472
rect 14240 7460 14246 7472
rect 14292 7460 14320 7500
rect 14240 7432 14333 7460
rect 14240 7420 14246 7432
rect 14366 7420 14372 7472
rect 14424 7469 14430 7472
rect 14424 7463 14443 7469
rect 14431 7429 14443 7463
rect 14476 7460 14504 7500
rect 14553 7497 14565 7531
rect 14599 7528 14611 7531
rect 14642 7528 14648 7540
rect 14599 7500 14648 7528
rect 14599 7497 14611 7500
rect 14553 7491 14611 7497
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 17862 7488 17868 7540
rect 17920 7528 17926 7540
rect 18325 7531 18383 7537
rect 18325 7528 18337 7531
rect 17920 7500 18337 7528
rect 17920 7488 17926 7500
rect 18325 7497 18337 7500
rect 18371 7497 18383 7531
rect 18325 7491 18383 7497
rect 19429 7531 19487 7537
rect 19429 7497 19441 7531
rect 19475 7497 19487 7531
rect 19429 7491 19487 7497
rect 14734 7460 14740 7472
rect 14476 7432 14740 7460
rect 14424 7423 14443 7429
rect 14424 7420 14430 7423
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 19444 7460 19472 7491
rect 19518 7488 19524 7540
rect 19576 7528 19582 7540
rect 20070 7528 20076 7540
rect 19576 7500 20076 7528
rect 19576 7488 19582 7500
rect 19720 7469 19748 7500
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 21910 7528 21916 7540
rect 21871 7500 21916 7528
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 25130 7488 25136 7540
rect 25188 7528 25194 7540
rect 25958 7528 25964 7540
rect 25188 7500 25964 7528
rect 25188 7488 25194 7500
rect 25958 7488 25964 7500
rect 26016 7488 26022 7540
rect 27249 7531 27307 7537
rect 27249 7497 27261 7531
rect 27295 7528 27307 7531
rect 27430 7528 27436 7540
rect 27295 7500 27436 7528
rect 27295 7497 27307 7500
rect 27249 7491 27307 7497
rect 27430 7488 27436 7500
rect 27488 7488 27494 7540
rect 27706 7528 27712 7540
rect 27667 7500 27712 7528
rect 27706 7488 27712 7500
rect 27764 7488 27770 7540
rect 18524 7432 19472 7460
rect 19705 7463 19763 7469
rect 16942 7392 16948 7404
rect 12952 7364 12997 7392
rect 14108 7364 16804 7392
rect 16903 7364 16948 7392
rect 12952 7352 12958 7364
rect 13170 7324 13176 7336
rect 12544 7296 13176 7324
rect 13170 7284 13176 7296
rect 13228 7324 13234 7336
rect 13357 7327 13415 7333
rect 13357 7324 13369 7327
rect 13228 7296 13369 7324
rect 13228 7284 13234 7296
rect 13357 7293 13369 7296
rect 13403 7293 13415 7327
rect 16666 7324 16672 7336
rect 16627 7296 16672 7324
rect 13357 7287 13415 7293
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 16776 7324 16804 7364
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 17218 7392 17224 7404
rect 17179 7364 17224 7392
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 17770 7392 17776 7404
rect 17731 7364 17776 7392
rect 17770 7352 17776 7364
rect 17828 7352 17834 7404
rect 18524 7401 18552 7432
rect 19705 7429 19717 7463
rect 19751 7429 19763 7463
rect 19705 7423 19763 7429
rect 19797 7463 19855 7469
rect 19797 7429 19809 7463
rect 19843 7460 19855 7463
rect 20438 7460 20444 7472
rect 19843 7432 20444 7460
rect 19843 7429 19855 7432
rect 19797 7423 19855 7429
rect 20438 7420 20444 7432
rect 20496 7420 20502 7472
rect 21177 7463 21235 7469
rect 21177 7429 21189 7463
rect 21223 7460 21235 7463
rect 22094 7460 22100 7472
rect 21223 7432 22100 7460
rect 21223 7429 21235 7432
rect 21177 7423 21235 7429
rect 18509 7395 18567 7401
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 18785 7395 18843 7401
rect 18785 7392 18797 7395
rect 18656 7364 18797 7392
rect 18656 7352 18662 7364
rect 18785 7361 18797 7364
rect 18831 7361 18843 7395
rect 18785 7355 18843 7361
rect 18969 7395 19027 7401
rect 18969 7361 18981 7395
rect 19015 7392 19027 7395
rect 19426 7392 19432 7404
rect 19015 7364 19432 7392
rect 19015 7361 19027 7364
rect 18969 7355 19027 7361
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 19610 7401 19616 7404
rect 19608 7392 19616 7401
rect 19571 7364 19616 7392
rect 19608 7355 19616 7364
rect 19610 7352 19616 7355
rect 19668 7352 19674 7404
rect 19980 7395 20038 7401
rect 19980 7361 19992 7395
rect 20026 7361 20038 7395
rect 19980 7355 20038 7361
rect 20073 7395 20131 7401
rect 20073 7361 20085 7395
rect 20119 7392 20131 7395
rect 20346 7392 20352 7404
rect 20119 7364 20352 7392
rect 20119 7361 20131 7364
rect 20073 7355 20131 7361
rect 17126 7324 17132 7336
rect 16776 7296 17132 7324
rect 17126 7284 17132 7296
rect 17184 7284 17190 7336
rect 19996 7324 20024 7355
rect 20346 7352 20352 7364
rect 20404 7392 20410 7404
rect 21192 7392 21220 7423
rect 22094 7420 22100 7432
rect 22152 7420 22158 7472
rect 28718 7460 28724 7472
rect 28679 7432 28724 7460
rect 28718 7420 28724 7432
rect 28776 7420 28782 7472
rect 22830 7392 22836 7404
rect 20404 7364 21220 7392
rect 22791 7364 22836 7392
rect 20404 7352 20410 7364
rect 22830 7352 22836 7364
rect 22888 7352 22894 7404
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7361 23535 7395
rect 23477 7355 23535 7361
rect 20625 7327 20683 7333
rect 20625 7324 20637 7327
rect 19306 7296 20637 7324
rect 12618 7256 12624 7268
rect 11747 7228 12624 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 15289 7259 15347 7265
rect 15289 7256 15301 7259
rect 13280 7228 15301 7256
rect 1854 7148 1860 7200
rect 1912 7188 1918 7200
rect 10134 7188 10140 7200
rect 1912 7160 10140 7188
rect 1912 7148 1918 7160
rect 10134 7148 10140 7160
rect 10192 7188 10198 7200
rect 10686 7188 10692 7200
rect 10192 7160 10692 7188
rect 10192 7148 10198 7160
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11238 7188 11244 7200
rect 11011 7160 11244 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11238 7148 11244 7160
rect 11296 7148 11302 7200
rect 11330 7148 11336 7200
rect 11388 7188 11394 7200
rect 12342 7188 12348 7200
rect 11388 7160 12348 7188
rect 11388 7148 11394 7160
rect 12342 7148 12348 7160
rect 12400 7188 12406 7200
rect 13280 7188 13308 7228
rect 15289 7225 15301 7228
rect 15335 7256 15347 7259
rect 15930 7256 15936 7268
rect 15335 7228 15936 7256
rect 15335 7225 15347 7228
rect 15289 7219 15347 7225
rect 15930 7216 15936 7228
rect 15988 7256 15994 7268
rect 19306 7256 19334 7296
rect 20625 7293 20637 7296
rect 20671 7324 20683 7327
rect 22646 7324 22652 7336
rect 20671 7296 22652 7324
rect 20671 7293 20683 7296
rect 20625 7287 20683 7293
rect 22646 7284 22652 7296
rect 22704 7284 22710 7336
rect 22741 7327 22799 7333
rect 22741 7293 22753 7327
rect 22787 7324 22799 7327
rect 23198 7324 23204 7336
rect 22787 7296 23204 7324
rect 22787 7293 22799 7296
rect 22741 7287 22799 7293
rect 23198 7284 23204 7296
rect 23256 7284 23262 7336
rect 15988 7228 19334 7256
rect 15988 7216 15994 7228
rect 20806 7216 20812 7268
rect 20864 7256 20870 7268
rect 23492 7256 23520 7355
rect 23566 7352 23572 7404
rect 23624 7392 23630 7404
rect 23624 7364 23669 7392
rect 23624 7352 23630 7364
rect 25498 7352 25504 7404
rect 25556 7392 25562 7404
rect 25685 7395 25743 7401
rect 25685 7392 25697 7395
rect 25556 7364 25697 7392
rect 25556 7352 25562 7364
rect 25685 7361 25697 7364
rect 25731 7392 25743 7395
rect 26973 7395 27031 7401
rect 26973 7392 26985 7395
rect 25731 7364 26985 7392
rect 25731 7361 25743 7364
rect 25685 7355 25743 7361
rect 26973 7361 26985 7364
rect 27019 7392 27031 7395
rect 27985 7395 28043 7401
rect 27985 7392 27997 7395
rect 27019 7364 27997 7392
rect 27019 7361 27031 7364
rect 26973 7355 27031 7361
rect 27985 7361 27997 7364
rect 28031 7361 28043 7395
rect 27985 7355 28043 7361
rect 25961 7327 26019 7333
rect 25961 7293 25973 7327
rect 26007 7324 26019 7327
rect 27154 7324 27160 7336
rect 26007 7296 27160 7324
rect 26007 7293 26019 7296
rect 25961 7287 26019 7293
rect 27154 7284 27160 7296
rect 27212 7324 27218 7336
rect 27249 7327 27307 7333
rect 27249 7324 27261 7327
rect 27212 7296 27261 7324
rect 27212 7284 27218 7296
rect 27249 7293 27261 7296
rect 27295 7324 27307 7327
rect 27709 7327 27767 7333
rect 27709 7324 27721 7327
rect 27295 7296 27721 7324
rect 27295 7293 27307 7296
rect 27249 7287 27307 7293
rect 27709 7293 27721 7296
rect 27755 7293 27767 7327
rect 27709 7287 27767 7293
rect 20864 7228 23520 7256
rect 20864 7216 20870 7228
rect 12400 7160 13308 7188
rect 12400 7148 12406 7160
rect 14090 7148 14096 7200
rect 14148 7188 14154 7200
rect 14369 7191 14427 7197
rect 14369 7188 14381 7191
rect 14148 7160 14381 7188
rect 14148 7148 14154 7160
rect 14369 7157 14381 7160
rect 14415 7157 14427 7191
rect 14369 7151 14427 7157
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 15841 7191 15899 7197
rect 15841 7188 15853 7191
rect 15804 7160 15853 7188
rect 15804 7148 15810 7160
rect 15841 7157 15853 7160
rect 15887 7188 15899 7191
rect 17034 7188 17040 7200
rect 15887 7160 17040 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 19334 7148 19340 7200
rect 19392 7188 19398 7200
rect 21174 7188 21180 7200
rect 19392 7160 21180 7188
rect 19392 7148 19398 7160
rect 21174 7148 21180 7160
rect 21232 7148 21238 7200
rect 21818 7148 21824 7200
rect 21876 7188 21882 7200
rect 22465 7191 22523 7197
rect 22465 7188 22477 7191
rect 21876 7160 22477 7188
rect 21876 7148 21882 7160
rect 22465 7157 22477 7160
rect 22511 7157 22523 7191
rect 22465 7151 22523 7157
rect 22833 7191 22891 7197
rect 22833 7157 22845 7191
rect 22879 7188 22891 7191
rect 23293 7191 23351 7197
rect 23293 7188 23305 7191
rect 22879 7160 23305 7188
rect 22879 7157 22891 7160
rect 22833 7151 22891 7157
rect 23293 7157 23305 7160
rect 23339 7157 23351 7191
rect 23293 7151 23351 7157
rect 25590 7148 25596 7200
rect 25648 7188 25654 7200
rect 25777 7191 25835 7197
rect 25777 7188 25789 7191
rect 25648 7160 25789 7188
rect 25648 7148 25654 7160
rect 25777 7157 25789 7160
rect 25823 7157 25835 7191
rect 27062 7188 27068 7200
rect 27023 7160 27068 7188
rect 25777 7151 25835 7157
rect 27062 7148 27068 7160
rect 27120 7148 27126 7200
rect 27890 7148 27896 7200
rect 27948 7188 27954 7200
rect 27948 7160 27993 7188
rect 27948 7148 27954 7160
rect 1104 7098 29440 7120
rect 1104 7046 4492 7098
rect 4544 7046 4556 7098
rect 4608 7046 4620 7098
rect 4672 7046 4684 7098
rect 4736 7046 4748 7098
rect 4800 7046 11576 7098
rect 11628 7046 11640 7098
rect 11692 7046 11704 7098
rect 11756 7046 11768 7098
rect 11820 7046 11832 7098
rect 11884 7046 18660 7098
rect 18712 7046 18724 7098
rect 18776 7046 18788 7098
rect 18840 7046 18852 7098
rect 18904 7046 18916 7098
rect 18968 7046 25744 7098
rect 25796 7046 25808 7098
rect 25860 7046 25872 7098
rect 25924 7046 25936 7098
rect 25988 7046 26000 7098
rect 26052 7046 29440 7098
rect 1104 7024 29440 7046
rect 4341 6987 4399 6993
rect 4341 6953 4353 6987
rect 4387 6953 4399 6987
rect 4890 6984 4896 6996
rect 4851 6956 4896 6984
rect 4341 6947 4399 6953
rect 4356 6916 4384 6947
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 9582 6984 9588 6996
rect 9272 6956 9588 6984
rect 9272 6944 9278 6956
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 11422 6944 11428 6996
rect 11480 6984 11486 6996
rect 11793 6987 11851 6993
rect 11793 6984 11805 6987
rect 11480 6956 11805 6984
rect 11480 6944 11486 6956
rect 11793 6953 11805 6956
rect 11839 6953 11851 6987
rect 11793 6947 11851 6953
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 13173 6987 13231 6993
rect 13173 6984 13185 6987
rect 12952 6956 13185 6984
rect 12952 6944 12958 6956
rect 13173 6953 13185 6956
rect 13219 6953 13231 6987
rect 13173 6947 13231 6953
rect 13906 6944 13912 6996
rect 13964 6984 13970 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 13964 6956 14105 6984
rect 13964 6944 13970 6956
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 9398 6916 9404 6928
rect 4356 6888 5028 6916
rect 9359 6888 9404 6916
rect 4246 6848 4252 6860
rect 4207 6820 4252 6848
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 4801 6783 4859 6789
rect 4801 6780 4813 6783
rect 4387 6752 4813 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4801 6749 4813 6752
rect 4847 6780 4859 6783
rect 4890 6780 4896 6792
rect 4847 6752 4896 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 5000 6789 5028 6888
rect 9398 6876 9404 6888
rect 9456 6876 9462 6928
rect 9766 6916 9772 6928
rect 9508 6888 9772 6916
rect 8386 6848 8392 6860
rect 7024 6820 8392 6848
rect 7024 6792 7052 6820
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 9508 6857 9536 6888
rect 9766 6876 9772 6888
rect 9824 6916 9830 6928
rect 10505 6919 10563 6925
rect 10505 6916 10517 6919
rect 9824 6888 10517 6916
rect 9824 6876 9830 6888
rect 10505 6885 10517 6888
rect 10551 6916 10563 6919
rect 10594 6916 10600 6928
rect 10551 6888 10600 6916
rect 10551 6885 10563 6888
rect 10505 6879 10563 6885
rect 10594 6876 10600 6888
rect 10652 6876 10658 6928
rect 12713 6919 12771 6925
rect 12713 6885 12725 6919
rect 12759 6885 12771 6919
rect 14108 6916 14136 6947
rect 14366 6944 14372 6996
rect 14424 6984 14430 6996
rect 14461 6987 14519 6993
rect 14461 6984 14473 6987
rect 14424 6956 14473 6984
rect 14424 6944 14430 6956
rect 14461 6953 14473 6956
rect 14507 6953 14519 6987
rect 14461 6947 14519 6953
rect 16853 6987 16911 6993
rect 16853 6953 16865 6987
rect 16899 6984 16911 6987
rect 17218 6984 17224 6996
rect 16899 6956 17224 6984
rect 16899 6953 16911 6956
rect 16853 6947 16911 6953
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 18693 6987 18751 6993
rect 18693 6984 18705 6987
rect 18564 6956 18705 6984
rect 18564 6944 18570 6956
rect 18693 6953 18705 6956
rect 18739 6953 18751 6987
rect 18693 6947 18751 6953
rect 21174 6944 21180 6996
rect 21232 6984 21238 6996
rect 22097 6987 22155 6993
rect 22097 6984 22109 6987
rect 21232 6956 22109 6984
rect 21232 6944 21238 6956
rect 22097 6953 22109 6956
rect 22143 6953 22155 6987
rect 22097 6947 22155 6953
rect 23477 6987 23535 6993
rect 23477 6953 23489 6987
rect 23523 6984 23535 6987
rect 23566 6984 23572 6996
rect 23523 6956 23572 6984
rect 23523 6953 23535 6956
rect 23477 6947 23535 6953
rect 14108 6888 14412 6916
rect 12713 6879 12771 6885
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 9600 6820 11652 6848
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6780 5043 6783
rect 5258 6780 5264 6792
rect 5031 6752 5264 6780
rect 5031 6749 5043 6752
rect 4985 6743 5043 6749
rect 5258 6740 5264 6752
rect 5316 6780 5322 6792
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5316 6752 5825 6780
rect 5316 6740 5322 6752
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 5902 6740 5908 6792
rect 5960 6780 5966 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5960 6752 6009 6780
rect 5960 6740 5966 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 7006 6780 7012 6792
rect 6967 6752 7012 6780
rect 6273 6743 6331 6749
rect 6288 6712 6316 6743
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 7190 6780 7196 6792
rect 7151 6752 7196 6780
rect 7190 6740 7196 6752
rect 7248 6780 7254 6792
rect 7653 6783 7711 6789
rect 7653 6780 7665 6783
rect 7248 6752 7665 6780
rect 7248 6740 7254 6752
rect 7653 6749 7665 6752
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9600 6789 9628 6820
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 9272 6752 9321 6780
rect 9272 6740 9278 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9574 6783 9632 6789
rect 9574 6749 9586 6783
rect 9620 6749 9632 6783
rect 9574 6743 9632 6749
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 9732 6752 10333 6780
rect 9732 6740 9738 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 7101 6715 7159 6721
rect 7101 6712 7113 6715
rect 6288 6684 7113 6712
rect 7101 6681 7113 6684
rect 7147 6681 7159 6715
rect 7101 6675 7159 6681
rect 8389 6715 8447 6721
rect 8389 6681 8401 6715
rect 8435 6712 8447 6715
rect 8478 6712 8484 6724
rect 8435 6684 8484 6712
rect 8435 6681 8447 6684
rect 8389 6675 8447 6681
rect 8478 6672 8484 6684
rect 8536 6672 8542 6724
rect 9125 6715 9183 6721
rect 9125 6681 9137 6715
rect 9171 6712 9183 6715
rect 9858 6712 9864 6724
rect 9171 6684 9864 6712
rect 9171 6681 9183 6684
rect 9125 6675 9183 6681
rect 9858 6672 9864 6684
rect 9916 6672 9922 6724
rect 10428 6712 10456 6743
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 10612 6789 10640 6820
rect 10597 6783 10655 6789
rect 10597 6780 10609 6783
rect 10560 6752 10609 6780
rect 10560 6740 10566 6752
rect 10597 6749 10609 6752
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 11238 6780 11244 6792
rect 10836 6752 10881 6780
rect 11199 6752 11244 6780
rect 10836 6740 10842 6752
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11624 6789 11652 6820
rect 11517 6783 11575 6789
rect 11388 6752 11433 6780
rect 11388 6740 11394 6752
rect 11517 6749 11529 6783
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 9968 6684 10456 6712
rect 11532 6712 11560 6743
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 12728 6780 12756 6879
rect 14274 6848 14280 6860
rect 14108 6820 14280 6848
rect 13173 6783 13231 6789
rect 13173 6780 13185 6783
rect 12492 6752 12537 6780
rect 12728 6752 13185 6780
rect 12492 6740 12498 6752
rect 13173 6749 13185 6752
rect 13219 6749 13231 6783
rect 13173 6743 13231 6749
rect 13262 6740 13268 6792
rect 13320 6780 13326 6792
rect 14108 6789 14136 6820
rect 14274 6808 14280 6820
rect 14332 6808 14338 6860
rect 14384 6848 14412 6888
rect 15838 6876 15844 6928
rect 15896 6916 15902 6928
rect 15933 6919 15991 6925
rect 15933 6916 15945 6919
rect 15896 6888 15945 6916
rect 15896 6876 15902 6888
rect 15933 6885 15945 6888
rect 15979 6885 15991 6919
rect 17770 6916 17776 6928
rect 15933 6879 15991 6885
rect 16868 6888 17776 6916
rect 16868 6848 16896 6888
rect 17770 6876 17776 6888
rect 17828 6876 17834 6928
rect 18340 6888 19334 6916
rect 14384 6820 15884 6848
rect 13357 6783 13415 6789
rect 13357 6780 13369 6783
rect 13320 6752 13369 6780
rect 13320 6740 13326 6752
rect 13357 6749 13369 6752
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 14182 6740 14188 6792
rect 14240 6780 14246 6792
rect 15654 6780 15660 6792
rect 14240 6752 15660 6780
rect 14240 6740 14246 6752
rect 15654 6740 15660 6752
rect 15712 6780 15718 6792
rect 15856 6789 15884 6820
rect 16132 6820 16896 6848
rect 16945 6851 17003 6857
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 15712 6752 15761 6780
rect 15712 6740 15718 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 16022 6780 16028 6792
rect 15983 6752 16028 6780
rect 15841 6743 15899 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 12713 6715 12771 6721
rect 12713 6712 12725 6715
rect 11532 6684 12725 6712
rect 3970 6644 3976 6656
rect 3931 6616 3976 6644
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5350 6644 5356 6656
rect 5215 6616 5356 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 6178 6644 6184 6656
rect 6139 6616 6184 6644
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 9968 6644 9996 6684
rect 12713 6681 12725 6684
rect 12759 6712 12771 6715
rect 13814 6712 13820 6724
rect 12759 6684 13820 6712
rect 12759 6681 12771 6684
rect 12713 6675 12771 6681
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 15565 6715 15623 6721
rect 15565 6681 15577 6715
rect 15611 6712 15623 6715
rect 16132 6712 16160 6820
rect 16945 6817 16957 6851
rect 16991 6848 17003 6851
rect 17494 6848 17500 6860
rect 16991 6820 17500 6848
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16669 6783 16727 6789
rect 16669 6780 16681 6783
rect 16255 6752 16681 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 16669 6749 16681 6752
rect 16715 6749 16727 6783
rect 16669 6743 16727 6749
rect 15611 6684 16160 6712
rect 16684 6712 16712 6743
rect 16758 6740 16764 6792
rect 16816 6780 16822 6792
rect 18230 6780 18236 6792
rect 16816 6752 16861 6780
rect 18143 6752 18236 6780
rect 16816 6740 16822 6752
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 18340 6789 18368 6888
rect 18506 6808 18512 6860
rect 18564 6848 18570 6860
rect 19306 6848 19334 6888
rect 19518 6848 19524 6860
rect 18564 6820 18736 6848
rect 19306 6820 19524 6848
rect 18564 6808 18570 6820
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18598 6780 18604 6792
rect 18559 6752 18604 6780
rect 18325 6743 18383 6749
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 18708 6789 18736 6820
rect 19518 6808 19524 6820
rect 19576 6808 19582 6860
rect 20714 6848 20720 6860
rect 20675 6820 20720 6848
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 22112 6848 22140 6947
rect 22649 6851 22707 6857
rect 22649 6848 22661 6851
rect 22112 6820 22661 6848
rect 22649 6817 22661 6820
rect 22695 6817 22707 6851
rect 22649 6811 22707 6817
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6780 18751 6783
rect 19242 6780 19248 6792
rect 18739 6752 19248 6780
rect 18739 6749 18751 6752
rect 18693 6743 18751 6749
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19610 6780 19616 6792
rect 19392 6752 19437 6780
rect 19571 6752 19616 6780
rect 19392 6740 19398 6752
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 19751 6783 19809 6789
rect 19751 6749 19763 6783
rect 19797 6749 19809 6783
rect 20438 6780 20444 6792
rect 20399 6752 20444 6780
rect 19751 6743 19809 6749
rect 17954 6712 17960 6724
rect 16684 6684 17960 6712
rect 15611 6681 15623 6684
rect 15565 6675 15623 6681
rect 17954 6672 17960 6684
rect 18012 6672 18018 6724
rect 10134 6644 10140 6656
rect 9456 6616 9996 6644
rect 10095 6616 10140 6644
rect 9456 6604 9462 6616
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 12529 6647 12587 6653
rect 12529 6644 12541 6647
rect 12400 6616 12541 6644
rect 12400 6604 12406 6616
rect 12529 6613 12541 6616
rect 12575 6613 12587 6647
rect 12529 6607 12587 6613
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 15013 6647 15071 6653
rect 15013 6644 15025 6647
rect 14792 6616 15025 6644
rect 14792 6604 14798 6616
rect 15013 6613 15025 6616
rect 15059 6644 15071 6647
rect 17494 6644 17500 6656
rect 15059 6616 17500 6644
rect 15059 6613 15071 6616
rect 15013 6607 15071 6613
rect 17494 6604 17500 6616
rect 17552 6604 17558 6656
rect 18248 6644 18276 6740
rect 18417 6715 18475 6721
rect 18417 6681 18429 6715
rect 18463 6712 18475 6715
rect 19518 6712 19524 6724
rect 18463 6684 19524 6712
rect 18463 6681 18475 6684
rect 18417 6675 18475 6681
rect 19518 6672 19524 6684
rect 19576 6672 19582 6724
rect 19764 6644 19792 6743
rect 20438 6740 20444 6752
rect 20496 6740 20502 6792
rect 20530 6740 20536 6792
rect 20588 6780 20594 6792
rect 20588 6752 20633 6780
rect 20588 6740 20594 6752
rect 20898 6740 20904 6792
rect 20956 6780 20962 6792
rect 22002 6780 22008 6792
rect 20956 6752 22008 6780
rect 20956 6740 20962 6752
rect 22002 6740 22008 6752
rect 22060 6740 22066 6792
rect 22189 6783 22247 6789
rect 22189 6749 22201 6783
rect 22235 6780 22247 6783
rect 22738 6780 22744 6792
rect 22235 6752 22744 6780
rect 22235 6749 22247 6752
rect 22189 6743 22247 6749
rect 22738 6740 22744 6752
rect 22796 6740 22802 6792
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6780 22891 6783
rect 23492 6780 23520 6947
rect 23566 6944 23572 6956
rect 23624 6944 23630 6996
rect 25590 6944 25596 6996
rect 25648 6984 25654 6996
rect 25685 6987 25743 6993
rect 25685 6984 25697 6987
rect 25648 6956 25697 6984
rect 25648 6944 25654 6956
rect 25685 6953 25697 6956
rect 25731 6953 25743 6987
rect 25685 6947 25743 6953
rect 27062 6944 27068 6996
rect 27120 6984 27126 6996
rect 27341 6987 27399 6993
rect 27341 6984 27353 6987
rect 27120 6956 27353 6984
rect 27120 6944 27126 6956
rect 27341 6953 27353 6956
rect 27387 6953 27399 6987
rect 27341 6947 27399 6953
rect 27801 6987 27859 6993
rect 27801 6953 27813 6987
rect 27847 6984 27859 6987
rect 27890 6984 27896 6996
rect 27847 6956 27896 6984
rect 27847 6953 27859 6956
rect 27801 6947 27859 6953
rect 27890 6944 27896 6956
rect 27948 6944 27954 6996
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6848 25191 6851
rect 26789 6851 26847 6857
rect 26789 6848 26801 6851
rect 25179 6820 26801 6848
rect 25179 6817 25191 6820
rect 25133 6811 25191 6817
rect 26789 6817 26801 6820
rect 26835 6848 26847 6851
rect 27522 6848 27528 6860
rect 26835 6820 27528 6848
rect 26835 6817 26847 6820
rect 26789 6811 26847 6817
rect 27522 6808 27528 6820
rect 27580 6808 27586 6860
rect 27614 6808 27620 6860
rect 27672 6848 27678 6860
rect 28074 6848 28080 6860
rect 27672 6820 28080 6848
rect 27672 6808 27678 6820
rect 28074 6808 28080 6820
rect 28132 6848 28138 6860
rect 28261 6851 28319 6857
rect 28261 6848 28273 6851
rect 28132 6820 28273 6848
rect 28132 6808 28138 6820
rect 28261 6817 28273 6820
rect 28307 6817 28319 6851
rect 28261 6811 28319 6817
rect 28350 6808 28356 6860
rect 28408 6848 28414 6860
rect 28408 6820 28453 6848
rect 28408 6808 28414 6820
rect 25317 6783 25375 6789
rect 22879 6752 23520 6780
rect 23584 6780 23888 6782
rect 25317 6780 25329 6783
rect 23584 6754 25329 6780
rect 22879 6749 22891 6752
rect 22833 6743 22891 6749
rect 20717 6715 20775 6721
rect 20717 6681 20729 6715
rect 20763 6712 20775 6715
rect 21266 6712 21272 6724
rect 20763 6684 21272 6712
rect 20763 6681 20775 6684
rect 20717 6675 20775 6681
rect 21266 6672 21272 6684
rect 21324 6672 21330 6724
rect 21358 6672 21364 6724
rect 21416 6712 21422 6724
rect 23584 6712 23612 6754
rect 23860 6752 25329 6754
rect 25317 6749 25329 6752
rect 25363 6780 25375 6783
rect 28442 6780 28448 6792
rect 25363 6752 28448 6780
rect 25363 6749 25375 6752
rect 25317 6743 25375 6749
rect 28442 6740 28448 6752
rect 28500 6740 28506 6792
rect 21416 6684 23612 6712
rect 21416 6672 21422 6684
rect 23658 6672 23664 6724
rect 23716 6712 23722 6724
rect 23716 6684 23761 6712
rect 23716 6672 23722 6684
rect 23842 6672 23848 6724
rect 23900 6712 23906 6724
rect 26881 6715 26939 6721
rect 23900 6684 23945 6712
rect 23900 6672 23906 6684
rect 26881 6681 26893 6715
rect 26927 6712 26939 6715
rect 28166 6712 28172 6724
rect 26927 6684 27200 6712
rect 28127 6684 28172 6712
rect 26927 6681 26939 6684
rect 26881 6675 26939 6681
rect 18248 6616 19792 6644
rect 19889 6647 19947 6653
rect 19889 6613 19901 6647
rect 19935 6644 19947 6647
rect 20806 6644 20812 6656
rect 19935 6616 20812 6644
rect 19935 6613 19947 6616
rect 19889 6607 19947 6613
rect 20806 6604 20812 6616
rect 20864 6604 20870 6656
rect 21082 6604 21088 6656
rect 21140 6644 21146 6656
rect 21177 6647 21235 6653
rect 21177 6644 21189 6647
rect 21140 6616 21189 6644
rect 21140 6604 21146 6616
rect 21177 6613 21189 6616
rect 21223 6613 21235 6647
rect 21177 6607 21235 6613
rect 22738 6604 22744 6656
rect 22796 6644 22802 6656
rect 23017 6647 23075 6653
rect 23017 6644 23029 6647
rect 22796 6616 23029 6644
rect 22796 6604 22802 6616
rect 23017 6613 23029 6616
rect 23063 6613 23075 6647
rect 23676 6644 23704 6672
rect 24397 6647 24455 6653
rect 24397 6644 24409 6647
rect 23676 6616 24409 6644
rect 23017 6607 23075 6613
rect 24397 6613 24409 6616
rect 24443 6613 24455 6647
rect 25222 6644 25228 6656
rect 25183 6616 25228 6644
rect 24397 6607 24455 6613
rect 25222 6604 25228 6616
rect 25280 6604 25286 6656
rect 26970 6604 26976 6656
rect 27028 6644 27034 6656
rect 27172 6644 27200 6684
rect 28166 6672 28172 6684
rect 28224 6672 28230 6724
rect 27706 6644 27712 6656
rect 27028 6616 27073 6644
rect 27172 6616 27712 6644
rect 27028 6604 27034 6616
rect 27706 6604 27712 6616
rect 27764 6644 27770 6656
rect 28258 6644 28264 6656
rect 27764 6616 28264 6644
rect 27764 6604 27770 6616
rect 28258 6604 28264 6616
rect 28316 6604 28322 6656
rect 1104 6554 29600 6576
rect 1104 6502 8034 6554
rect 8086 6502 8098 6554
rect 8150 6502 8162 6554
rect 8214 6502 8226 6554
rect 8278 6502 8290 6554
rect 8342 6502 15118 6554
rect 15170 6502 15182 6554
rect 15234 6502 15246 6554
rect 15298 6502 15310 6554
rect 15362 6502 15374 6554
rect 15426 6502 22202 6554
rect 22254 6502 22266 6554
rect 22318 6502 22330 6554
rect 22382 6502 22394 6554
rect 22446 6502 22458 6554
rect 22510 6502 29286 6554
rect 29338 6502 29350 6554
rect 29402 6502 29414 6554
rect 29466 6502 29478 6554
rect 29530 6502 29542 6554
rect 29594 6502 29600 6554
rect 1104 6480 29600 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 5500 6412 5580 6440
rect 5500 6400 5506 6412
rect 3970 6332 3976 6384
rect 4028 6372 4034 6384
rect 4028 6344 5488 6372
rect 4028 6332 4034 6344
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6264 1458 6316
rect 5166 6304 5172 6316
rect 5127 6276 5172 6304
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 5350 6304 5356 6316
rect 5311 6276 5356 6304
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5460 6313 5488 6344
rect 5552 6313 5580 6412
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6546 6440 6552 6452
rect 5960 6412 6552 6440
rect 5960 6400 5966 6412
rect 6546 6400 6552 6412
rect 6604 6440 6610 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 6604 6412 6837 6440
rect 6604 6400 6610 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 8665 6443 8723 6449
rect 8665 6409 8677 6443
rect 8711 6440 8723 6443
rect 9214 6440 9220 6452
rect 8711 6412 9220 6440
rect 8711 6409 8723 6412
rect 8665 6403 8723 6409
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 11330 6440 11336 6452
rect 10643 6412 11336 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 11885 6443 11943 6449
rect 11885 6409 11897 6443
rect 11931 6440 11943 6443
rect 12342 6440 12348 6452
rect 11931 6412 12348 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 12621 6443 12679 6449
rect 12621 6409 12633 6443
rect 12667 6440 12679 6443
rect 12710 6440 12716 6452
rect 12667 6412 12716 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 13262 6440 13268 6452
rect 13223 6412 13268 6440
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 14090 6440 14096 6452
rect 14051 6412 14096 6440
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 14550 6440 14556 6452
rect 14511 6412 14556 6440
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 15841 6443 15899 6449
rect 15841 6409 15853 6443
rect 15887 6440 15899 6443
rect 16758 6440 16764 6452
rect 15887 6412 16764 6440
rect 15887 6409 15899 6412
rect 15841 6403 15899 6409
rect 16758 6400 16764 6412
rect 16816 6400 16822 6452
rect 18414 6440 18420 6452
rect 18375 6412 18420 6440
rect 18414 6400 18420 6412
rect 18472 6400 18478 6452
rect 18598 6400 18604 6452
rect 18656 6440 18662 6452
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 18656 6412 19073 6440
rect 18656 6400 18662 6412
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 19061 6403 19119 6409
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 19613 6443 19671 6449
rect 19613 6440 19625 6443
rect 19300 6412 19625 6440
rect 19300 6400 19306 6412
rect 19613 6409 19625 6412
rect 19659 6409 19671 6443
rect 19613 6403 19671 6409
rect 19886 6400 19892 6452
rect 19944 6440 19950 6452
rect 20530 6440 20536 6452
rect 19944 6412 20536 6440
rect 19944 6400 19950 6412
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 22002 6400 22008 6452
rect 22060 6440 22066 6452
rect 23201 6443 23259 6449
rect 23201 6440 23213 6443
rect 22060 6412 23213 6440
rect 22060 6400 22066 6412
rect 23201 6409 23213 6412
rect 23247 6440 23259 6443
rect 23842 6440 23848 6452
rect 23247 6412 23848 6440
rect 23247 6409 23259 6412
rect 23201 6403 23259 6409
rect 23842 6400 23848 6412
rect 23900 6440 23906 6452
rect 24121 6443 24179 6449
rect 24121 6440 24133 6443
rect 23900 6412 24133 6440
rect 23900 6400 23906 6412
rect 24121 6409 24133 6412
rect 24167 6409 24179 6443
rect 24121 6403 24179 6409
rect 24210 6400 24216 6452
rect 24268 6440 24274 6452
rect 26421 6443 26479 6449
rect 26421 6440 26433 6443
rect 24268 6412 26433 6440
rect 24268 6400 24274 6412
rect 26421 6409 26433 6412
rect 26467 6440 26479 6443
rect 26970 6440 26976 6452
rect 26467 6412 26976 6440
rect 26467 6409 26479 6412
rect 26421 6403 26479 6409
rect 26970 6400 26976 6412
rect 27028 6400 27034 6452
rect 27065 6443 27123 6449
rect 27065 6409 27077 6443
rect 27111 6440 27123 6443
rect 27706 6440 27712 6452
rect 27111 6412 27712 6440
rect 27111 6409 27123 6412
rect 27065 6403 27123 6409
rect 27706 6400 27712 6412
rect 27764 6400 27770 6452
rect 28074 6440 28080 6452
rect 28035 6412 28080 6440
rect 28074 6400 28080 6412
rect 28132 6400 28138 6452
rect 6178 6332 6184 6384
rect 6236 6372 6242 6384
rect 6730 6372 6736 6384
rect 6236 6344 6736 6372
rect 6236 6332 6242 6344
rect 6730 6332 6736 6344
rect 6788 6372 6794 6384
rect 9585 6375 9643 6381
rect 6788 6344 7972 6372
rect 6788 6332 6794 6344
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 7006 6304 7012 6316
rect 6967 6276 7012 6304
rect 5537 6267 5595 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7190 6304 7196 6316
rect 7151 6276 7196 6304
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 7944 6313 7972 6344
rect 9585 6341 9597 6375
rect 9631 6372 9643 6375
rect 10229 6375 10287 6381
rect 10229 6372 10241 6375
rect 9631 6344 10241 6372
rect 9631 6341 9643 6344
rect 9585 6335 9643 6341
rect 10229 6341 10241 6344
rect 10275 6372 10287 6375
rect 10962 6372 10968 6384
rect 10275 6344 10968 6372
rect 10275 6341 10287 6344
rect 10229 6335 10287 6341
rect 10962 6332 10968 6344
rect 11020 6332 11026 6384
rect 13280 6372 13308 6400
rect 14568 6372 14596 6400
rect 15470 6372 15476 6384
rect 12728 6344 13308 6372
rect 13372 6344 14596 6372
rect 15383 6344 15476 6372
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8536 6276 8861 6304
rect 8536 6264 8542 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 9030 6304 9036 6316
rect 8991 6276 9036 6304
rect 8849 6267 8907 6273
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 9364 6276 10057 6304
rect 9364 6264 9370 6276
rect 10045 6273 10057 6276
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 10870 6304 10876 6316
rect 10459 6276 10876 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6236 7343 6239
rect 7837 6239 7895 6245
rect 7837 6236 7849 6239
rect 7331 6208 7849 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 7837 6205 7849 6208
rect 7883 6205 7895 6239
rect 10336 6236 10364 6267
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 12728 6313 12756 6344
rect 12529 6307 12587 6313
rect 12529 6304 12541 6307
rect 12492 6276 12541 6304
rect 12492 6264 12498 6276
rect 12529 6273 12541 6276
rect 12575 6273 12587 6307
rect 12529 6267 12587 6273
rect 12713 6307 12771 6313
rect 12713 6273 12725 6307
rect 12759 6273 12771 6307
rect 13170 6304 13176 6316
rect 13131 6276 13176 6304
rect 12713 6267 12771 6273
rect 10594 6236 10600 6248
rect 10336 6208 10600 6236
rect 7837 6199 7895 6205
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 10778 6196 10784 6248
rect 10836 6236 10842 6248
rect 10962 6236 10968 6248
rect 10836 6208 10968 6236
rect 10836 6196 10842 6208
rect 10962 6196 10968 6208
rect 11020 6236 11026 6248
rect 12544 6236 12572 6267
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 13262 6264 13268 6316
rect 13320 6304 13326 6316
rect 13372 6313 13400 6344
rect 13357 6307 13415 6313
rect 13357 6304 13369 6307
rect 13320 6276 13369 6304
rect 13320 6264 13326 6276
rect 13357 6273 13369 6276
rect 13403 6273 13415 6307
rect 13357 6267 13415 6273
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6304 13875 6307
rect 14182 6304 14188 6316
rect 13863 6276 14188 6304
rect 13863 6273 13875 6276
rect 13817 6267 13875 6273
rect 13832 6236 13860 6267
rect 14182 6264 14188 6276
rect 14240 6264 14246 6316
rect 15396 6313 15424 6344
rect 15470 6332 15476 6344
rect 15528 6372 15534 6384
rect 16022 6372 16028 6384
rect 15528 6344 16028 6372
rect 15528 6332 15534 6344
rect 16022 6332 16028 6344
rect 16080 6372 16086 6384
rect 16669 6375 16727 6381
rect 16669 6372 16681 6375
rect 16080 6344 16681 6372
rect 16080 6332 16086 6344
rect 16669 6341 16681 6344
rect 16715 6341 16727 6375
rect 17957 6375 18015 6381
rect 17957 6372 17969 6375
rect 16669 6335 16727 6341
rect 16868 6344 17969 6372
rect 16868 6316 16896 6344
rect 17957 6341 17969 6344
rect 18003 6372 18015 6375
rect 18046 6372 18052 6384
rect 18003 6344 18052 6372
rect 18003 6341 18015 6344
rect 17957 6335 18015 6341
rect 18046 6332 18052 6344
rect 18104 6332 18110 6384
rect 19334 6372 19340 6384
rect 19168 6344 19340 6372
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6273 15439 6307
rect 15654 6304 15660 6316
rect 15615 6276 15660 6304
rect 15381 6267 15439 6273
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 16850 6304 16856 6316
rect 16811 6276 16856 6304
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 17034 6304 17040 6316
rect 16995 6276 17040 6304
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6304 18291 6307
rect 18322 6304 18328 6316
rect 18279 6276 18328 6304
rect 18279 6273 18291 6276
rect 18233 6267 18291 6273
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 19168 6313 19196 6344
rect 19334 6332 19340 6344
rect 19392 6372 19398 6384
rect 19392 6344 20484 6372
rect 19392 6332 19398 6344
rect 20456 6316 20484 6344
rect 20714 6332 20720 6384
rect 20772 6372 20778 6384
rect 22649 6375 22707 6381
rect 20772 6344 22232 6372
rect 20772 6332 20778 6344
rect 19153 6307 19211 6313
rect 19153 6273 19165 6307
rect 19199 6273 19211 6307
rect 19153 6267 19211 6273
rect 20070 6264 20076 6316
rect 20128 6304 20134 6316
rect 20349 6307 20407 6313
rect 20349 6304 20361 6307
rect 20128 6276 20361 6304
rect 20128 6264 20134 6276
rect 20349 6273 20361 6276
rect 20395 6273 20407 6307
rect 20349 6267 20407 6273
rect 11020 6208 12434 6236
rect 12544 6208 13860 6236
rect 14093 6239 14151 6245
rect 11020 6196 11026 6208
rect 5813 6171 5871 6177
rect 5813 6137 5825 6171
rect 5859 6168 5871 6171
rect 5859 6140 10088 6168
rect 5859 6137 5871 6140
rect 5813 6131 5871 6137
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 4396 6072 4629 6100
rect 4396 6060 4402 6072
rect 4617 6069 4629 6072
rect 4663 6100 4675 6103
rect 6178 6100 6184 6112
rect 4663 6072 6184 6100
rect 4663 6069 4675 6072
rect 4617 6063 4675 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 10060 6100 10088 6140
rect 10134 6128 10140 6180
rect 10192 6168 10198 6180
rect 12406 6168 12434 6208
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 14274 6236 14280 6248
rect 14139 6208 14280 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 15473 6239 15531 6245
rect 15473 6205 15485 6239
rect 15519 6236 15531 6239
rect 15838 6236 15844 6248
rect 15519 6208 15844 6236
rect 15519 6205 15531 6208
rect 15473 6199 15531 6205
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 18141 6239 18199 6245
rect 18141 6205 18153 6239
rect 18187 6236 18199 6239
rect 19058 6236 19064 6248
rect 18187 6208 19064 6236
rect 18187 6205 18199 6208
rect 18141 6199 18199 6205
rect 19058 6196 19064 6208
rect 19116 6196 19122 6248
rect 19978 6196 19984 6248
rect 20036 6236 20042 6248
rect 20165 6239 20223 6245
rect 20165 6236 20177 6239
rect 20036 6208 20177 6236
rect 20036 6196 20042 6208
rect 20165 6205 20177 6208
rect 20211 6236 20223 6239
rect 20364 6236 20392 6267
rect 20438 6264 20444 6316
rect 20496 6304 20502 6316
rect 22204 6313 22232 6344
rect 22649 6341 22661 6375
rect 22695 6372 22707 6375
rect 22830 6372 22836 6384
rect 22695 6344 22836 6372
rect 22695 6341 22707 6344
rect 22649 6335 22707 6341
rect 22830 6332 22836 6344
rect 22888 6372 22894 6384
rect 23658 6372 23664 6384
rect 22888 6344 23664 6372
rect 22888 6332 22894 6344
rect 23658 6332 23664 6344
rect 23716 6332 23722 6384
rect 25869 6375 25927 6381
rect 25869 6341 25881 6375
rect 25915 6372 25927 6375
rect 27614 6372 27620 6384
rect 25915 6344 27620 6372
rect 25915 6341 25927 6344
rect 25869 6335 25927 6341
rect 27614 6332 27620 6344
rect 27672 6372 27678 6384
rect 28350 6372 28356 6384
rect 27672 6344 28356 6372
rect 27672 6332 27678 6344
rect 28350 6332 28356 6344
rect 28408 6372 28414 6384
rect 28629 6375 28687 6381
rect 28629 6372 28641 6375
rect 28408 6344 28641 6372
rect 28408 6332 28414 6344
rect 28629 6341 28641 6344
rect 28675 6341 28687 6375
rect 28629 6335 28687 6341
rect 20533 6307 20591 6313
rect 20533 6304 20545 6307
rect 20496 6276 20545 6304
rect 20496 6264 20502 6276
rect 20533 6273 20545 6276
rect 20579 6304 20591 6307
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 20579 6276 22017 6304
rect 20579 6273 20591 6276
rect 20533 6267 20591 6273
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6304 22247 6307
rect 22738 6304 22744 6316
rect 22235 6276 22744 6304
rect 22235 6273 22247 6276
rect 22189 6267 22247 6273
rect 22738 6264 22744 6276
rect 22796 6264 22802 6316
rect 20806 6236 20812 6248
rect 20211 6208 20300 6236
rect 20364 6208 20812 6236
rect 20211 6205 20223 6208
rect 20165 6199 20223 6205
rect 12710 6168 12716 6180
rect 10192 6140 11928 6168
rect 12406 6140 12716 6168
rect 10192 6128 10198 6140
rect 11422 6100 11428 6112
rect 10060 6072 11428 6100
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 11900 6100 11928 6140
rect 12710 6128 12716 6140
rect 12768 6128 12774 6180
rect 15565 6171 15623 6177
rect 15565 6168 15577 6171
rect 13924 6140 15577 6168
rect 13924 6112 13952 6140
rect 15565 6137 15577 6140
rect 15611 6137 15623 6171
rect 15565 6131 15623 6137
rect 17770 6128 17776 6180
rect 17828 6168 17834 6180
rect 19886 6168 19892 6180
rect 17828 6140 19892 6168
rect 17828 6128 17834 6140
rect 19886 6128 19892 6140
rect 19944 6128 19950 6180
rect 20272 6168 20300 6208
rect 20806 6196 20812 6208
rect 20864 6236 20870 6248
rect 21358 6236 21364 6248
rect 20864 6208 21364 6236
rect 20864 6196 20870 6208
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 20272 6140 20392 6168
rect 13906 6100 13912 6112
rect 11900 6072 13912 6100
rect 13906 6060 13912 6072
rect 13964 6060 13970 6112
rect 18233 6103 18291 6109
rect 18233 6069 18245 6103
rect 18279 6100 18291 6103
rect 19242 6100 19248 6112
rect 18279 6072 19248 6100
rect 18279 6069 18291 6072
rect 18233 6063 18291 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 20364 6100 20392 6140
rect 20530 6128 20536 6180
rect 20588 6168 20594 6180
rect 20588 6140 22048 6168
rect 20588 6128 20594 6140
rect 21082 6100 21088 6112
rect 20364 6072 21088 6100
rect 21082 6060 21088 6072
rect 21140 6060 21146 6112
rect 21174 6060 21180 6112
rect 21232 6100 21238 6112
rect 22020 6109 22048 6140
rect 22462 6128 22468 6180
rect 22520 6168 22526 6180
rect 22922 6168 22928 6180
rect 22520 6140 22928 6168
rect 22520 6128 22526 6140
rect 22922 6128 22928 6140
rect 22980 6168 22986 6180
rect 24857 6171 24915 6177
rect 24857 6168 24869 6171
rect 22980 6140 24869 6168
rect 22980 6128 22986 6140
rect 24857 6137 24869 6140
rect 24903 6168 24915 6171
rect 25222 6168 25228 6180
rect 24903 6140 25228 6168
rect 24903 6137 24915 6140
rect 24857 6131 24915 6137
rect 25222 6128 25228 6140
rect 25280 6128 25286 6180
rect 21821 6103 21879 6109
rect 21821 6100 21833 6103
rect 21232 6072 21833 6100
rect 21232 6060 21238 6072
rect 21821 6069 21833 6072
rect 21867 6069 21879 6103
rect 21821 6063 21879 6069
rect 22005 6103 22063 6109
rect 22005 6069 22017 6103
rect 22051 6069 22063 6103
rect 22005 6063 22063 6069
rect 1104 6010 29440 6032
rect 1104 5958 4492 6010
rect 4544 5958 4556 6010
rect 4608 5958 4620 6010
rect 4672 5958 4684 6010
rect 4736 5958 4748 6010
rect 4800 5958 11576 6010
rect 11628 5958 11640 6010
rect 11692 5958 11704 6010
rect 11756 5958 11768 6010
rect 11820 5958 11832 6010
rect 11884 5958 18660 6010
rect 18712 5958 18724 6010
rect 18776 5958 18788 6010
rect 18840 5958 18852 6010
rect 18904 5958 18916 6010
rect 18968 5958 25744 6010
rect 25796 5958 25808 6010
rect 25860 5958 25872 6010
rect 25924 5958 25936 6010
rect 25988 5958 26000 6010
rect 26052 5958 29440 6010
rect 1104 5936 29440 5958
rect 1394 5896 1400 5908
rect 1355 5868 1400 5896
rect 1394 5856 1400 5868
rect 1452 5856 1458 5908
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5721 5899 5779 5905
rect 5721 5896 5733 5899
rect 5224 5868 5733 5896
rect 5224 5856 5230 5868
rect 5721 5865 5733 5868
rect 5767 5865 5779 5899
rect 5721 5859 5779 5865
rect 6178 5856 6184 5908
rect 6236 5896 6242 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 6236 5868 7205 5896
rect 6236 5856 6242 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 9030 5856 9036 5908
rect 9088 5896 9094 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 9088 5868 9137 5896
rect 9088 5856 9094 5868
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 10594 5896 10600 5908
rect 10555 5868 10600 5896
rect 9125 5859 9183 5865
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 13081 5899 13139 5905
rect 13081 5865 13093 5899
rect 13127 5896 13139 5899
rect 14182 5896 14188 5908
rect 13127 5868 14188 5896
rect 13127 5865 13139 5868
rect 13081 5859 13139 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 14458 5856 14464 5908
rect 14516 5896 14522 5908
rect 15102 5896 15108 5908
rect 14516 5868 15108 5896
rect 14516 5856 14522 5868
rect 15102 5856 15108 5868
rect 15160 5896 15166 5908
rect 15197 5899 15255 5905
rect 15197 5896 15209 5899
rect 15160 5868 15209 5896
rect 15160 5856 15166 5868
rect 15197 5865 15209 5868
rect 15243 5865 15255 5899
rect 15197 5859 15255 5865
rect 15749 5899 15807 5905
rect 15749 5865 15761 5899
rect 15795 5896 15807 5899
rect 15838 5896 15844 5908
rect 15795 5868 15844 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 17126 5856 17132 5908
rect 17184 5896 17190 5908
rect 18325 5899 18383 5905
rect 18325 5896 18337 5899
rect 17184 5868 18337 5896
rect 17184 5856 17190 5868
rect 18325 5865 18337 5868
rect 18371 5896 18383 5899
rect 19518 5896 19524 5908
rect 18371 5868 19524 5896
rect 18371 5865 18383 5868
rect 18325 5859 18383 5865
rect 19518 5856 19524 5868
rect 19576 5896 19582 5908
rect 19889 5899 19947 5905
rect 19889 5896 19901 5899
rect 19576 5868 19901 5896
rect 19576 5856 19582 5868
rect 19889 5865 19901 5868
rect 19935 5865 19947 5899
rect 19889 5859 19947 5865
rect 21177 5899 21235 5905
rect 21177 5865 21189 5899
rect 21223 5896 21235 5899
rect 21266 5896 21272 5908
rect 21223 5868 21272 5896
rect 21223 5865 21235 5868
rect 21177 5859 21235 5865
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 22554 5896 22560 5908
rect 22515 5868 22560 5896
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 26786 5856 26792 5908
rect 26844 5896 26850 5908
rect 28537 5899 28595 5905
rect 28537 5896 28549 5899
rect 26844 5868 28549 5896
rect 26844 5856 26850 5868
rect 28537 5865 28549 5868
rect 28583 5865 28595 5899
rect 28537 5859 28595 5865
rect 4890 5788 4896 5840
rect 4948 5828 4954 5840
rect 6549 5831 6607 5837
rect 6549 5828 6561 5831
rect 4948 5800 6561 5828
rect 4948 5788 4954 5800
rect 6549 5797 6561 5800
rect 6595 5797 6607 5831
rect 13814 5828 13820 5840
rect 6549 5791 6607 5797
rect 12406 5800 13820 5828
rect 6012 5732 6684 5760
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5902 5692 5908 5704
rect 5863 5664 5908 5692
rect 5537 5655 5595 5661
rect 5552 5624 5580 5655
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6012 5701 6040 5732
rect 6656 5704 6684 5732
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 6454 5692 6460 5704
rect 6415 5664 6460 5692
rect 5997 5655 6055 5661
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6638 5692 6644 5704
rect 6599 5664 6644 5692
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 7926 5692 7932 5704
rect 7839 5664 7932 5692
rect 7926 5652 7932 5664
rect 7984 5692 7990 5704
rect 9030 5692 9036 5704
rect 7984 5664 9036 5692
rect 7984 5652 7990 5664
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 6472 5624 6500 5652
rect 5552 5596 6500 5624
rect 11149 5627 11207 5633
rect 11149 5593 11161 5627
rect 11195 5624 11207 5627
rect 12069 5627 12127 5633
rect 12069 5624 12081 5627
rect 11195 5596 12081 5624
rect 11195 5593 11207 5596
rect 11149 5587 11207 5593
rect 12069 5593 12081 5596
rect 12115 5624 12127 5627
rect 12406 5624 12434 5800
rect 13814 5788 13820 5800
rect 13872 5828 13878 5840
rect 17681 5831 17739 5837
rect 17681 5828 17693 5831
rect 13872 5800 17693 5828
rect 13872 5788 13878 5800
rect 17681 5797 17693 5800
rect 17727 5797 17739 5831
rect 17681 5791 17739 5797
rect 13280 5732 13768 5760
rect 13280 5704 13308 5732
rect 13262 5692 13268 5704
rect 13223 5664 13268 5692
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13449 5695 13507 5701
rect 13449 5661 13461 5695
rect 13495 5661 13507 5695
rect 13740 5692 13768 5732
rect 15102 5720 15108 5772
rect 15160 5760 15166 5772
rect 16117 5763 16175 5769
rect 16117 5760 16129 5763
rect 15160 5732 16129 5760
rect 15160 5720 15166 5732
rect 16117 5729 16129 5732
rect 16163 5760 16175 5763
rect 16577 5763 16635 5769
rect 16577 5760 16589 5763
rect 16163 5732 16589 5760
rect 16163 5729 16175 5732
rect 16117 5723 16175 5729
rect 16577 5729 16589 5732
rect 16623 5760 16635 5763
rect 16850 5760 16856 5772
rect 16623 5732 16856 5760
rect 16623 5729 16635 5732
rect 16577 5723 16635 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 17696 5760 17724 5791
rect 17954 5788 17960 5840
rect 18012 5828 18018 5840
rect 19245 5831 19303 5837
rect 19245 5828 19257 5831
rect 18012 5800 19257 5828
rect 18012 5788 18018 5800
rect 19245 5797 19257 5800
rect 19291 5797 19303 5831
rect 19245 5791 19303 5797
rect 21361 5831 21419 5837
rect 21361 5797 21373 5831
rect 21407 5828 21419 5831
rect 21910 5828 21916 5840
rect 21407 5800 21916 5828
rect 21407 5797 21419 5800
rect 21361 5791 21419 5797
rect 21910 5788 21916 5800
rect 21968 5788 21974 5840
rect 27985 5831 28043 5837
rect 27985 5797 27997 5831
rect 28031 5828 28043 5831
rect 28166 5828 28172 5840
rect 28031 5800 28172 5828
rect 28031 5797 28043 5800
rect 27985 5791 28043 5797
rect 28166 5788 28172 5800
rect 28224 5788 28230 5840
rect 18506 5760 18512 5772
rect 17696 5732 18512 5760
rect 18506 5720 18512 5732
rect 18564 5720 18570 5772
rect 19334 5760 19340 5772
rect 19260 5732 19340 5760
rect 13814 5692 13820 5704
rect 13740 5664 13820 5692
rect 13449 5655 13507 5661
rect 12115 5596 12434 5624
rect 12115 5593 12127 5596
rect 12069 5587 12127 5593
rect 13170 5584 13176 5636
rect 13228 5624 13234 5636
rect 13464 5624 13492 5655
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5692 15991 5695
rect 17034 5692 17040 5704
rect 15979 5664 17040 5692
rect 15979 5661 15991 5664
rect 15933 5655 15991 5661
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 19260 5701 19288 5732
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 19610 5720 19616 5772
rect 19668 5760 19674 5772
rect 20530 5760 20536 5772
rect 19668 5732 20536 5760
rect 19668 5720 19674 5732
rect 20530 5720 20536 5732
rect 20588 5760 20594 5772
rect 22830 5760 22836 5772
rect 20588 5732 22836 5760
rect 20588 5720 20594 5732
rect 22830 5720 22836 5732
rect 22888 5720 22894 5772
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5661 19303 5695
rect 19426 5692 19432 5704
rect 19387 5664 19432 5692
rect 19245 5655 19303 5661
rect 19426 5652 19432 5664
rect 19484 5652 19490 5704
rect 21821 5695 21879 5701
rect 21821 5692 21833 5695
rect 21008 5664 21833 5692
rect 14185 5627 14243 5633
rect 14185 5624 14197 5627
rect 13228 5596 14197 5624
rect 13228 5584 13234 5596
rect 14185 5593 14197 5596
rect 14231 5624 14243 5627
rect 14737 5627 14795 5633
rect 14737 5624 14749 5627
rect 14231 5596 14749 5624
rect 14231 5593 14243 5596
rect 14185 5587 14243 5593
rect 14737 5593 14749 5596
rect 14783 5624 14795 5627
rect 15470 5624 15476 5636
rect 14783 5596 15476 5624
rect 14783 5593 14795 5596
rect 14737 5587 14795 5593
rect 15470 5584 15476 5596
rect 15528 5584 15534 5636
rect 17494 5584 17500 5636
rect 17552 5624 17558 5636
rect 21008 5633 21036 5664
rect 21821 5661 21833 5664
rect 21867 5661 21879 5695
rect 28718 5692 28724 5704
rect 28679 5664 28724 5692
rect 21821 5655 21879 5661
rect 28718 5652 28724 5664
rect 28776 5652 28782 5704
rect 20993 5627 21051 5633
rect 20993 5624 21005 5627
rect 17552 5596 21005 5624
rect 17552 5584 17558 5596
rect 20993 5593 21005 5596
rect 21039 5593 21051 5627
rect 20993 5587 21051 5593
rect 21174 5584 21180 5636
rect 21232 5633 21238 5636
rect 21232 5627 21251 5633
rect 21239 5593 21251 5627
rect 21232 5587 21251 5593
rect 21232 5584 21238 5587
rect 7834 5556 7840 5568
rect 7795 5528 7840 5556
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 17034 5516 17040 5568
rect 17092 5556 17098 5568
rect 17221 5559 17279 5565
rect 17221 5556 17233 5559
rect 17092 5528 17233 5556
rect 17092 5516 17098 5528
rect 17221 5525 17233 5528
rect 17267 5556 17279 5559
rect 17770 5556 17776 5568
rect 17267 5528 17776 5556
rect 17267 5525 17279 5528
rect 17221 5519 17279 5525
rect 17770 5516 17776 5528
rect 17828 5556 17834 5568
rect 22462 5556 22468 5568
rect 17828 5528 22468 5556
rect 17828 5516 17834 5528
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 1104 5466 29600 5488
rect 1104 5414 8034 5466
rect 8086 5414 8098 5466
rect 8150 5414 8162 5466
rect 8214 5414 8226 5466
rect 8278 5414 8290 5466
rect 8342 5414 15118 5466
rect 15170 5414 15182 5466
rect 15234 5414 15246 5466
rect 15298 5414 15310 5466
rect 15362 5414 15374 5466
rect 15426 5414 22202 5466
rect 22254 5414 22266 5466
rect 22318 5414 22330 5466
rect 22382 5414 22394 5466
rect 22446 5414 22458 5466
rect 22510 5414 29286 5466
rect 29338 5414 29350 5466
rect 29402 5414 29414 5466
rect 29466 5414 29478 5466
rect 29530 5414 29542 5466
rect 29594 5414 29600 5466
rect 1104 5392 29600 5414
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 6696 5324 6837 5352
rect 6696 5312 6702 5324
rect 6825 5321 6837 5324
rect 6871 5321 6883 5355
rect 6825 5315 6883 5321
rect 7926 5312 7932 5364
rect 7984 5352 7990 5364
rect 8021 5355 8079 5361
rect 8021 5352 8033 5355
rect 7984 5324 8033 5352
rect 7984 5312 7990 5324
rect 8021 5321 8033 5324
rect 8067 5321 8079 5355
rect 10042 5352 10048 5364
rect 10003 5324 10048 5352
rect 8021 5315 8079 5321
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 10870 5352 10876 5364
rect 10831 5324 10876 5352
rect 10870 5312 10876 5324
rect 10928 5312 10934 5364
rect 13814 5352 13820 5364
rect 13775 5324 13820 5352
rect 13814 5312 13820 5324
rect 13872 5352 13878 5364
rect 14366 5352 14372 5364
rect 13872 5324 14372 5352
rect 13872 5312 13878 5324
rect 14366 5312 14372 5324
rect 14424 5352 14430 5364
rect 14645 5355 14703 5361
rect 14645 5352 14657 5355
rect 14424 5324 14657 5352
rect 14424 5312 14430 5324
rect 14645 5321 14657 5324
rect 14691 5321 14703 5355
rect 14645 5315 14703 5321
rect 15473 5355 15531 5361
rect 15473 5321 15485 5355
rect 15519 5352 15531 5355
rect 17034 5352 17040 5364
rect 15519 5324 17040 5352
rect 15519 5321 15531 5324
rect 15473 5315 15531 5321
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 17865 5355 17923 5361
rect 17865 5321 17877 5355
rect 17911 5352 17923 5355
rect 18046 5352 18052 5364
rect 17911 5324 18052 5352
rect 17911 5321 17923 5324
rect 17865 5315 17923 5321
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 18322 5312 18328 5364
rect 18380 5352 18386 5364
rect 18601 5355 18659 5361
rect 18601 5352 18613 5355
rect 18380 5324 18613 5352
rect 18380 5312 18386 5324
rect 18601 5321 18613 5324
rect 18647 5321 18659 5355
rect 22554 5352 22560 5364
rect 18601 5315 18659 5321
rect 22112 5324 22560 5352
rect 22112 5293 22140 5324
rect 22554 5312 22560 5324
rect 22612 5352 22618 5364
rect 23014 5352 23020 5364
rect 22612 5324 23020 5352
rect 22612 5312 22618 5324
rect 23014 5312 23020 5324
rect 23072 5312 23078 5364
rect 28718 5352 28724 5364
rect 28679 5324 28724 5352
rect 28718 5312 28724 5324
rect 28776 5312 28782 5364
rect 22097 5287 22155 5293
rect 22097 5253 22109 5287
rect 22143 5253 22155 5287
rect 22097 5247 22155 5253
rect 7190 5216 7196 5228
rect 7151 5188 7196 5216
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 21818 5216 21824 5228
rect 21779 5188 21824 5216
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 21910 5176 21916 5228
rect 21968 5216 21974 5228
rect 21968 5188 22013 5216
rect 21968 5176 21974 5188
rect 7098 5148 7104 5160
rect 7011 5120 7104 5148
rect 7098 5108 7104 5120
rect 7156 5148 7162 5160
rect 7834 5148 7840 5160
rect 7156 5120 7840 5148
rect 7156 5108 7162 5120
rect 7834 5108 7840 5120
rect 7892 5108 7898 5160
rect 15930 5108 15936 5160
rect 15988 5148 15994 5160
rect 22112 5148 22140 5247
rect 22186 5244 22192 5296
rect 22244 5284 22250 5296
rect 22244 5256 22289 5284
rect 22244 5244 22250 5256
rect 22281 5219 22339 5225
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 22554 5216 22560 5228
rect 22327 5188 22560 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 22554 5176 22560 5188
rect 22612 5176 22618 5228
rect 23382 5176 23388 5228
rect 23440 5216 23446 5228
rect 23661 5219 23719 5225
rect 23661 5216 23673 5219
rect 23440 5188 23673 5216
rect 23440 5176 23446 5188
rect 23661 5185 23673 5188
rect 23707 5185 23719 5219
rect 23661 5179 23719 5185
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 24121 5219 24179 5225
rect 24121 5216 24133 5219
rect 23808 5188 24133 5216
rect 23808 5176 23814 5188
rect 24121 5185 24133 5188
rect 24167 5216 24179 5219
rect 24673 5219 24731 5225
rect 24673 5216 24685 5219
rect 24167 5188 24685 5216
rect 24167 5185 24179 5188
rect 24121 5179 24179 5185
rect 24673 5185 24685 5188
rect 24719 5185 24731 5219
rect 24673 5179 24731 5185
rect 22925 5151 22983 5157
rect 22925 5148 22937 5151
rect 15988 5120 22140 5148
rect 22480 5120 22937 5148
rect 15988 5108 15994 5120
rect 22480 5092 22508 5120
rect 22925 5117 22937 5120
rect 22971 5117 22983 5151
rect 22925 5111 22983 5117
rect 22462 5080 22468 5092
rect 22375 5052 22468 5080
rect 22462 5040 22468 5052
rect 22520 5040 22526 5092
rect 23385 5083 23443 5089
rect 23385 5049 23397 5083
rect 23431 5080 23443 5083
rect 23474 5080 23480 5092
rect 23431 5052 23480 5080
rect 23431 5049 23443 5052
rect 23385 5043 23443 5049
rect 23474 5040 23480 5052
rect 23532 5040 23538 5092
rect 5813 5015 5871 5021
rect 5813 4981 5825 5015
rect 5859 5012 5871 5015
rect 6730 5012 6736 5024
rect 5859 4984 6736 5012
rect 5859 4981 5871 4984
rect 5813 4975 5871 4981
rect 6730 4972 6736 4984
rect 6788 5012 6794 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 6788 4984 7205 5012
rect 6788 4972 6794 4984
rect 7193 4981 7205 4984
rect 7239 5012 7251 5015
rect 8478 5012 8484 5024
rect 7239 4984 8484 5012
rect 7239 4981 7251 4984
rect 7193 4975 7251 4981
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 19150 5012 19156 5024
rect 19111 4984 19156 5012
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 19242 4972 19248 5024
rect 19300 5012 19306 5024
rect 19797 5015 19855 5021
rect 19797 5012 19809 5015
rect 19300 4984 19809 5012
rect 19300 4972 19306 4984
rect 19797 4981 19809 4984
rect 19843 5012 19855 5015
rect 23106 5012 23112 5024
rect 19843 4984 23112 5012
rect 19843 4981 19855 4984
rect 19797 4975 19855 4981
rect 23106 4972 23112 4984
rect 23164 4972 23170 5024
rect 1104 4922 29440 4944
rect 1104 4870 4492 4922
rect 4544 4870 4556 4922
rect 4608 4870 4620 4922
rect 4672 4870 4684 4922
rect 4736 4870 4748 4922
rect 4800 4870 11576 4922
rect 11628 4870 11640 4922
rect 11692 4870 11704 4922
rect 11756 4870 11768 4922
rect 11820 4870 11832 4922
rect 11884 4870 18660 4922
rect 18712 4870 18724 4922
rect 18776 4870 18788 4922
rect 18840 4870 18852 4922
rect 18904 4870 18916 4922
rect 18968 4870 25744 4922
rect 25796 4870 25808 4922
rect 25860 4870 25872 4922
rect 25924 4870 25936 4922
rect 25988 4870 26000 4922
rect 26052 4870 29440 4922
rect 1104 4848 29440 4870
rect 2133 4811 2191 4817
rect 2133 4777 2145 4811
rect 2179 4808 2191 4811
rect 4338 4808 4344 4820
rect 2179 4780 4344 4808
rect 2179 4777 2191 4780
rect 2133 4771 2191 4777
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 6641 4811 6699 4817
rect 6641 4808 6653 4811
rect 6512 4780 6653 4808
rect 6512 4768 6518 4780
rect 6641 4777 6653 4780
rect 6687 4777 6699 4811
rect 6641 4771 6699 4777
rect 6730 4768 6736 4820
rect 6788 4808 6794 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 6788 4780 7297 4808
rect 6788 4768 6794 4780
rect 7285 4777 7297 4780
rect 7331 4777 7343 4811
rect 10502 4808 10508 4820
rect 10463 4780 10508 4808
rect 7285 4771 7343 4777
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 14366 4808 14372 4820
rect 14327 4780 14372 4808
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15470 4808 15476 4820
rect 15252 4780 15476 4808
rect 15252 4768 15258 4780
rect 15470 4768 15476 4780
rect 15528 4808 15534 4820
rect 15749 4811 15807 4817
rect 15749 4808 15761 4811
rect 15528 4780 15761 4808
rect 15528 4768 15534 4780
rect 15749 4777 15761 4780
rect 15795 4808 15807 4811
rect 19242 4808 19248 4820
rect 15795 4780 19248 4808
rect 15795 4777 15807 4780
rect 15749 4771 15807 4777
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 19889 4811 19947 4817
rect 19889 4777 19901 4811
rect 19935 4808 19947 4811
rect 20254 4808 20260 4820
rect 19935 4780 20260 4808
rect 19935 4777 19947 4780
rect 19889 4771 19947 4777
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 23382 4808 23388 4820
rect 21100 4780 23388 4808
rect 14384 4740 14412 4768
rect 14458 4740 14464 4752
rect 14371 4712 14464 4740
rect 14458 4700 14464 4712
rect 14516 4740 14522 4752
rect 16209 4743 16267 4749
rect 16209 4740 16221 4743
rect 14516 4712 16221 4740
rect 14516 4700 14522 4712
rect 16209 4709 16221 4712
rect 16255 4709 16267 4743
rect 17770 4740 17776 4752
rect 17731 4712 17776 4740
rect 16209 4703 16267 4709
rect 17770 4700 17776 4712
rect 17828 4700 17834 4752
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4672 6607 4675
rect 7190 4672 7196 4684
rect 6595 4644 7196 4672
rect 6595 4641 6607 4644
rect 6549 4635 6607 4641
rect 7190 4632 7196 4644
rect 7248 4672 7254 4684
rect 9306 4672 9312 4684
rect 7248 4644 9312 4672
rect 7248 4632 7254 4644
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 9766 4672 9772 4684
rect 9508 4644 9772 4672
rect 6825 4607 6883 4613
rect 6825 4573 6837 4607
rect 6871 4604 6883 4607
rect 7098 4604 7104 4616
rect 6871 4576 7104 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 7098 4564 7104 4576
rect 7156 4564 7162 4616
rect 9508 4613 9536 4644
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 12618 4672 12624 4684
rect 12406 4644 12624 4672
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4604 9735 4607
rect 10502 4604 10508 4616
rect 9723 4576 10508 4604
rect 9723 4573 9735 4576
rect 9677 4567 9735 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 1578 4496 1584 4548
rect 1636 4536 1642 4548
rect 1857 4539 1915 4545
rect 1857 4536 1869 4539
rect 1636 4508 1869 4536
rect 1636 4496 1642 4508
rect 1857 4505 1869 4508
rect 1903 4505 1915 4539
rect 1857 4499 1915 4505
rect 10042 4496 10048 4548
rect 10100 4536 10106 4548
rect 10137 4539 10195 4545
rect 10137 4536 10149 4539
rect 10100 4508 10149 4536
rect 10100 4496 10106 4508
rect 10137 4505 10149 4508
rect 10183 4505 10195 4539
rect 10137 4499 10195 4505
rect 10321 4539 10379 4545
rect 10321 4505 10333 4539
rect 10367 4536 10379 4539
rect 10594 4536 10600 4548
rect 10367 4508 10600 4536
rect 10367 4505 10379 4508
rect 10321 4499 10379 4505
rect 10594 4496 10600 4508
rect 10652 4536 10658 4548
rect 10965 4539 11023 4545
rect 10965 4536 10977 4539
rect 10652 4508 10977 4536
rect 10652 4496 10658 4508
rect 10965 4505 10977 4508
rect 11011 4536 11023 4539
rect 12406 4536 12434 4644
rect 12618 4632 12624 4644
rect 12676 4672 12682 4684
rect 19150 4672 19156 4684
rect 12676 4644 19156 4672
rect 12676 4632 12682 4644
rect 19150 4632 19156 4644
rect 19208 4632 19214 4684
rect 20530 4672 20536 4684
rect 20491 4644 20536 4672
rect 20530 4632 20536 4644
rect 20588 4672 20594 4684
rect 20993 4675 21051 4681
rect 20993 4672 21005 4675
rect 20588 4644 21005 4672
rect 20588 4632 20594 4644
rect 20993 4641 21005 4644
rect 21039 4641 21051 4675
rect 20993 4635 21051 4641
rect 14185 4607 14243 4613
rect 14185 4573 14197 4607
rect 14231 4604 14243 4607
rect 14274 4604 14280 4616
rect 14231 4576 14280 4604
rect 14231 4573 14243 4576
rect 14185 4567 14243 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4604 14427 4607
rect 14550 4604 14556 4616
rect 14415 4576 14556 4604
rect 14415 4573 14427 4576
rect 14369 4567 14427 4573
rect 14550 4564 14556 4576
rect 14608 4604 14614 4616
rect 15105 4607 15163 4613
rect 15105 4604 15117 4607
rect 14608 4576 15117 4604
rect 14608 4564 14614 4576
rect 15105 4573 15117 4576
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 15194 4564 15200 4616
rect 15252 4604 15258 4616
rect 20070 4604 20076 4616
rect 15252 4576 15297 4604
rect 20031 4576 20076 4604
rect 15252 4564 15258 4576
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20395 4607 20453 4613
rect 20395 4573 20407 4607
rect 20441 4604 20453 4607
rect 20622 4604 20628 4616
rect 20441 4576 20628 4604
rect 20441 4573 20453 4576
rect 20395 4567 20453 4573
rect 20622 4564 20628 4576
rect 20680 4604 20686 4616
rect 21100 4604 21128 4780
rect 23382 4768 23388 4780
rect 23440 4768 23446 4820
rect 22002 4740 22008 4752
rect 21963 4712 22008 4740
rect 22002 4700 22008 4712
rect 22060 4740 22066 4752
rect 23658 4740 23664 4752
rect 22060 4712 23664 4740
rect 22060 4700 22066 4712
rect 20680 4576 21128 4604
rect 20680 4564 20686 4576
rect 22462 4564 22468 4616
rect 22520 4604 22526 4616
rect 22756 4613 22784 4712
rect 23216 4613 23244 4712
rect 23658 4700 23664 4712
rect 23716 4740 23722 4752
rect 24397 4743 24455 4749
rect 24397 4740 24409 4743
rect 23716 4712 24409 4740
rect 23716 4700 23722 4712
rect 24397 4709 24409 4712
rect 24443 4709 24455 4743
rect 24397 4703 24455 4709
rect 22557 4607 22615 4613
rect 22557 4604 22569 4607
rect 22520 4576 22569 4604
rect 22520 4564 22526 4576
rect 22557 4573 22569 4576
rect 22603 4573 22615 4607
rect 22557 4567 22615 4573
rect 22741 4607 22799 4613
rect 22741 4573 22753 4607
rect 22787 4573 22799 4607
rect 22741 4567 22799 4573
rect 23201 4607 23259 4613
rect 23201 4573 23213 4607
rect 23247 4573 23259 4607
rect 23201 4567 23259 4573
rect 11011 4508 12434 4536
rect 11011 4505 11023 4508
rect 10965 4499 11023 4505
rect 19334 4496 19340 4548
rect 19392 4536 19398 4548
rect 20165 4539 20223 4545
rect 20165 4536 20177 4539
rect 19392 4508 20177 4536
rect 19392 4496 19398 4508
rect 20165 4505 20177 4508
rect 20211 4505 20223 4539
rect 20165 4499 20223 4505
rect 20257 4539 20315 4545
rect 20257 4505 20269 4539
rect 20303 4505 20315 4539
rect 20257 4499 20315 4505
rect 14366 4428 14372 4480
rect 14424 4468 14430 4480
rect 14553 4471 14611 4477
rect 14553 4468 14565 4471
rect 14424 4440 14565 4468
rect 14424 4428 14430 4440
rect 14553 4437 14565 4440
rect 14599 4437 14611 4471
rect 20272 4468 20300 4499
rect 20714 4468 20720 4480
rect 20272 4440 20720 4468
rect 14553 4431 14611 4437
rect 20714 4428 20720 4440
rect 20772 4428 20778 4480
rect 22741 4471 22799 4477
rect 22741 4437 22753 4471
rect 22787 4468 22799 4471
rect 23198 4468 23204 4480
rect 22787 4440 23204 4468
rect 22787 4437 22799 4440
rect 22741 4431 22799 4437
rect 23198 4428 23204 4440
rect 23256 4428 23262 4480
rect 1104 4378 29600 4400
rect 1104 4326 8034 4378
rect 8086 4326 8098 4378
rect 8150 4326 8162 4378
rect 8214 4326 8226 4378
rect 8278 4326 8290 4378
rect 8342 4326 15118 4378
rect 15170 4326 15182 4378
rect 15234 4326 15246 4378
rect 15298 4326 15310 4378
rect 15362 4326 15374 4378
rect 15426 4326 22202 4378
rect 22254 4326 22266 4378
rect 22318 4326 22330 4378
rect 22382 4326 22394 4378
rect 22446 4326 22458 4378
rect 22510 4326 29286 4378
rect 29338 4326 29350 4378
rect 29402 4326 29414 4378
rect 29466 4326 29478 4378
rect 29530 4326 29542 4378
rect 29594 4326 29600 4378
rect 1104 4304 29600 4326
rect 10594 4224 10600 4276
rect 10652 4264 10658 4276
rect 10873 4267 10931 4273
rect 10873 4264 10885 4267
rect 10652 4236 10885 4264
rect 10652 4224 10658 4236
rect 10873 4233 10885 4236
rect 10919 4233 10931 4267
rect 10873 4227 10931 4233
rect 12713 4267 12771 4273
rect 12713 4233 12725 4267
rect 12759 4264 12771 4267
rect 15930 4264 15936 4276
rect 12759 4236 13032 4264
rect 12759 4233 12771 4236
rect 12713 4227 12771 4233
rect 1578 4196 1584 4208
rect 1539 4168 1584 4196
rect 1578 4156 1584 4168
rect 1636 4156 1642 4208
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2455 4100 2774 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2746 4060 2774 4100
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9824 4100 10057 4128
rect 9824 4088 9830 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 10612 4128 10640 4224
rect 10459 4100 10640 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 2958 4060 2964 4072
rect 2746 4032 2964 4060
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 10244 4060 10272 4091
rect 10962 4088 10968 4140
rect 11020 4128 11026 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11020 4100 11529 4128
rect 11020 4088 11026 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 11716 4060 11744 4091
rect 11974 4088 11980 4140
rect 12032 4128 12038 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12032 4100 12909 4128
rect 12032 4088 12038 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 13004 4128 13032 4236
rect 15396 4236 15936 4264
rect 13173 4199 13231 4205
rect 13173 4165 13185 4199
rect 13219 4196 13231 4199
rect 14918 4196 14924 4208
rect 13219 4168 14924 4196
rect 13219 4165 13231 4168
rect 13173 4159 13231 4165
rect 14918 4156 14924 4168
rect 14976 4156 14982 4208
rect 15194 4205 15200 4208
rect 15181 4199 15200 4205
rect 15181 4165 15193 4199
rect 15181 4159 15200 4165
rect 15194 4156 15200 4159
rect 15252 4156 15258 4208
rect 15396 4205 15424 4236
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 20625 4267 20683 4273
rect 20625 4233 20637 4267
rect 20671 4264 20683 4267
rect 20714 4264 20720 4276
rect 20671 4236 20720 4264
rect 20671 4233 20683 4236
rect 20625 4227 20683 4233
rect 20714 4224 20720 4236
rect 20772 4224 20778 4276
rect 22281 4267 22339 4273
rect 22281 4233 22293 4267
rect 22327 4264 22339 4267
rect 22554 4264 22560 4276
rect 22327 4236 22560 4264
rect 22327 4233 22339 4236
rect 22281 4227 22339 4233
rect 22554 4224 22560 4236
rect 22612 4224 22618 4276
rect 15381 4199 15439 4205
rect 15381 4165 15393 4199
rect 15427 4165 15439 4199
rect 15381 4159 15439 4165
rect 16758 4156 16764 4208
rect 16816 4196 16822 4208
rect 16853 4199 16911 4205
rect 16853 4196 16865 4199
rect 16816 4168 16865 4196
rect 16816 4156 16822 4168
rect 16853 4165 16865 4168
rect 16899 4196 16911 4199
rect 17770 4196 17776 4208
rect 16899 4168 17776 4196
rect 16899 4165 16911 4168
rect 16853 4159 16911 4165
rect 14274 4128 14280 4140
rect 13004 4100 13676 4128
rect 14235 4100 14280 4128
rect 12897 4091 12955 4097
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 10060 4032 12173 4060
rect 10060 4004 10088 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4060 13139 4063
rect 13538 4060 13544 4072
rect 13127 4032 13544 4060
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 9585 3995 9643 4001
rect 9585 3961 9597 3995
rect 9631 3992 9643 3995
rect 10042 3992 10048 4004
rect 9631 3964 10048 3992
rect 9631 3961 9643 3964
rect 9585 3955 9643 3961
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 11422 3952 11428 4004
rect 11480 3992 11486 4004
rect 13648 3992 13676 4100
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 14550 4128 14556 4140
rect 14511 4100 14556 4128
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 17328 4137 17356 4168
rect 17770 4156 17776 4168
rect 17828 4156 17834 4208
rect 18046 4156 18052 4208
rect 18104 4196 18110 4208
rect 23385 4199 23443 4205
rect 18104 4168 19104 4196
rect 18104 4156 18110 4168
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 17954 4128 17960 4140
rect 17543 4100 17960 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17954 4088 17960 4100
rect 18012 4128 18018 4140
rect 19076 4137 19104 4168
rect 23385 4165 23397 4199
rect 23431 4196 23443 4199
rect 23431 4168 23520 4196
rect 23431 4165 23443 4168
rect 23385 4159 23443 4165
rect 18141 4131 18199 4137
rect 18141 4128 18153 4131
rect 18012 4100 18153 4128
rect 18012 4088 18018 4100
rect 18141 4097 18153 4100
rect 18187 4097 18199 4131
rect 18141 4091 18199 4097
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4128 19119 4131
rect 19521 4131 19579 4137
rect 19521 4128 19533 4131
rect 19107 4100 19533 4128
rect 19107 4097 19119 4100
rect 19061 4091 19119 4097
rect 19521 4097 19533 4100
rect 19567 4097 19579 4131
rect 20898 4128 20904 4140
rect 20859 4100 20904 4128
rect 19521 4091 19579 4097
rect 20898 4088 20904 4100
rect 20956 4088 20962 4140
rect 21818 4128 21824 4140
rect 21779 4100 21824 4128
rect 21818 4088 21824 4100
rect 21876 4088 21882 4140
rect 21910 4088 21916 4140
rect 21968 4128 21974 4140
rect 22097 4131 22155 4137
rect 21968 4100 22013 4128
rect 21968 4088 21974 4100
rect 22097 4097 22109 4131
rect 22143 4097 22155 4131
rect 23198 4128 23204 4140
rect 23159 4100 23204 4128
rect 22097 4091 22155 4097
rect 14458 4060 14464 4072
rect 14419 4032 14464 4060
rect 14458 4020 14464 4032
rect 14516 4020 14522 4072
rect 14844 4032 16436 4060
rect 14844 3992 14872 4032
rect 15010 3992 15016 4004
rect 11480 3964 12434 3992
rect 13648 3964 14872 3992
rect 14971 3964 15016 3992
rect 11480 3952 11486 3964
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 2225 3927 2283 3933
rect 2225 3924 2237 3927
rect 1728 3896 2237 3924
rect 1728 3884 1734 3896
rect 2225 3893 2237 3896
rect 2271 3893 2283 3927
rect 2225 3887 2283 3893
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11020 3896 11529 3924
rect 11020 3884 11026 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 12406 3924 12434 3964
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 16408 3992 16436 4032
rect 17770 4020 17776 4072
rect 17828 4060 17834 4072
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 17828 4032 18337 4060
rect 17828 4020 17834 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 18325 4023 18383 4029
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4060 18475 4063
rect 18969 4063 19027 4069
rect 18969 4060 18981 4063
rect 18463 4032 18981 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 18969 4029 18981 4032
rect 19015 4029 19027 4063
rect 18969 4023 19027 4029
rect 20625 4063 20683 4069
rect 20625 4029 20637 4063
rect 20671 4029 20683 4063
rect 20806 4060 20812 4072
rect 20767 4032 20812 4060
rect 20625 4023 20683 4029
rect 19334 3992 19340 4004
rect 16408 3964 19340 3992
rect 19334 3952 19340 3964
rect 19392 3952 19398 4004
rect 20640 3992 20668 4023
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 21450 4020 21456 4072
rect 21508 4060 21514 4072
rect 22112 4060 22140 4091
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 23290 4088 23296 4140
rect 23348 4128 23354 4140
rect 23492 4128 23520 4168
rect 23348 4100 23393 4128
rect 23492 4100 23796 4128
rect 23348 4088 23354 4100
rect 23658 4060 23664 4072
rect 21508 4032 22140 4060
rect 23619 4032 23664 4060
rect 21508 4020 21514 4032
rect 23658 4020 23664 4032
rect 23716 4020 23722 4072
rect 23768 4060 23796 4100
rect 23842 4088 23848 4140
rect 23900 4128 23906 4140
rect 24121 4131 24179 4137
rect 24121 4128 24133 4131
rect 23900 4100 24133 4128
rect 23900 4088 23906 4100
rect 24121 4097 24133 4100
rect 24167 4097 24179 4131
rect 24121 4091 24179 4097
rect 24305 4131 24363 4137
rect 24305 4097 24317 4131
rect 24351 4128 24363 4131
rect 24765 4131 24823 4137
rect 24765 4128 24777 4131
rect 24351 4100 24777 4128
rect 24351 4097 24363 4100
rect 24305 4091 24363 4097
rect 24765 4097 24777 4100
rect 24811 4097 24823 4131
rect 24765 4091 24823 4097
rect 24213 4063 24271 4069
rect 24213 4060 24225 4063
rect 23768 4032 24225 4060
rect 24213 4029 24225 4032
rect 24259 4029 24271 4063
rect 24213 4023 24271 4029
rect 20990 3992 20996 4004
rect 20640 3964 20996 3992
rect 20990 3952 20996 3964
rect 21048 3992 21054 4004
rect 22738 3992 22744 4004
rect 21048 3964 22744 3992
rect 21048 3952 21054 3964
rect 22738 3952 22744 3964
rect 22796 3952 22802 4004
rect 23014 3952 23020 4004
rect 23072 3992 23078 4004
rect 24320 3992 24348 4091
rect 23072 3964 24348 3992
rect 23072 3952 23078 3964
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 12406 3896 12909 3924
rect 11517 3887 11575 3893
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 14090 3924 14096 3936
rect 14051 3896 14096 3924
rect 12897 3887 12955 3893
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 15197 3927 15255 3933
rect 15197 3893 15209 3927
rect 15243 3924 15255 3927
rect 15286 3924 15292 3936
rect 15243 3896 15292 3924
rect 15243 3893 15255 3896
rect 15197 3887 15255 3893
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 15838 3884 15844 3936
rect 15896 3924 15902 3936
rect 17218 3924 17224 3936
rect 15896 3896 17224 3924
rect 15896 3884 15902 3896
rect 17218 3884 17224 3896
rect 17276 3884 17282 3936
rect 17497 3927 17555 3933
rect 17497 3893 17509 3927
rect 17543 3924 17555 3927
rect 17862 3924 17868 3936
rect 17543 3896 17868 3924
rect 17543 3893 17555 3896
rect 17497 3887 17555 3893
rect 17862 3884 17868 3896
rect 17920 3884 17926 3936
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 22922 3924 22928 3936
rect 18012 3896 18057 3924
rect 22883 3896 22928 3924
rect 18012 3884 18018 3896
rect 22922 3884 22928 3896
rect 22980 3884 22986 3936
rect 23474 3884 23480 3936
rect 23532 3924 23538 3936
rect 23569 3927 23627 3933
rect 23569 3924 23581 3927
rect 23532 3896 23581 3924
rect 23532 3884 23538 3896
rect 23569 3893 23581 3896
rect 23615 3893 23627 3927
rect 28626 3924 28632 3936
rect 28587 3896 28632 3924
rect 23569 3887 23627 3893
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 1104 3834 29440 3856
rect 1104 3782 4492 3834
rect 4544 3782 4556 3834
rect 4608 3782 4620 3834
rect 4672 3782 4684 3834
rect 4736 3782 4748 3834
rect 4800 3782 11576 3834
rect 11628 3782 11640 3834
rect 11692 3782 11704 3834
rect 11756 3782 11768 3834
rect 11820 3782 11832 3834
rect 11884 3782 18660 3834
rect 18712 3782 18724 3834
rect 18776 3782 18788 3834
rect 18840 3782 18852 3834
rect 18904 3782 18916 3834
rect 18968 3782 25744 3834
rect 25796 3782 25808 3834
rect 25860 3782 25872 3834
rect 25924 3782 25936 3834
rect 25988 3782 26000 3834
rect 26052 3782 29440 3834
rect 1104 3760 29440 3782
rect 10965 3723 11023 3729
rect 10965 3689 10977 3723
rect 11011 3720 11023 3723
rect 13538 3720 13544 3732
rect 11011 3692 11652 3720
rect 13499 3692 13544 3720
rect 11011 3689 11023 3692
rect 10965 3683 11023 3689
rect 10962 3584 10968 3596
rect 10520 3556 10968 3584
rect 1670 3516 1676 3528
rect 1631 3488 1676 3516
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 10520 3525 10548 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11422 3544 11428 3596
rect 11480 3584 11486 3596
rect 11517 3587 11575 3593
rect 11517 3584 11529 3587
rect 11480 3556 11529 3584
rect 11480 3544 11486 3556
rect 11517 3553 11529 3556
rect 11563 3553 11575 3587
rect 11517 3547 11575 3553
rect 11624 3525 11652 3692
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 13630 3680 13636 3732
rect 13688 3720 13694 3732
rect 14185 3723 14243 3729
rect 14185 3720 14197 3723
rect 13688 3692 14197 3720
rect 13688 3680 13694 3692
rect 14185 3689 14197 3692
rect 14231 3689 14243 3723
rect 14185 3683 14243 3689
rect 14645 3723 14703 3729
rect 14645 3689 14657 3723
rect 14691 3720 14703 3723
rect 15194 3720 15200 3732
rect 14691 3692 15200 3720
rect 14691 3689 14703 3692
rect 14645 3683 14703 3689
rect 15194 3680 15200 3692
rect 15252 3720 15258 3732
rect 15657 3723 15715 3729
rect 15657 3720 15669 3723
rect 15252 3692 15669 3720
rect 15252 3680 15258 3692
rect 15657 3689 15669 3692
rect 15703 3720 15715 3723
rect 16574 3720 16580 3732
rect 15703 3692 16580 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 16853 3723 16911 3729
rect 16853 3689 16865 3723
rect 16899 3720 16911 3723
rect 20070 3720 20076 3732
rect 16899 3692 19932 3720
rect 20031 3692 20076 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 11977 3655 12035 3661
rect 11977 3621 11989 3655
rect 12023 3652 12035 3655
rect 12023 3624 13308 3652
rect 12023 3621 12035 3624
rect 11977 3615 12035 3621
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3485 10563 3519
rect 10505 3479 10563 3485
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3485 10839 3519
rect 10781 3479 10839 3485
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3516 11667 3519
rect 11974 3516 11980 3528
rect 11655 3488 11980 3516
rect 11655 3485 11667 3488
rect 11609 3479 11667 3485
rect 10594 3448 10600 3460
rect 10555 3420 10600 3448
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 10796 3448 10824 3479
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12618 3516 12624 3528
rect 12579 3488 12624 3516
rect 12618 3476 12624 3488
rect 12676 3476 12682 3528
rect 13280 3525 13308 3624
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13265 3519 13323 3525
rect 13265 3485 13277 3519
rect 13311 3516 13323 3519
rect 13354 3516 13360 3528
rect 13311 3488 13360 3516
rect 13311 3485 13323 3488
rect 13265 3479 13323 3485
rect 11514 3448 11520 3460
rect 10796 3420 11520 3448
rect 11514 3408 11520 3420
rect 11572 3448 11578 3460
rect 13096 3448 13124 3479
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 13556 3516 13584 3680
rect 15838 3652 15844 3664
rect 15799 3624 15844 3652
rect 15838 3612 15844 3624
rect 15896 3612 15902 3664
rect 17310 3652 17316 3664
rect 17271 3624 17316 3652
rect 17310 3612 17316 3624
rect 17368 3612 17374 3664
rect 18138 3612 18144 3664
rect 18196 3652 18202 3664
rect 18601 3655 18659 3661
rect 18601 3652 18613 3655
rect 18196 3624 18613 3652
rect 18196 3612 18202 3624
rect 18601 3621 18613 3624
rect 18647 3621 18659 3655
rect 18601 3615 18659 3621
rect 16574 3544 16580 3596
rect 16632 3584 16638 3596
rect 16632 3556 16677 3584
rect 16632 3544 16638 3556
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 17589 3587 17647 3593
rect 17589 3584 17601 3587
rect 17276 3556 17601 3584
rect 17276 3544 17282 3556
rect 17589 3553 17601 3556
rect 17635 3553 17647 3587
rect 19521 3587 19579 3593
rect 19521 3584 19533 3587
rect 17589 3547 17647 3553
rect 17788 3556 19533 3584
rect 13906 3516 13912 3528
rect 13556 3488 13912 3516
rect 13906 3476 13912 3488
rect 13964 3516 13970 3528
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13964 3488 14105 3516
rect 13964 3476 13970 3488
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 14458 3516 14464 3528
rect 14419 3488 14464 3516
rect 14093 3479 14151 3485
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 16390 3516 16396 3528
rect 16351 3488 16396 3516
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3485 16543 3519
rect 16485 3479 16543 3485
rect 16672 3519 16730 3525
rect 16672 3485 16684 3519
rect 16718 3518 16730 3519
rect 16718 3516 16804 3518
rect 17678 3516 17684 3528
rect 16718 3490 16896 3516
rect 16718 3485 16730 3490
rect 16776 3488 16896 3490
rect 17639 3488 17684 3516
rect 16672 3479 16730 3485
rect 14476 3448 14504 3476
rect 11572 3420 14504 3448
rect 15473 3451 15531 3457
rect 11572 3408 11578 3420
rect 15473 3417 15485 3451
rect 15519 3448 15531 3451
rect 16500 3448 16528 3479
rect 15519 3420 16528 3448
rect 15519 3417 15531 3420
rect 15473 3411 15531 3417
rect 1486 3380 1492 3392
rect 1447 3352 1492 3380
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 12526 3380 12532 3392
rect 12487 3352 12532 3380
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 13357 3383 13415 3389
rect 13357 3349 13369 3383
rect 13403 3380 13415 3383
rect 15286 3380 15292 3392
rect 13403 3352 15292 3380
rect 13403 3349 13415 3352
rect 13357 3343 13415 3349
rect 15286 3340 15292 3352
rect 15344 3380 15350 3392
rect 15488 3380 15516 3411
rect 15344 3352 15516 3380
rect 15344 3340 15350 3352
rect 15562 3340 15568 3392
rect 15620 3380 15626 3392
rect 15683 3383 15741 3389
rect 15683 3380 15695 3383
rect 15620 3352 15695 3380
rect 15620 3340 15626 3352
rect 15683 3349 15695 3352
rect 15729 3380 15741 3383
rect 16868 3380 16896 3488
rect 17678 3476 17684 3488
rect 17736 3476 17742 3528
rect 17788 3380 17816 3556
rect 19521 3553 19533 3556
rect 19567 3553 19579 3587
rect 19904 3584 19932 3692
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20806 3720 20812 3732
rect 20767 3692 20812 3720
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 21729 3723 21787 3729
rect 21729 3689 21741 3723
rect 21775 3720 21787 3723
rect 22094 3720 22100 3732
rect 21775 3692 22100 3720
rect 21775 3689 21787 3692
rect 21729 3683 21787 3689
rect 22094 3680 22100 3692
rect 22152 3680 22158 3732
rect 23290 3720 23296 3732
rect 23251 3692 23296 3720
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 23658 3680 23664 3732
rect 23716 3720 23722 3732
rect 24397 3723 24455 3729
rect 24397 3720 24409 3723
rect 23716 3692 24409 3720
rect 23716 3680 23722 3692
rect 24397 3689 24409 3692
rect 24443 3689 24455 3723
rect 24397 3683 24455 3689
rect 23106 3612 23112 3664
rect 23164 3652 23170 3664
rect 28445 3655 28503 3661
rect 28445 3652 28457 3655
rect 23164 3624 28457 3652
rect 23164 3612 23170 3624
rect 28445 3621 28457 3624
rect 28491 3621 28503 3655
rect 28445 3615 28503 3621
rect 21818 3584 21824 3596
rect 19904 3556 21824 3584
rect 19521 3547 19579 3553
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18325 3519 18383 3525
rect 18325 3516 18337 3519
rect 17920 3488 18337 3516
rect 17920 3476 17926 3488
rect 18325 3485 18337 3488
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 18966 3476 18972 3528
rect 19024 3516 19030 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 19024 3488 19441 3516
rect 19024 3476 19030 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19948 3519 20006 3525
rect 19948 3516 19960 3519
rect 19429 3479 19487 3485
rect 19628 3488 19960 3516
rect 17954 3408 17960 3460
rect 18012 3448 18018 3460
rect 18601 3451 18659 3457
rect 18601 3448 18613 3451
rect 18012 3420 18613 3448
rect 18012 3408 18018 3420
rect 18601 3417 18613 3420
rect 18647 3448 18659 3451
rect 19628 3448 19656 3488
rect 19948 3485 19960 3488
rect 19994 3516 20006 3519
rect 20898 3516 20904 3528
rect 19994 3488 20760 3516
rect 20859 3488 20904 3516
rect 19994 3485 20006 3488
rect 19948 3479 20006 3485
rect 18647 3420 19656 3448
rect 18647 3417 18659 3420
rect 18601 3411 18659 3417
rect 15729 3352 17816 3380
rect 15729 3349 15741 3352
rect 15683 3343 15741 3349
rect 18046 3340 18052 3392
rect 18104 3380 18110 3392
rect 18417 3383 18475 3389
rect 18417 3380 18429 3383
rect 18104 3352 18429 3380
rect 18104 3340 18110 3352
rect 18417 3349 18429 3352
rect 18463 3349 18475 3383
rect 18417 3343 18475 3349
rect 19889 3383 19947 3389
rect 19889 3349 19901 3383
rect 19935 3380 19947 3383
rect 20530 3380 20536 3392
rect 19935 3352 20536 3380
rect 19935 3349 19947 3352
rect 19889 3343 19947 3349
rect 20530 3340 20536 3352
rect 20588 3380 20594 3392
rect 20625 3383 20683 3389
rect 20625 3380 20637 3383
rect 20588 3352 20637 3380
rect 20588 3340 20594 3352
rect 20625 3349 20637 3352
rect 20671 3349 20683 3383
rect 20732 3380 20760 3488
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 20990 3476 20996 3528
rect 21048 3516 21054 3528
rect 21450 3516 21456 3528
rect 21048 3488 21093 3516
rect 21411 3488 21456 3516
rect 21048 3476 21054 3488
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 21652 3525 21680 3556
rect 21818 3544 21824 3556
rect 21876 3544 21882 3596
rect 22281 3587 22339 3593
rect 22281 3584 22293 3587
rect 22066 3556 22293 3584
rect 21637 3519 21695 3525
rect 21637 3485 21649 3519
rect 21683 3485 21695 3519
rect 21637 3479 21695 3485
rect 21729 3519 21787 3525
rect 21729 3485 21741 3519
rect 21775 3516 21787 3519
rect 21910 3516 21916 3528
rect 21775 3488 21916 3516
rect 21775 3485 21787 3488
rect 21729 3479 21787 3485
rect 21910 3476 21916 3488
rect 21968 3516 21974 3528
rect 22066 3516 22094 3556
rect 22281 3553 22293 3556
rect 22327 3553 22339 3587
rect 22281 3547 22339 3553
rect 23474 3544 23480 3596
rect 23532 3584 23538 3596
rect 23753 3587 23811 3593
rect 23753 3584 23765 3587
rect 23532 3556 23765 3584
rect 23532 3544 23538 3556
rect 23753 3553 23765 3556
rect 23799 3553 23811 3587
rect 23753 3547 23811 3553
rect 21968 3488 22094 3516
rect 22189 3519 22247 3525
rect 21968 3476 21974 3488
rect 22189 3485 22201 3519
rect 22235 3485 22247 3519
rect 22189 3479 22247 3485
rect 22204 3380 22232 3479
rect 22738 3476 22744 3528
rect 22796 3516 22802 3528
rect 22925 3519 22983 3525
rect 22925 3516 22937 3519
rect 22796 3488 22937 3516
rect 22796 3476 22802 3488
rect 22925 3485 22937 3488
rect 22971 3516 22983 3519
rect 23842 3516 23848 3528
rect 22971 3488 23848 3516
rect 22971 3485 22983 3488
rect 22925 3479 22983 3485
rect 23842 3476 23848 3488
rect 23900 3476 23906 3528
rect 23014 3408 23020 3460
rect 23072 3448 23078 3460
rect 23109 3451 23167 3457
rect 23109 3448 23121 3451
rect 23072 3420 23121 3448
rect 23072 3408 23078 3420
rect 23109 3417 23121 3420
rect 23155 3417 23167 3451
rect 28629 3451 28687 3457
rect 28629 3448 28641 3451
rect 23109 3411 23167 3417
rect 27908 3420 28641 3448
rect 20732 3352 22232 3380
rect 20625 3343 20683 3349
rect 27430 3340 27436 3392
rect 27488 3380 27494 3392
rect 27908 3389 27936 3420
rect 28629 3417 28641 3420
rect 28675 3417 28687 3451
rect 28629 3411 28687 3417
rect 27893 3383 27951 3389
rect 27893 3380 27905 3383
rect 27488 3352 27905 3380
rect 27488 3340 27494 3352
rect 27893 3349 27905 3352
rect 27939 3349 27951 3383
rect 27893 3343 27951 3349
rect 1104 3290 29600 3312
rect 1104 3238 8034 3290
rect 8086 3238 8098 3290
rect 8150 3238 8162 3290
rect 8214 3238 8226 3290
rect 8278 3238 8290 3290
rect 8342 3238 15118 3290
rect 15170 3238 15182 3290
rect 15234 3238 15246 3290
rect 15298 3238 15310 3290
rect 15362 3238 15374 3290
rect 15426 3238 22202 3290
rect 22254 3238 22266 3290
rect 22318 3238 22330 3290
rect 22382 3238 22394 3290
rect 22446 3238 22458 3290
rect 22510 3238 29286 3290
rect 29338 3238 29350 3290
rect 29402 3238 29414 3290
rect 29466 3238 29478 3290
rect 29530 3238 29542 3290
rect 29594 3238 29600 3290
rect 1104 3216 29600 3238
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 10321 3179 10379 3185
rect 10321 3176 10333 3179
rect 10100 3148 10333 3176
rect 10100 3136 10106 3148
rect 10321 3145 10333 3148
rect 10367 3145 10379 3179
rect 10321 3139 10379 3145
rect 2406 3068 2412 3120
rect 2464 3108 2470 3120
rect 10336 3108 10364 3139
rect 10594 3136 10600 3188
rect 10652 3176 10658 3188
rect 10873 3179 10931 3185
rect 10873 3176 10885 3179
rect 10652 3148 10885 3176
rect 10652 3136 10658 3148
rect 10873 3145 10885 3148
rect 10919 3145 10931 3179
rect 11514 3176 11520 3188
rect 11475 3148 11520 3176
rect 10873 3139 10931 3145
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 12713 3179 12771 3185
rect 12713 3176 12725 3179
rect 12676 3148 12725 3176
rect 12676 3136 12682 3148
rect 12713 3145 12725 3148
rect 12759 3145 12771 3179
rect 13906 3176 13912 3188
rect 13867 3148 13912 3176
rect 12713 3139 12771 3145
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 14458 3136 14464 3188
rect 14516 3176 14522 3188
rect 14921 3179 14979 3185
rect 14921 3176 14933 3179
rect 14516 3148 14933 3176
rect 14516 3136 14522 3148
rect 14921 3145 14933 3148
rect 14967 3145 14979 3179
rect 14921 3139 14979 3145
rect 17678 3136 17684 3188
rect 17736 3176 17742 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 17736 3148 18061 3176
rect 17736 3136 17742 3148
rect 18049 3145 18061 3148
rect 18095 3176 18107 3179
rect 20717 3179 20775 3185
rect 20717 3176 20729 3179
rect 18095 3148 19196 3176
rect 18095 3145 18107 3148
rect 18049 3139 18107 3145
rect 2464 3080 2774 3108
rect 10336 3080 11928 3108
rect 2464 3068 2470 3080
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 2038 3040 2044 3052
rect 1719 3012 2044 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 2038 3000 2044 3012
rect 2096 3000 2102 3052
rect 2746 2972 2774 3080
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 11900 3049 11928 3080
rect 14090 3068 14096 3120
rect 14148 3108 14154 3120
rect 15105 3111 15163 3117
rect 15105 3108 15117 3111
rect 14148 3080 15117 3108
rect 14148 3068 14154 3080
rect 15105 3077 15117 3080
rect 15151 3077 15163 3111
rect 18966 3108 18972 3120
rect 15105 3071 15163 3077
rect 17236 3080 18972 3108
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 10928 3012 11713 3040
rect 10928 3000 10934 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12526 3040 12532 3052
rect 12023 3012 12532 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 14366 3040 14372 3052
rect 14327 3012 14372 3040
rect 14366 3000 14372 3012
rect 14424 3040 14430 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14424 3012 14841 3040
rect 14424 3000 14430 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 17236 3040 17264 3080
rect 18966 3068 18972 3080
rect 19024 3068 19030 3120
rect 19168 3117 19196 3148
rect 19352 3148 20729 3176
rect 19352 3117 19380 3148
rect 20717 3145 20729 3148
rect 20763 3176 20775 3179
rect 21450 3176 21456 3188
rect 20763 3148 21456 3176
rect 20763 3145 20775 3148
rect 20717 3139 20775 3145
rect 21450 3136 21456 3148
rect 21508 3136 21514 3188
rect 23014 3136 23020 3188
rect 23072 3176 23078 3188
rect 23385 3179 23443 3185
rect 23385 3176 23397 3179
rect 23072 3148 23397 3176
rect 23072 3136 23078 3148
rect 23385 3145 23397 3148
rect 23431 3145 23443 3179
rect 23385 3139 23443 3145
rect 19153 3111 19211 3117
rect 19153 3077 19165 3111
rect 19199 3077 19211 3111
rect 19153 3071 19211 3077
rect 19337 3111 19395 3117
rect 19337 3077 19349 3111
rect 19383 3077 19395 3111
rect 19337 3071 19395 3077
rect 19444 3080 20852 3108
rect 18138 3040 18144 3052
rect 14976 3012 17264 3040
rect 18099 3012 18144 3040
rect 14976 3000 14982 3012
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 18230 3000 18236 3052
rect 18288 3040 18294 3052
rect 19444 3040 19472 3080
rect 20530 3040 20536 3052
rect 18288 3012 19472 3040
rect 20491 3012 20536 3040
rect 18288 3000 18294 3012
rect 20530 3000 20536 3012
rect 20588 3000 20594 3052
rect 20714 3040 20720 3052
rect 20675 3012 20720 3040
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 20824 3040 20852 3080
rect 20990 3068 20996 3120
rect 21048 3108 21054 3120
rect 21269 3111 21327 3117
rect 21269 3108 21281 3111
rect 21048 3080 21281 3108
rect 21048 3068 21054 3080
rect 21269 3077 21281 3080
rect 21315 3108 21327 3111
rect 28445 3111 28503 3117
rect 28445 3108 28457 3111
rect 21315 3080 28457 3108
rect 21315 3077 21327 3080
rect 21269 3071 21327 3077
rect 28445 3077 28457 3080
rect 28491 3077 28503 3111
rect 28445 3071 28503 3077
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 20824 3012 27169 3040
rect 27157 3009 27169 3012
rect 27203 3040 27215 3043
rect 27709 3043 27767 3049
rect 27709 3040 27721 3043
rect 27203 3012 27721 3040
rect 27203 3009 27215 3012
rect 27157 3003 27215 3009
rect 27709 3009 27721 3012
rect 27755 3009 27767 3043
rect 28626 3040 28632 3052
rect 28587 3012 28632 3040
rect 27709 3003 27767 3009
rect 28626 3000 28632 3012
rect 28684 3000 28690 3052
rect 21818 2972 21824 2984
rect 2746 2944 21824 2972
rect 21818 2932 21824 2944
rect 21876 2932 21882 2984
rect 15105 2907 15163 2913
rect 15105 2873 15117 2907
rect 15151 2904 15163 2907
rect 15562 2904 15568 2916
rect 15151 2876 15568 2904
rect 15151 2873 15163 2876
rect 15105 2867 15163 2873
rect 15562 2864 15568 2876
rect 15620 2864 15626 2916
rect 27893 2907 27951 2913
rect 27893 2873 27905 2907
rect 27939 2904 27951 2907
rect 29638 2904 29644 2916
rect 27939 2876 29644 2904
rect 27939 2873 27951 2876
rect 27893 2867 27951 2873
rect 29638 2864 29644 2876
rect 29696 2864 29702 2916
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 72 2808 1501 2836
rect 72 2796 78 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 14090 2836 14096 2848
rect 14051 2808 14096 2836
rect 1489 2799 1547 2805
rect 14090 2796 14096 2808
rect 14148 2796 14154 2848
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 16853 2839 16911 2845
rect 16853 2836 16865 2839
rect 16816 2808 16865 2836
rect 16816 2796 16822 2808
rect 16853 2805 16865 2808
rect 16899 2805 16911 2839
rect 16853 2799 16911 2805
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 19797 2839 19855 2845
rect 19797 2836 19809 2839
rect 19300 2808 19809 2836
rect 19300 2796 19306 2808
rect 19797 2805 19809 2808
rect 19843 2805 19855 2839
rect 19797 2799 19855 2805
rect 1104 2746 29440 2768
rect 1104 2694 4492 2746
rect 4544 2694 4556 2746
rect 4608 2694 4620 2746
rect 4672 2694 4684 2746
rect 4736 2694 4748 2746
rect 4800 2694 11576 2746
rect 11628 2694 11640 2746
rect 11692 2694 11704 2746
rect 11756 2694 11768 2746
rect 11820 2694 11832 2746
rect 11884 2694 18660 2746
rect 18712 2694 18724 2746
rect 18776 2694 18788 2746
rect 18840 2694 18852 2746
rect 18904 2694 18916 2746
rect 18968 2694 25744 2746
rect 25796 2694 25808 2746
rect 25860 2694 25872 2746
rect 25924 2694 25936 2746
rect 25988 2694 26000 2746
rect 26052 2694 29440 2746
rect 1104 2672 29440 2694
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 6730 2632 6736 2644
rect 6595 2604 6736 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14369 2635 14427 2641
rect 14369 2632 14381 2635
rect 14056 2604 14381 2632
rect 14056 2592 14062 2604
rect 14369 2601 14381 2604
rect 14415 2632 14427 2635
rect 14918 2632 14924 2644
rect 14415 2604 14924 2632
rect 14415 2601 14427 2604
rect 14369 2595 14427 2601
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 17221 2635 17279 2641
rect 17221 2601 17233 2635
rect 17267 2632 17279 2635
rect 19610 2632 19616 2644
rect 17267 2604 19616 2632
rect 17267 2601 17279 2604
rect 17221 2595 17279 2601
rect 19610 2592 19616 2604
rect 19668 2592 19674 2644
rect 20898 2632 20904 2644
rect 20859 2604 20904 2632
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 27982 2632 27988 2644
rect 27943 2604 27988 2632
rect 27982 2592 27988 2604
rect 28040 2592 28046 2644
rect 2409 2567 2467 2573
rect 2409 2533 2421 2567
rect 2455 2564 2467 2567
rect 22922 2564 22928 2576
rect 2455 2536 10640 2564
rect 2455 2533 2467 2536
rect 2409 2527 2467 2533
rect 4246 2428 4252 2440
rect 4207 2400 4252 2428
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5828 2400 6377 2428
rect 1581 2363 1639 2369
rect 1581 2329 1593 2363
rect 1627 2360 1639 2363
rect 1946 2360 1952 2372
rect 1627 2332 1952 2360
rect 1627 2329 1639 2332
rect 1581 2323 1639 2329
rect 1946 2320 1952 2332
rect 2004 2360 2010 2372
rect 2133 2363 2191 2369
rect 2133 2360 2145 2363
rect 2004 2332 2145 2360
rect 2004 2320 2010 2332
rect 2133 2329 2145 2332
rect 2179 2329 2191 2363
rect 2133 2323 2191 2329
rect 5828 2304 5856 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8628 2400 8953 2428
rect 8628 2388 8634 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3936 2264 4077 2292
rect 3936 2252 3942 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 5810 2292 5816 2304
rect 5771 2264 5816 2292
rect 4065 2255 4123 2261
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8444 2264 9137 2292
rect 8444 2252 8450 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10505 2295 10563 2301
rect 10505 2292 10517 2295
rect 10376 2264 10517 2292
rect 10376 2252 10382 2264
rect 10505 2261 10517 2264
rect 10551 2261 10563 2295
rect 10612 2292 10640 2536
rect 10704 2536 22928 2564
rect 10704 2437 10732 2536
rect 22922 2524 22928 2536
rect 22980 2524 22986 2576
rect 23569 2567 23627 2573
rect 23569 2533 23581 2567
rect 23615 2564 23627 2567
rect 24026 2564 24032 2576
rect 23615 2536 24032 2564
rect 23615 2533 23627 2536
rect 23569 2527 23627 2533
rect 24026 2524 24032 2536
rect 24084 2524 24090 2576
rect 12713 2499 12771 2505
rect 12713 2465 12725 2499
rect 12759 2496 12771 2499
rect 18230 2496 18236 2508
rect 12759 2468 18092 2496
rect 18191 2468 18236 2496
rect 12759 2465 12771 2468
rect 12713 2459 12771 2465
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2397 10747 2431
rect 14918 2428 14924 2440
rect 14879 2400 14924 2428
rect 10689 2391 10747 2397
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 11885 2363 11943 2369
rect 11885 2329 11897 2363
rect 11931 2360 11943 2363
rect 12250 2360 12256 2372
rect 11931 2332 12256 2360
rect 11931 2329 11943 2332
rect 11885 2323 11943 2329
rect 12250 2320 12256 2332
rect 12308 2360 12314 2372
rect 12437 2363 12495 2369
rect 12437 2360 12449 2363
rect 12308 2332 12449 2360
rect 12308 2320 12314 2332
rect 12437 2329 12449 2332
rect 12483 2329 12495 2363
rect 16574 2360 16580 2372
rect 12437 2323 12495 2329
rect 12544 2332 16580 2360
rect 12544 2292 12572 2332
rect 16574 2320 16580 2332
rect 16632 2320 16638 2372
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16816 2332 17141 2360
rect 16816 2320 16822 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 18064 2360 18092 2468
rect 18230 2456 18236 2468
rect 18288 2456 18294 2508
rect 19150 2456 19156 2508
rect 19208 2496 19214 2508
rect 19521 2499 19579 2505
rect 19208 2468 19380 2496
rect 19208 2456 19214 2468
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 19242 2428 19248 2440
rect 18748 2400 19248 2428
rect 18748 2388 18754 2400
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 19352 2428 19380 2468
rect 19521 2465 19533 2499
rect 19567 2496 19579 2499
rect 19794 2496 19800 2508
rect 19567 2468 19800 2496
rect 19567 2465 19579 2468
rect 19521 2459 19579 2465
rect 19794 2456 19800 2468
rect 19852 2456 19858 2508
rect 25225 2499 25283 2505
rect 25225 2496 25237 2499
rect 19904 2468 25237 2496
rect 19904 2428 19932 2468
rect 25225 2465 25237 2468
rect 25271 2465 25283 2499
rect 25225 2459 25283 2465
rect 20990 2428 20996 2440
rect 19352 2400 19932 2428
rect 20951 2400 20996 2428
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 21818 2428 21824 2440
rect 21779 2400 21824 2428
rect 21818 2388 21824 2400
rect 21876 2388 21882 2440
rect 19886 2360 19892 2372
rect 18064 2332 19892 2360
rect 17129 2323 17187 2329
rect 19886 2320 19892 2332
rect 19944 2320 19950 2372
rect 22833 2363 22891 2369
rect 22833 2329 22845 2363
rect 22879 2360 22891 2363
rect 23198 2360 23204 2372
rect 22879 2332 23204 2360
rect 22879 2329 22891 2332
rect 22833 2323 22891 2329
rect 23198 2320 23204 2332
rect 23256 2360 23262 2372
rect 23385 2363 23443 2369
rect 23385 2360 23397 2363
rect 23256 2332 23397 2360
rect 23256 2320 23262 2332
rect 23385 2329 23397 2332
rect 23431 2329 23443 2363
rect 23385 2323 23443 2329
rect 24765 2363 24823 2369
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 25130 2360 25136 2372
rect 24811 2332 25136 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 25130 2320 25136 2332
rect 25188 2360 25194 2372
rect 25409 2363 25467 2369
rect 25409 2360 25421 2363
rect 25188 2332 25421 2360
rect 25188 2320 25194 2332
rect 25409 2329 25421 2332
rect 25455 2329 25467 2363
rect 25409 2323 25467 2329
rect 27341 2363 27399 2369
rect 27341 2329 27353 2363
rect 27387 2360 27399 2363
rect 27706 2360 27712 2372
rect 27387 2332 27712 2360
rect 27387 2329 27399 2332
rect 27341 2323 27399 2329
rect 27706 2320 27712 2332
rect 27764 2360 27770 2372
rect 27893 2363 27951 2369
rect 27893 2360 27905 2363
rect 27764 2332 27905 2360
rect 27764 2320 27770 2332
rect 27893 2329 27905 2332
rect 27939 2329 27951 2363
rect 27893 2323 27951 2329
rect 10612 2264 12572 2292
rect 10505 2255 10563 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14884 2264 15117 2292
rect 14884 2252 14890 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21324 2264 22017 2292
rect 21324 2252 21330 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 1104 2202 29600 2224
rect 1104 2150 8034 2202
rect 8086 2150 8098 2202
rect 8150 2150 8162 2202
rect 8214 2150 8226 2202
rect 8278 2150 8290 2202
rect 8342 2150 15118 2202
rect 15170 2150 15182 2202
rect 15234 2150 15246 2202
rect 15298 2150 15310 2202
rect 15362 2150 15374 2202
rect 15426 2150 22202 2202
rect 22254 2150 22266 2202
rect 22318 2150 22330 2202
rect 22382 2150 22394 2202
rect 22446 2150 22458 2202
rect 22510 2150 29286 2202
rect 29338 2150 29350 2202
rect 29402 2150 29414 2202
rect 29466 2150 29478 2202
rect 29530 2150 29542 2202
rect 29594 2150 29600 2202
rect 1104 2128 29600 2150
<< via1 >>
rect 8034 30438 8086 30490
rect 8098 30438 8150 30490
rect 8162 30438 8214 30490
rect 8226 30438 8278 30490
rect 8290 30438 8342 30490
rect 15118 30438 15170 30490
rect 15182 30438 15234 30490
rect 15246 30438 15298 30490
rect 15310 30438 15362 30490
rect 15374 30438 15426 30490
rect 22202 30438 22254 30490
rect 22266 30438 22318 30490
rect 22330 30438 22382 30490
rect 22394 30438 22446 30490
rect 22458 30438 22510 30490
rect 29286 30438 29338 30490
rect 29350 30438 29402 30490
rect 29414 30438 29466 30490
rect 29478 30438 29530 30490
rect 29542 30438 29594 30490
rect 664 30268 716 30320
rect 1308 30268 1360 30320
rect 2596 30268 2648 30320
rect 13544 30311 13596 30320
rect 5540 30243 5592 30252
rect 5540 30209 5549 30243
rect 5549 30209 5583 30243
rect 5583 30209 5592 30243
rect 5540 30200 5592 30209
rect 7104 30200 7156 30252
rect 7840 30200 7892 30252
rect 11336 30200 11388 30252
rect 13544 30277 13553 30311
rect 13553 30277 13587 30311
rect 13587 30277 13596 30311
rect 13544 30268 13596 30277
rect 15476 30268 15528 30320
rect 18052 30200 18104 30252
rect 19984 30200 20036 30252
rect 21916 30200 21968 30252
rect 24492 30200 24544 30252
rect 26332 30200 26384 30252
rect 27620 30200 27672 30252
rect 28264 30200 28316 30252
rect 2044 30107 2096 30116
rect 2044 30073 2053 30107
rect 2053 30073 2087 30107
rect 2087 30073 2096 30107
rect 2044 30064 2096 30073
rect 5172 30064 5224 30116
rect 9036 30064 9088 30116
rect 11612 30064 11664 30116
rect 10968 29996 11020 30048
rect 13084 30064 13136 30116
rect 13912 30132 13964 30184
rect 13360 30064 13412 30116
rect 17960 30064 18012 30116
rect 22652 30064 22704 30116
rect 26424 30064 26476 30116
rect 28356 30064 28408 30116
rect 16028 29996 16080 30048
rect 20076 29996 20128 30048
rect 22008 29996 22060 30048
rect 24400 29996 24452 30048
rect 26332 30039 26384 30048
rect 26332 30005 26341 30039
rect 26341 30005 26375 30039
rect 26375 30005 26384 30039
rect 26332 29996 26384 30005
rect 27896 30039 27948 30048
rect 27896 30005 27905 30039
rect 27905 30005 27939 30039
rect 27939 30005 27948 30039
rect 27896 29996 27948 30005
rect 4492 29894 4544 29946
rect 4556 29894 4608 29946
rect 4620 29894 4672 29946
rect 4684 29894 4736 29946
rect 4748 29894 4800 29946
rect 11576 29894 11628 29946
rect 11640 29894 11692 29946
rect 11704 29894 11756 29946
rect 11768 29894 11820 29946
rect 11832 29894 11884 29946
rect 18660 29894 18712 29946
rect 18724 29894 18776 29946
rect 18788 29894 18840 29946
rect 18852 29894 18904 29946
rect 18916 29894 18968 29946
rect 25744 29894 25796 29946
rect 25808 29894 25860 29946
rect 25872 29894 25924 29946
rect 25936 29894 25988 29946
rect 26000 29894 26052 29946
rect 2596 29835 2648 29844
rect 2596 29801 2605 29835
rect 2605 29801 2639 29835
rect 2639 29801 2648 29835
rect 2596 29792 2648 29801
rect 19984 29835 20036 29844
rect 19984 29801 19993 29835
rect 19993 29801 20027 29835
rect 20027 29801 20036 29835
rect 19984 29792 20036 29801
rect 22100 29792 22152 29844
rect 24492 29835 24544 29844
rect 24492 29801 24501 29835
rect 24501 29801 24535 29835
rect 24535 29801 24544 29835
rect 24492 29792 24544 29801
rect 1308 29724 1360 29776
rect 13360 29724 13412 29776
rect 15660 29724 15712 29776
rect 12992 29656 13044 29708
rect 2136 29588 2188 29640
rect 12900 29588 12952 29640
rect 18236 29656 18288 29708
rect 22836 29699 22888 29708
rect 22836 29665 22845 29699
rect 22845 29665 22879 29699
rect 22879 29665 22888 29699
rect 22836 29656 22888 29665
rect 16856 29588 16908 29640
rect 17868 29631 17920 29640
rect 17868 29597 17877 29631
rect 17877 29597 17911 29631
rect 17911 29597 17920 29631
rect 17868 29588 17920 29597
rect 17960 29631 18012 29640
rect 17960 29597 17969 29631
rect 17969 29597 18003 29631
rect 18003 29597 18012 29631
rect 17960 29588 18012 29597
rect 20168 29588 20220 29640
rect 22652 29588 22704 29640
rect 30288 29588 30340 29640
rect 1492 29495 1544 29504
rect 1492 29461 1501 29495
rect 1501 29461 1535 29495
rect 1535 29461 1544 29495
rect 1492 29452 1544 29461
rect 8760 29452 8812 29504
rect 9404 29452 9456 29504
rect 11336 29452 11388 29504
rect 17224 29452 17276 29504
rect 27620 29495 27672 29504
rect 27620 29461 27629 29495
rect 27629 29461 27663 29495
rect 27663 29461 27672 29495
rect 27620 29452 27672 29461
rect 28816 29452 28868 29504
rect 8034 29350 8086 29402
rect 8098 29350 8150 29402
rect 8162 29350 8214 29402
rect 8226 29350 8278 29402
rect 8290 29350 8342 29402
rect 15118 29350 15170 29402
rect 15182 29350 15234 29402
rect 15246 29350 15298 29402
rect 15310 29350 15362 29402
rect 15374 29350 15426 29402
rect 22202 29350 22254 29402
rect 22266 29350 22318 29402
rect 22330 29350 22382 29402
rect 22394 29350 22446 29402
rect 22458 29350 22510 29402
rect 29286 29350 29338 29402
rect 29350 29350 29402 29402
rect 29414 29350 29466 29402
rect 29478 29350 29530 29402
rect 29542 29350 29594 29402
rect 12992 29291 13044 29300
rect 12992 29257 13001 29291
rect 13001 29257 13035 29291
rect 13035 29257 13044 29291
rect 12992 29248 13044 29257
rect 16856 29248 16908 29300
rect 1860 29223 1912 29232
rect 1860 29189 1869 29223
rect 1869 29189 1903 29223
rect 1903 29189 1912 29223
rect 1860 29180 1912 29189
rect 6736 29155 6788 29164
rect 6736 29121 6745 29155
rect 6745 29121 6779 29155
rect 6779 29121 6788 29155
rect 6736 29112 6788 29121
rect 8668 29180 8720 29232
rect 12900 29223 12952 29232
rect 12900 29189 12909 29223
rect 12909 29189 12943 29223
rect 12943 29189 12952 29223
rect 12900 29180 12952 29189
rect 2136 29044 2188 29096
rect 8300 29112 8352 29164
rect 8760 29155 8812 29164
rect 8760 29121 8769 29155
rect 8769 29121 8803 29155
rect 8803 29121 8812 29155
rect 8760 29112 8812 29121
rect 16580 29180 16632 29232
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 16856 29112 16908 29121
rect 16948 29155 17000 29164
rect 16948 29121 16957 29155
rect 16957 29121 16991 29155
rect 16991 29121 17000 29155
rect 16948 29112 17000 29121
rect 17224 29155 17276 29164
rect 17224 29121 17233 29155
rect 17233 29121 17267 29155
rect 17267 29121 17276 29155
rect 17224 29112 17276 29121
rect 17960 29112 18012 29164
rect 19156 29180 19208 29232
rect 8392 29044 8444 29096
rect 10140 29044 10192 29096
rect 12992 29044 13044 29096
rect 15660 29087 15712 29096
rect 4988 28976 5040 29028
rect 5816 28976 5868 29028
rect 9312 28976 9364 29028
rect 12624 28976 12676 29028
rect 9128 28951 9180 28960
rect 9128 28917 9137 28951
rect 9137 28917 9171 28951
rect 9171 28917 9180 28951
rect 9128 28908 9180 28917
rect 10232 28951 10284 28960
rect 10232 28917 10241 28951
rect 10241 28917 10275 28951
rect 10275 28917 10284 28951
rect 10232 28908 10284 28917
rect 13636 28908 13688 28960
rect 15660 29053 15669 29087
rect 15669 29053 15703 29087
rect 15703 29053 15712 29087
rect 15660 29044 15712 29053
rect 17868 29044 17920 29096
rect 19616 29112 19668 29164
rect 21456 29112 21508 29164
rect 22008 29112 22060 29164
rect 22652 29112 22704 29164
rect 15476 28908 15528 28960
rect 19248 28976 19300 29028
rect 19984 28976 20036 29028
rect 28264 29019 28316 29028
rect 28264 28985 28273 29019
rect 28273 28985 28307 29019
rect 28307 28985 28316 29019
rect 28264 28976 28316 28985
rect 19800 28951 19852 28960
rect 19800 28917 19809 28951
rect 19809 28917 19843 28951
rect 19843 28917 19852 28951
rect 19800 28908 19852 28917
rect 21272 28951 21324 28960
rect 21272 28917 21281 28951
rect 21281 28917 21315 28951
rect 21315 28917 21324 28951
rect 21272 28908 21324 28917
rect 22836 28908 22888 28960
rect 23020 28908 23072 28960
rect 23756 28951 23808 28960
rect 23756 28917 23765 28951
rect 23765 28917 23799 28951
rect 23799 28917 23808 28951
rect 23756 28908 23808 28917
rect 4492 28806 4544 28858
rect 4556 28806 4608 28858
rect 4620 28806 4672 28858
rect 4684 28806 4736 28858
rect 4748 28806 4800 28858
rect 11576 28806 11628 28858
rect 11640 28806 11692 28858
rect 11704 28806 11756 28858
rect 11768 28806 11820 28858
rect 11832 28806 11884 28858
rect 18660 28806 18712 28858
rect 18724 28806 18776 28858
rect 18788 28806 18840 28858
rect 18852 28806 18904 28858
rect 18916 28806 18968 28858
rect 25744 28806 25796 28858
rect 25808 28806 25860 28858
rect 25872 28806 25924 28858
rect 25936 28806 25988 28858
rect 26000 28806 26052 28858
rect 1860 28704 1912 28756
rect 6736 28704 6788 28756
rect 7840 28704 7892 28756
rect 8392 28704 8444 28756
rect 10232 28704 10284 28756
rect 19616 28747 19668 28756
rect 19616 28713 19625 28747
rect 19625 28713 19659 28747
rect 19659 28713 19668 28747
rect 19616 28704 19668 28713
rect 8668 28636 8720 28688
rect 16212 28679 16264 28688
rect 16212 28645 16221 28679
rect 16221 28645 16255 28679
rect 16255 28645 16264 28679
rect 16212 28636 16264 28645
rect 19248 28636 19300 28688
rect 9128 28568 9180 28620
rect 12440 28568 12492 28620
rect 13820 28568 13872 28620
rect 14832 28611 14884 28620
rect 14832 28577 14841 28611
rect 14841 28577 14875 28611
rect 14875 28577 14884 28611
rect 14832 28568 14884 28577
rect 18236 28611 18288 28620
rect 18236 28577 18245 28611
rect 18245 28577 18279 28611
rect 18279 28577 18288 28611
rect 18236 28568 18288 28577
rect 19156 28568 19208 28620
rect 21272 28568 21324 28620
rect 21824 28568 21876 28620
rect 5540 28500 5592 28552
rect 7104 28543 7156 28552
rect 7104 28509 7113 28543
rect 7113 28509 7147 28543
rect 7147 28509 7156 28543
rect 7104 28500 7156 28509
rect 8944 28500 8996 28552
rect 9312 28543 9364 28552
rect 9312 28509 9321 28543
rect 9321 28509 9355 28543
rect 9355 28509 9364 28543
rect 9312 28500 9364 28509
rect 11796 28543 11848 28552
rect 11796 28509 11805 28543
rect 11805 28509 11839 28543
rect 11839 28509 11848 28543
rect 11796 28500 11848 28509
rect 12900 28500 12952 28552
rect 13360 28500 13412 28552
rect 14556 28543 14608 28552
rect 14556 28509 14565 28543
rect 14565 28509 14599 28543
rect 14599 28509 14608 28543
rect 14556 28500 14608 28509
rect 15844 28500 15896 28552
rect 16304 28543 16356 28552
rect 16304 28509 16313 28543
rect 16313 28509 16347 28543
rect 16347 28509 16356 28543
rect 16304 28500 16356 28509
rect 8300 28475 8352 28484
rect 8300 28441 8309 28475
rect 8309 28441 8343 28475
rect 8343 28441 8352 28475
rect 8300 28432 8352 28441
rect 9220 28432 9272 28484
rect 16212 28432 16264 28484
rect 16948 28432 17000 28484
rect 22100 28543 22152 28552
rect 22100 28509 22109 28543
rect 22109 28509 22143 28543
rect 22143 28509 22152 28543
rect 22100 28500 22152 28509
rect 23020 28500 23072 28552
rect 6644 28364 6696 28416
rect 10140 28364 10192 28416
rect 11152 28407 11204 28416
rect 11152 28373 11161 28407
rect 11161 28373 11195 28407
rect 11195 28373 11204 28407
rect 11152 28364 11204 28373
rect 12164 28407 12216 28416
rect 12164 28373 12173 28407
rect 12173 28373 12207 28407
rect 12207 28373 12216 28407
rect 12164 28364 12216 28373
rect 12532 28364 12584 28416
rect 12992 28407 13044 28416
rect 12992 28373 13001 28407
rect 13001 28373 13035 28407
rect 13035 28373 13044 28407
rect 12992 28364 13044 28373
rect 19156 28364 19208 28416
rect 23204 28432 23256 28484
rect 23664 28432 23716 28484
rect 19984 28364 20036 28416
rect 21272 28407 21324 28416
rect 21272 28373 21281 28407
rect 21281 28373 21315 28407
rect 21315 28373 21324 28407
rect 21272 28364 21324 28373
rect 22560 28364 22612 28416
rect 23756 28364 23808 28416
rect 24492 28407 24544 28416
rect 24492 28373 24501 28407
rect 24501 28373 24535 28407
rect 24535 28373 24544 28407
rect 24492 28364 24544 28373
rect 8034 28262 8086 28314
rect 8098 28262 8150 28314
rect 8162 28262 8214 28314
rect 8226 28262 8278 28314
rect 8290 28262 8342 28314
rect 15118 28262 15170 28314
rect 15182 28262 15234 28314
rect 15246 28262 15298 28314
rect 15310 28262 15362 28314
rect 15374 28262 15426 28314
rect 22202 28262 22254 28314
rect 22266 28262 22318 28314
rect 22330 28262 22382 28314
rect 22394 28262 22446 28314
rect 22458 28262 22510 28314
rect 29286 28262 29338 28314
rect 29350 28262 29402 28314
rect 29414 28262 29466 28314
rect 29478 28262 29530 28314
rect 29542 28262 29594 28314
rect 7840 28203 7892 28212
rect 7840 28169 7849 28203
rect 7849 28169 7883 28203
rect 7883 28169 7892 28203
rect 7840 28160 7892 28169
rect 8944 28203 8996 28212
rect 8944 28169 8953 28203
rect 8953 28169 8987 28203
rect 8987 28169 8996 28203
rect 8944 28160 8996 28169
rect 10232 28160 10284 28212
rect 15476 28160 15528 28212
rect 15844 28203 15896 28212
rect 15844 28169 15853 28203
rect 15853 28169 15887 28203
rect 15887 28169 15896 28203
rect 15844 28160 15896 28169
rect 19800 28160 19852 28212
rect 20720 28160 20772 28212
rect 12164 28092 12216 28144
rect 7656 28067 7708 28076
rect 7656 28033 7665 28067
rect 7665 28033 7699 28067
rect 7699 28033 7708 28067
rect 7656 28024 7708 28033
rect 9312 28024 9364 28076
rect 11796 28024 11848 28076
rect 12900 28067 12952 28076
rect 12900 28033 12909 28067
rect 12909 28033 12943 28067
rect 12943 28033 12952 28067
rect 12900 28024 12952 28033
rect 12992 28067 13044 28076
rect 12992 28033 13001 28067
rect 13001 28033 13035 28067
rect 13035 28033 13044 28067
rect 14832 28092 14884 28144
rect 12992 28024 13044 28033
rect 9220 27999 9272 28008
rect 9220 27965 9229 27999
rect 9229 27965 9263 27999
rect 9263 27965 9272 27999
rect 9220 27956 9272 27965
rect 10692 27956 10744 28008
rect 13728 28024 13780 28076
rect 14924 28024 14976 28076
rect 21364 28092 21416 28144
rect 21548 28092 21600 28144
rect 16672 27999 16724 28008
rect 7748 27888 7800 27940
rect 16672 27965 16681 27999
rect 16681 27965 16715 27999
rect 16715 27965 16724 27999
rect 16672 27956 16724 27965
rect 19156 28067 19208 28076
rect 19156 28033 19165 28067
rect 19165 28033 19199 28067
rect 19199 28033 19208 28067
rect 20168 28067 20220 28076
rect 19156 28024 19208 28033
rect 20168 28033 20177 28067
rect 20177 28033 20211 28067
rect 20211 28033 20220 28067
rect 20168 28024 20220 28033
rect 21272 28024 21324 28076
rect 22100 28067 22152 28076
rect 22100 28033 22106 28067
rect 22106 28033 22140 28067
rect 22140 28033 22152 28067
rect 22652 28092 22704 28144
rect 23204 28160 23256 28212
rect 24676 28160 24728 28212
rect 23112 28092 23164 28144
rect 24584 28135 24636 28144
rect 22560 28067 22612 28076
rect 22100 28024 22152 28033
rect 22560 28033 22569 28067
rect 22569 28033 22603 28067
rect 22603 28033 22612 28067
rect 22560 28024 22612 28033
rect 23480 28024 23532 28076
rect 23664 28024 23716 28076
rect 24584 28101 24593 28135
rect 24593 28101 24627 28135
rect 24627 28101 24636 28135
rect 24584 28092 24636 28101
rect 28632 28067 28684 28076
rect 28632 28033 28641 28067
rect 28641 28033 28675 28067
rect 28675 28033 28684 28067
rect 28632 28024 28684 28033
rect 19616 27956 19668 28008
rect 24492 27956 24544 28008
rect 21732 27888 21784 27940
rect 10140 27820 10192 27872
rect 11060 27820 11112 27872
rect 13820 27820 13872 27872
rect 18512 27820 18564 27872
rect 19892 27820 19944 27872
rect 20168 27820 20220 27872
rect 23940 27888 23992 27940
rect 26148 27888 26200 27940
rect 22744 27820 22796 27872
rect 23480 27820 23532 27872
rect 24308 27820 24360 27872
rect 4492 27718 4544 27770
rect 4556 27718 4608 27770
rect 4620 27718 4672 27770
rect 4684 27718 4736 27770
rect 4748 27718 4800 27770
rect 11576 27718 11628 27770
rect 11640 27718 11692 27770
rect 11704 27718 11756 27770
rect 11768 27718 11820 27770
rect 11832 27718 11884 27770
rect 18660 27718 18712 27770
rect 18724 27718 18776 27770
rect 18788 27718 18840 27770
rect 18852 27718 18904 27770
rect 18916 27718 18968 27770
rect 25744 27718 25796 27770
rect 25808 27718 25860 27770
rect 25872 27718 25924 27770
rect 25936 27718 25988 27770
rect 26000 27718 26052 27770
rect 12900 27616 12952 27668
rect 14556 27616 14608 27668
rect 14648 27659 14700 27668
rect 14648 27625 14657 27659
rect 14657 27625 14691 27659
rect 14691 27625 14700 27659
rect 19616 27659 19668 27668
rect 14648 27616 14700 27625
rect 19616 27625 19625 27659
rect 19625 27625 19659 27659
rect 19659 27625 19668 27659
rect 19616 27616 19668 27625
rect 25504 27659 25556 27668
rect 10692 27591 10744 27600
rect 10692 27557 10701 27591
rect 10701 27557 10735 27591
rect 10735 27557 10744 27591
rect 10692 27548 10744 27557
rect 15660 27548 15712 27600
rect 19708 27548 19760 27600
rect 21548 27548 21600 27600
rect 21732 27591 21784 27600
rect 21732 27557 21741 27591
rect 21741 27557 21775 27591
rect 21775 27557 21784 27591
rect 21732 27548 21784 27557
rect 10048 27480 10100 27532
rect 11244 27412 11296 27464
rect 13728 27480 13780 27532
rect 19248 27480 19300 27532
rect 25504 27625 25513 27659
rect 25513 27625 25547 27659
rect 25547 27625 25556 27659
rect 25504 27616 25556 27625
rect 12624 27455 12676 27464
rect 12624 27421 12633 27455
rect 12633 27421 12667 27455
rect 12667 27421 12676 27455
rect 12624 27412 12676 27421
rect 13820 27412 13872 27464
rect 16120 27412 16172 27464
rect 19800 27455 19852 27464
rect 19800 27421 19809 27455
rect 19809 27421 19843 27455
rect 19843 27421 19852 27455
rect 19800 27412 19852 27421
rect 19892 27455 19944 27464
rect 19892 27421 19901 27455
rect 19901 27421 19935 27455
rect 19935 27421 19944 27455
rect 19892 27412 19944 27421
rect 10876 27344 10928 27396
rect 11060 27344 11112 27396
rect 12072 27344 12124 27396
rect 20444 27412 20496 27464
rect 24676 27480 24728 27532
rect 23204 27455 23256 27464
rect 23204 27421 23213 27455
rect 23213 27421 23247 27455
rect 23247 27421 23256 27455
rect 23204 27412 23256 27421
rect 23664 27455 23716 27464
rect 23664 27421 23673 27455
rect 23673 27421 23707 27455
rect 23707 27421 23716 27455
rect 23664 27412 23716 27421
rect 24308 27412 24360 27464
rect 24584 27455 24636 27464
rect 24584 27421 24593 27455
rect 24593 27421 24627 27455
rect 24627 27421 24636 27455
rect 24584 27412 24636 27421
rect 25136 27455 25188 27464
rect 25136 27421 25145 27455
rect 25145 27421 25179 27455
rect 25179 27421 25188 27455
rect 25136 27412 25188 27421
rect 25596 27455 25648 27464
rect 25596 27421 25605 27455
rect 25605 27421 25639 27455
rect 25639 27421 25648 27455
rect 25596 27412 25648 27421
rect 8392 27276 8444 27328
rect 9404 27276 9456 27328
rect 11152 27276 11204 27328
rect 15844 27276 15896 27328
rect 16212 27319 16264 27328
rect 16212 27285 16221 27319
rect 16221 27285 16255 27319
rect 16255 27285 16264 27319
rect 16212 27276 16264 27285
rect 19616 27276 19668 27328
rect 20168 27276 20220 27328
rect 20996 27319 21048 27328
rect 20996 27285 21005 27319
rect 21005 27285 21039 27319
rect 21039 27285 21048 27319
rect 20996 27276 21048 27285
rect 22652 27344 22704 27396
rect 8034 27174 8086 27226
rect 8098 27174 8150 27226
rect 8162 27174 8214 27226
rect 8226 27174 8278 27226
rect 8290 27174 8342 27226
rect 15118 27174 15170 27226
rect 15182 27174 15234 27226
rect 15246 27174 15298 27226
rect 15310 27174 15362 27226
rect 15374 27174 15426 27226
rect 22202 27174 22254 27226
rect 22266 27174 22318 27226
rect 22330 27174 22382 27226
rect 22394 27174 22446 27226
rect 22458 27174 22510 27226
rect 29286 27174 29338 27226
rect 29350 27174 29402 27226
rect 29414 27174 29466 27226
rect 29478 27174 29530 27226
rect 29542 27174 29594 27226
rect 7656 27072 7708 27124
rect 1584 26936 1636 26988
rect 5540 26936 5592 26988
rect 8944 26936 8996 26988
rect 10232 26936 10284 26988
rect 11152 27072 11204 27124
rect 11244 27004 11296 27056
rect 12992 27072 13044 27124
rect 11980 27004 12032 27056
rect 12440 27004 12492 27056
rect 7196 26868 7248 26920
rect 11060 26868 11112 26920
rect 11980 26868 12032 26920
rect 12348 26936 12400 26988
rect 12716 26979 12768 26988
rect 12716 26945 12725 26979
rect 12725 26945 12759 26979
rect 12759 26945 12768 26979
rect 12716 26936 12768 26945
rect 15660 27072 15712 27124
rect 15844 27072 15896 27124
rect 19616 27072 19668 27124
rect 20444 27115 20496 27124
rect 14372 27004 14424 27056
rect 16580 27004 16632 27056
rect 16672 27004 16724 27056
rect 19432 27004 19484 27056
rect 20444 27081 20453 27115
rect 20453 27081 20487 27115
rect 20487 27081 20496 27115
rect 20444 27072 20496 27081
rect 24676 27072 24728 27124
rect 25136 27072 25188 27124
rect 20352 27004 20404 27056
rect 21272 27004 21324 27056
rect 23940 27004 23992 27056
rect 25044 27047 25096 27056
rect 25044 27013 25053 27047
rect 25053 27013 25087 27047
rect 25087 27013 25096 27047
rect 25044 27004 25096 27013
rect 15200 26936 15252 26988
rect 15384 26979 15436 26988
rect 15384 26945 15393 26979
rect 15393 26945 15427 26979
rect 15427 26945 15436 26979
rect 15384 26936 15436 26945
rect 15568 26979 15620 26988
rect 15568 26945 15577 26979
rect 15577 26945 15611 26979
rect 15611 26945 15620 26979
rect 15568 26936 15620 26945
rect 19248 26936 19300 26988
rect 19708 26936 19760 26988
rect 20168 26979 20220 26988
rect 20168 26945 20177 26979
rect 20177 26945 20211 26979
rect 20211 26945 20220 26979
rect 20168 26936 20220 26945
rect 20260 26979 20312 26988
rect 20260 26945 20268 26979
rect 20268 26945 20302 26979
rect 20302 26945 20312 26979
rect 20260 26936 20312 26945
rect 22744 26979 22796 26988
rect 1860 26732 1912 26784
rect 5356 26732 5408 26784
rect 8760 26800 8812 26852
rect 10324 26843 10376 26852
rect 10324 26809 10333 26843
rect 10333 26809 10367 26843
rect 10367 26809 10376 26843
rect 15016 26868 15068 26920
rect 20904 26868 20956 26920
rect 22744 26945 22753 26979
rect 22753 26945 22787 26979
rect 22787 26945 22796 26979
rect 22744 26936 22796 26945
rect 24860 26979 24912 26988
rect 21272 26911 21324 26920
rect 21272 26877 21281 26911
rect 21281 26877 21315 26911
rect 21315 26877 21324 26911
rect 21272 26868 21324 26877
rect 24308 26911 24360 26920
rect 24308 26877 24317 26911
rect 24317 26877 24351 26911
rect 24351 26877 24360 26911
rect 24308 26868 24360 26877
rect 24860 26945 24869 26979
rect 24869 26945 24903 26979
rect 24903 26945 24912 26979
rect 24860 26936 24912 26945
rect 26148 26979 26200 26988
rect 24584 26868 24636 26920
rect 26148 26945 26157 26979
rect 26157 26945 26191 26979
rect 26191 26945 26200 26979
rect 26148 26936 26200 26945
rect 10324 26800 10376 26809
rect 14832 26800 14884 26852
rect 8300 26775 8352 26784
rect 8300 26741 8309 26775
rect 8309 26741 8343 26775
rect 8343 26741 8352 26775
rect 8300 26732 8352 26741
rect 10876 26775 10928 26784
rect 10876 26741 10885 26775
rect 10885 26741 10919 26775
rect 10919 26741 10928 26775
rect 10876 26732 10928 26741
rect 12808 26732 12860 26784
rect 14096 26775 14148 26784
rect 14096 26741 14105 26775
rect 14105 26741 14139 26775
rect 14139 26741 14148 26775
rect 14096 26732 14148 26741
rect 15292 26732 15344 26784
rect 19616 26800 19668 26852
rect 17132 26775 17184 26784
rect 17132 26741 17141 26775
rect 17141 26741 17175 26775
rect 17175 26741 17184 26775
rect 17132 26732 17184 26741
rect 18144 26732 18196 26784
rect 18420 26732 18472 26784
rect 19064 26732 19116 26784
rect 21548 26732 21600 26784
rect 22192 26800 22244 26852
rect 22376 26732 22428 26784
rect 22560 26775 22612 26784
rect 22560 26741 22569 26775
rect 22569 26741 22603 26775
rect 22603 26741 22612 26775
rect 22560 26732 22612 26741
rect 23296 26775 23348 26784
rect 23296 26741 23305 26775
rect 23305 26741 23339 26775
rect 23339 26741 23348 26775
rect 23296 26732 23348 26741
rect 24308 26732 24360 26784
rect 25136 26732 25188 26784
rect 28632 26775 28684 26784
rect 28632 26741 28641 26775
rect 28641 26741 28675 26775
rect 28675 26741 28684 26775
rect 28632 26732 28684 26741
rect 4492 26630 4544 26682
rect 4556 26630 4608 26682
rect 4620 26630 4672 26682
rect 4684 26630 4736 26682
rect 4748 26630 4800 26682
rect 11576 26630 11628 26682
rect 11640 26630 11692 26682
rect 11704 26630 11756 26682
rect 11768 26630 11820 26682
rect 11832 26630 11884 26682
rect 18660 26630 18712 26682
rect 18724 26630 18776 26682
rect 18788 26630 18840 26682
rect 18852 26630 18904 26682
rect 18916 26630 18968 26682
rect 25744 26630 25796 26682
rect 25808 26630 25860 26682
rect 25872 26630 25924 26682
rect 25936 26630 25988 26682
rect 26000 26630 26052 26682
rect 1584 26571 1636 26580
rect 1584 26537 1593 26571
rect 1593 26537 1627 26571
rect 1627 26537 1636 26571
rect 1584 26528 1636 26537
rect 5540 26571 5592 26580
rect 5540 26537 5549 26571
rect 5549 26537 5583 26571
rect 5583 26537 5592 26571
rect 5540 26528 5592 26537
rect 7104 26571 7156 26580
rect 7104 26537 7113 26571
rect 7113 26537 7147 26571
rect 7147 26537 7156 26571
rect 7104 26528 7156 26537
rect 7748 26528 7800 26580
rect 11980 26571 12032 26580
rect 11980 26537 11989 26571
rect 11989 26537 12023 26571
rect 12023 26537 12032 26571
rect 11980 26528 12032 26537
rect 12348 26528 12400 26580
rect 14372 26528 14424 26580
rect 15200 26571 15252 26580
rect 15200 26537 15209 26571
rect 15209 26537 15243 26571
rect 15243 26537 15252 26571
rect 15200 26528 15252 26537
rect 16304 26528 16356 26580
rect 5724 26460 5776 26512
rect 10048 26460 10100 26512
rect 5080 26367 5132 26376
rect 5080 26333 5089 26367
rect 5089 26333 5123 26367
rect 5123 26333 5132 26367
rect 5080 26324 5132 26333
rect 5540 26367 5592 26376
rect 5540 26333 5549 26367
rect 5549 26333 5583 26367
rect 5583 26333 5592 26367
rect 5540 26324 5592 26333
rect 5724 26367 5776 26376
rect 5724 26333 5733 26367
rect 5733 26333 5767 26367
rect 5767 26333 5776 26367
rect 5724 26324 5776 26333
rect 7012 26367 7064 26376
rect 7012 26333 7021 26367
rect 7021 26333 7055 26367
rect 7055 26333 7064 26367
rect 7012 26324 7064 26333
rect 8300 26392 8352 26444
rect 8484 26392 8536 26444
rect 8392 26324 8444 26376
rect 10876 26392 10928 26444
rect 11244 26435 11296 26444
rect 11244 26401 11253 26435
rect 11253 26401 11287 26435
rect 11287 26401 11296 26435
rect 11244 26392 11296 26401
rect 12348 26392 12400 26444
rect 5356 26256 5408 26308
rect 9864 26256 9916 26308
rect 7840 26188 7892 26240
rect 8300 26231 8352 26240
rect 8300 26197 8309 26231
rect 8309 26197 8343 26231
rect 8343 26197 8352 26231
rect 8300 26188 8352 26197
rect 10508 26324 10560 26376
rect 10232 26299 10284 26308
rect 10232 26265 10237 26299
rect 10237 26265 10271 26299
rect 10271 26265 10284 26299
rect 11520 26324 11572 26376
rect 12256 26367 12308 26376
rect 12256 26333 12265 26367
rect 12265 26333 12299 26367
rect 12299 26333 12308 26367
rect 12716 26460 12768 26512
rect 19800 26528 19852 26580
rect 20996 26571 21048 26580
rect 20996 26537 21005 26571
rect 21005 26537 21039 26571
rect 21039 26537 21048 26571
rect 20996 26528 21048 26537
rect 22376 26528 22428 26580
rect 23572 26528 23624 26580
rect 23664 26528 23716 26580
rect 17408 26460 17460 26512
rect 18328 26460 18380 26512
rect 18972 26460 19024 26512
rect 15568 26392 15620 26444
rect 19432 26460 19484 26512
rect 20352 26460 20404 26512
rect 21548 26460 21600 26512
rect 23112 26503 23164 26512
rect 12256 26324 12308 26333
rect 12808 26324 12860 26376
rect 10232 26256 10284 26265
rect 12716 26256 12768 26308
rect 10416 26188 10468 26240
rect 12256 26188 12308 26240
rect 15292 26324 15344 26376
rect 15660 26324 15712 26376
rect 15844 26324 15896 26376
rect 16672 26367 16724 26376
rect 16672 26333 16681 26367
rect 16681 26333 16715 26367
rect 16715 26333 16724 26367
rect 16672 26324 16724 26333
rect 14096 26299 14148 26308
rect 14096 26265 14105 26299
rect 14105 26265 14139 26299
rect 14139 26265 14148 26299
rect 14096 26256 14148 26265
rect 14280 26299 14332 26308
rect 14280 26265 14289 26299
rect 14289 26265 14323 26299
rect 14323 26265 14332 26299
rect 14280 26256 14332 26265
rect 13912 26188 13964 26240
rect 16580 26256 16632 26308
rect 16948 26367 17000 26376
rect 16948 26333 16957 26367
rect 16957 26333 16991 26367
rect 16991 26333 17000 26367
rect 17132 26367 17184 26376
rect 16948 26324 17000 26333
rect 17132 26333 17141 26367
rect 17141 26333 17175 26367
rect 17175 26333 17184 26367
rect 17132 26324 17184 26333
rect 18144 26256 18196 26308
rect 15660 26188 15712 26240
rect 16212 26188 16264 26240
rect 18328 26367 18380 26376
rect 18328 26333 18337 26367
rect 18337 26333 18371 26367
rect 18371 26333 18380 26367
rect 18328 26324 18380 26333
rect 19064 26324 19116 26376
rect 18880 26256 18932 26308
rect 18972 26256 19024 26308
rect 19892 26392 19944 26444
rect 23112 26469 23121 26503
rect 23121 26469 23155 26503
rect 23155 26469 23164 26503
rect 23112 26460 23164 26469
rect 19616 26367 19668 26376
rect 19616 26333 19625 26367
rect 19625 26333 19659 26367
rect 19659 26333 19668 26367
rect 19616 26324 19668 26333
rect 19800 26367 19852 26376
rect 19800 26333 19814 26367
rect 19814 26333 19848 26367
rect 19848 26333 19852 26367
rect 20444 26367 20496 26376
rect 19800 26324 19852 26333
rect 20444 26333 20453 26367
rect 20453 26333 20487 26367
rect 20487 26333 20496 26367
rect 20444 26324 20496 26333
rect 20812 26367 20864 26376
rect 20812 26333 20821 26367
rect 20821 26333 20855 26367
rect 20855 26333 20864 26367
rect 20812 26324 20864 26333
rect 19708 26299 19760 26308
rect 19708 26265 19717 26299
rect 19717 26265 19751 26299
rect 19751 26265 19760 26299
rect 19708 26256 19760 26265
rect 22192 26392 22244 26444
rect 24860 26392 24912 26444
rect 24492 26324 24544 26376
rect 26148 26392 26200 26444
rect 19248 26188 19300 26240
rect 25964 26367 26016 26376
rect 25964 26333 25973 26367
rect 25973 26333 26007 26367
rect 26007 26333 26016 26367
rect 25964 26324 26016 26333
rect 28356 26256 28408 26308
rect 28632 26299 28684 26308
rect 28632 26265 28641 26299
rect 28641 26265 28675 26299
rect 28675 26265 28684 26299
rect 28632 26256 28684 26265
rect 21364 26188 21416 26240
rect 25596 26188 25648 26240
rect 8034 26086 8086 26138
rect 8098 26086 8150 26138
rect 8162 26086 8214 26138
rect 8226 26086 8278 26138
rect 8290 26086 8342 26138
rect 15118 26086 15170 26138
rect 15182 26086 15234 26138
rect 15246 26086 15298 26138
rect 15310 26086 15362 26138
rect 15374 26086 15426 26138
rect 22202 26086 22254 26138
rect 22266 26086 22318 26138
rect 22330 26086 22382 26138
rect 22394 26086 22446 26138
rect 22458 26086 22510 26138
rect 29286 26086 29338 26138
rect 29350 26086 29402 26138
rect 29414 26086 29466 26138
rect 29478 26086 29530 26138
rect 29542 26086 29594 26138
rect 5080 25984 5132 26036
rect 7012 25984 7064 26036
rect 7196 26027 7248 26036
rect 7196 25993 7205 26027
rect 7205 25993 7239 26027
rect 7239 25993 7248 26027
rect 7196 25984 7248 25993
rect 8760 26027 8812 26036
rect 8760 25993 8769 26027
rect 8769 25993 8803 26027
rect 8803 25993 8812 26027
rect 8760 25984 8812 25993
rect 9864 25984 9916 26036
rect 10508 25984 10560 26036
rect 11520 26027 11572 26036
rect 11520 25993 11529 26027
rect 11529 25993 11563 26027
rect 11563 25993 11572 26027
rect 11520 25984 11572 25993
rect 13360 26027 13412 26036
rect 13360 25993 13369 26027
rect 13369 25993 13403 26027
rect 13403 25993 13412 26027
rect 13360 25984 13412 25993
rect 13912 25984 13964 26036
rect 14280 25984 14332 26036
rect 15016 26027 15068 26036
rect 15016 25993 15025 26027
rect 15025 25993 15059 26027
rect 15059 25993 15068 26027
rect 15016 25984 15068 25993
rect 19248 25984 19300 26036
rect 20260 25984 20312 26036
rect 20812 25984 20864 26036
rect 23572 25984 23624 26036
rect 4344 25891 4396 25900
rect 4344 25857 4353 25891
rect 4353 25857 4387 25891
rect 4387 25857 4396 25891
rect 4344 25848 4396 25857
rect 5080 25848 5132 25900
rect 5264 25848 5316 25900
rect 5632 25891 5684 25900
rect 5632 25857 5641 25891
rect 5641 25857 5675 25891
rect 5675 25857 5684 25891
rect 5632 25848 5684 25857
rect 4252 25823 4304 25832
rect 4252 25789 4261 25823
rect 4261 25789 4295 25823
rect 4295 25789 4304 25823
rect 4252 25780 4304 25789
rect 6736 25823 6788 25832
rect 6736 25789 6745 25823
rect 6745 25789 6779 25823
rect 6779 25789 6788 25823
rect 6736 25780 6788 25789
rect 7012 25891 7064 25900
rect 7012 25857 7021 25891
rect 7021 25857 7055 25891
rect 7055 25857 7064 25891
rect 7012 25848 7064 25857
rect 7196 25848 7248 25900
rect 7840 25891 7892 25900
rect 7840 25857 7849 25891
rect 7849 25857 7883 25891
rect 7883 25857 7892 25891
rect 7840 25848 7892 25857
rect 7932 25848 7984 25900
rect 10968 25916 11020 25968
rect 8392 25848 8444 25900
rect 8668 25891 8720 25900
rect 8668 25857 8677 25891
rect 8677 25857 8711 25891
rect 8711 25857 8720 25891
rect 8668 25848 8720 25857
rect 9220 25848 9272 25900
rect 10416 25891 10468 25900
rect 10416 25857 10425 25891
rect 10425 25857 10459 25891
rect 10459 25857 10468 25891
rect 10416 25848 10468 25857
rect 12072 25916 12124 25968
rect 12624 25916 12676 25968
rect 14004 25916 14056 25968
rect 12532 25848 12584 25900
rect 14096 25848 14148 25900
rect 14372 25891 14424 25900
rect 14372 25857 14381 25891
rect 14381 25857 14415 25891
rect 14415 25857 14424 25891
rect 14372 25848 14424 25857
rect 14464 25848 14516 25900
rect 16764 25916 16816 25968
rect 18328 25916 18380 25968
rect 18880 25916 18932 25968
rect 20444 25916 20496 25968
rect 15292 25891 15344 25900
rect 15292 25857 15301 25891
rect 15301 25857 15335 25891
rect 15335 25857 15344 25891
rect 15292 25848 15344 25857
rect 15568 25891 15620 25900
rect 5540 25712 5592 25764
rect 8208 25712 8260 25764
rect 10232 25712 10284 25764
rect 12164 25780 12216 25832
rect 14832 25780 14884 25832
rect 15568 25857 15576 25891
rect 15576 25857 15610 25891
rect 15610 25857 15620 25891
rect 15568 25848 15620 25857
rect 19156 25848 19208 25900
rect 17224 25823 17276 25832
rect 15384 25712 15436 25764
rect 6828 25687 6880 25696
rect 6828 25653 6837 25687
rect 6837 25653 6871 25687
rect 6871 25653 6880 25687
rect 6828 25644 6880 25653
rect 12256 25644 12308 25696
rect 12900 25644 12952 25696
rect 17224 25789 17233 25823
rect 17233 25789 17267 25823
rect 17267 25789 17276 25823
rect 17224 25780 17276 25789
rect 18052 25780 18104 25832
rect 19708 25848 19760 25900
rect 21364 25916 21416 25968
rect 20904 25891 20956 25900
rect 20904 25857 20913 25891
rect 20913 25857 20947 25891
rect 20947 25857 20956 25891
rect 20904 25848 20956 25857
rect 26148 25984 26200 26036
rect 24952 25916 25004 25968
rect 25964 25916 26016 25968
rect 26884 25916 26936 25968
rect 19892 25780 19944 25832
rect 16764 25755 16816 25764
rect 16764 25721 16773 25755
rect 16773 25721 16807 25755
rect 16807 25721 16816 25755
rect 16764 25712 16816 25721
rect 19800 25712 19852 25764
rect 22744 25712 22796 25764
rect 23296 25712 23348 25764
rect 27712 25712 27764 25764
rect 18236 25644 18288 25696
rect 26148 25644 26200 25696
rect 27620 25687 27672 25696
rect 27620 25653 27629 25687
rect 27629 25653 27663 25687
rect 27663 25653 27672 25687
rect 27620 25644 27672 25653
rect 28540 25644 28592 25696
rect 4492 25542 4544 25594
rect 4556 25542 4608 25594
rect 4620 25542 4672 25594
rect 4684 25542 4736 25594
rect 4748 25542 4800 25594
rect 11576 25542 11628 25594
rect 11640 25542 11692 25594
rect 11704 25542 11756 25594
rect 11768 25542 11820 25594
rect 11832 25542 11884 25594
rect 18660 25542 18712 25594
rect 18724 25542 18776 25594
rect 18788 25542 18840 25594
rect 18852 25542 18904 25594
rect 18916 25542 18968 25594
rect 25744 25542 25796 25594
rect 25808 25542 25860 25594
rect 25872 25542 25924 25594
rect 25936 25542 25988 25594
rect 26000 25542 26052 25594
rect 4252 25440 4304 25492
rect 5264 25483 5316 25492
rect 5264 25449 5273 25483
rect 5273 25449 5307 25483
rect 5307 25449 5316 25483
rect 5264 25440 5316 25449
rect 7012 25440 7064 25492
rect 8208 25483 8260 25492
rect 8208 25449 8217 25483
rect 8217 25449 8251 25483
rect 8251 25449 8260 25483
rect 8208 25440 8260 25449
rect 14096 25440 14148 25492
rect 15568 25440 15620 25492
rect 16120 25440 16172 25492
rect 17408 25483 17460 25492
rect 17408 25449 17417 25483
rect 17417 25449 17451 25483
rect 17451 25449 17460 25483
rect 17408 25440 17460 25449
rect 18236 25440 18288 25492
rect 19248 25483 19300 25492
rect 19248 25449 19257 25483
rect 19257 25449 19291 25483
rect 19291 25449 19300 25483
rect 19248 25440 19300 25449
rect 20904 25440 20956 25492
rect 21364 25440 21416 25492
rect 23112 25440 23164 25492
rect 23296 25440 23348 25492
rect 26884 25483 26936 25492
rect 26884 25449 26893 25483
rect 26893 25449 26927 25483
rect 26927 25449 26936 25483
rect 26884 25440 26936 25449
rect 27620 25440 27672 25492
rect 28448 25440 28500 25492
rect 7748 25304 7800 25356
rect 4620 25279 4672 25288
rect 4620 25245 4629 25279
rect 4629 25245 4663 25279
rect 4663 25245 4672 25279
rect 4620 25236 4672 25245
rect 5080 25279 5132 25288
rect 5080 25245 5089 25279
rect 5089 25245 5123 25279
rect 5123 25245 5132 25279
rect 5080 25236 5132 25245
rect 5264 25279 5316 25288
rect 5264 25245 5273 25279
rect 5273 25245 5307 25279
rect 5307 25245 5316 25279
rect 5264 25236 5316 25245
rect 6828 25236 6880 25288
rect 7840 25279 7892 25288
rect 7196 25168 7248 25220
rect 7840 25245 7849 25279
rect 7849 25245 7883 25279
rect 7883 25245 7892 25279
rect 7840 25236 7892 25245
rect 8668 25304 8720 25356
rect 16672 25304 16724 25356
rect 9312 25236 9364 25288
rect 12164 25279 12216 25288
rect 12164 25245 12173 25279
rect 12173 25245 12207 25279
rect 12207 25245 12216 25279
rect 12164 25236 12216 25245
rect 13544 25236 13596 25288
rect 10416 25211 10468 25220
rect 10416 25177 10425 25211
rect 10425 25177 10459 25211
rect 10459 25177 10468 25211
rect 10416 25168 10468 25177
rect 12256 25168 12308 25220
rect 5080 25100 5132 25152
rect 6460 25100 6512 25152
rect 6736 25100 6788 25152
rect 10876 25100 10928 25152
rect 12532 25100 12584 25152
rect 13912 25100 13964 25152
rect 15660 25236 15712 25288
rect 25044 25372 25096 25424
rect 19524 25236 19576 25288
rect 22008 25304 22060 25356
rect 19800 25236 19852 25288
rect 22836 25304 22888 25356
rect 22560 25279 22612 25288
rect 17684 25168 17736 25220
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 22560 25236 22612 25245
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 25136 25236 25188 25288
rect 25688 25279 25740 25288
rect 25688 25245 25697 25279
rect 25697 25245 25731 25279
rect 25731 25245 25740 25279
rect 25688 25236 25740 25245
rect 26148 25304 26200 25356
rect 20996 25168 21048 25220
rect 21272 25168 21324 25220
rect 23388 25168 23440 25220
rect 25596 25168 25648 25220
rect 26240 25236 26292 25288
rect 16396 25100 16448 25152
rect 18236 25100 18288 25152
rect 22928 25100 22980 25152
rect 28264 25100 28316 25152
rect 8034 24998 8086 25050
rect 8098 24998 8150 25050
rect 8162 24998 8214 25050
rect 8226 24998 8278 25050
rect 8290 24998 8342 25050
rect 15118 24998 15170 25050
rect 15182 24998 15234 25050
rect 15246 24998 15298 25050
rect 15310 24998 15362 25050
rect 15374 24998 15426 25050
rect 22202 24998 22254 25050
rect 22266 24998 22318 25050
rect 22330 24998 22382 25050
rect 22394 24998 22446 25050
rect 22458 24998 22510 25050
rect 29286 24998 29338 25050
rect 29350 24998 29402 25050
rect 29414 24998 29466 25050
rect 29478 24998 29530 25050
rect 29542 24998 29594 25050
rect 4988 24896 5040 24948
rect 5172 24896 5224 24948
rect 7932 24896 7984 24948
rect 10876 24896 10928 24948
rect 14832 24939 14884 24948
rect 14832 24905 14841 24939
rect 14841 24905 14875 24939
rect 14875 24905 14884 24939
rect 14832 24896 14884 24905
rect 22560 24896 22612 24948
rect 25688 24896 25740 24948
rect 1400 24803 1452 24812
rect 1400 24769 1409 24803
rect 1409 24769 1443 24803
rect 1443 24769 1452 24803
rect 1400 24760 1452 24769
rect 4896 24760 4948 24812
rect 5264 24760 5316 24812
rect 7840 24828 7892 24880
rect 7748 24760 7800 24812
rect 8208 24803 8260 24812
rect 8208 24769 8217 24803
rect 8217 24769 8251 24803
rect 8251 24769 8260 24803
rect 8208 24760 8260 24769
rect 4620 24692 4672 24744
rect 5080 24692 5132 24744
rect 11428 24692 11480 24744
rect 9496 24624 9548 24676
rect 12808 24760 12860 24812
rect 13268 24760 13320 24812
rect 15476 24828 15528 24880
rect 22928 24828 22980 24880
rect 13912 24803 13964 24812
rect 13912 24769 13921 24803
rect 13921 24769 13955 24803
rect 13955 24769 13964 24803
rect 21824 24803 21876 24812
rect 13912 24760 13964 24769
rect 21824 24769 21833 24803
rect 21833 24769 21867 24803
rect 21867 24769 21876 24803
rect 21824 24760 21876 24769
rect 23388 24803 23440 24812
rect 23388 24769 23397 24803
rect 23397 24769 23431 24803
rect 23431 24769 23440 24803
rect 23388 24760 23440 24769
rect 24952 24760 25004 24812
rect 13360 24692 13412 24744
rect 14004 24735 14056 24744
rect 14004 24701 14013 24735
rect 14013 24701 14047 24735
rect 14047 24701 14056 24735
rect 14004 24692 14056 24701
rect 25320 24692 25372 24744
rect 1584 24599 1636 24608
rect 1584 24565 1593 24599
rect 1593 24565 1627 24599
rect 1627 24565 1636 24599
rect 1584 24556 1636 24565
rect 5540 24556 5592 24608
rect 7196 24556 7248 24608
rect 8852 24556 8904 24608
rect 10048 24556 10100 24608
rect 14740 24624 14792 24676
rect 17224 24556 17276 24608
rect 19064 24556 19116 24608
rect 19800 24556 19852 24608
rect 24216 24556 24268 24608
rect 25688 24760 25740 24812
rect 25596 24556 25648 24608
rect 26976 24599 27028 24608
rect 26976 24565 26985 24599
rect 26985 24565 27019 24599
rect 27019 24565 27028 24599
rect 26976 24556 27028 24565
rect 28540 24556 28592 24608
rect 4492 24454 4544 24506
rect 4556 24454 4608 24506
rect 4620 24454 4672 24506
rect 4684 24454 4736 24506
rect 4748 24454 4800 24506
rect 11576 24454 11628 24506
rect 11640 24454 11692 24506
rect 11704 24454 11756 24506
rect 11768 24454 11820 24506
rect 11832 24454 11884 24506
rect 18660 24454 18712 24506
rect 18724 24454 18776 24506
rect 18788 24454 18840 24506
rect 18852 24454 18904 24506
rect 18916 24454 18968 24506
rect 25744 24454 25796 24506
rect 25808 24454 25860 24506
rect 25872 24454 25924 24506
rect 25936 24454 25988 24506
rect 26000 24454 26052 24506
rect 1400 24395 1452 24404
rect 1400 24361 1409 24395
rect 1409 24361 1443 24395
rect 1443 24361 1452 24395
rect 1400 24352 1452 24361
rect 1584 24352 1636 24404
rect 10048 24352 10100 24404
rect 5632 24327 5684 24336
rect 5632 24293 5641 24327
rect 5641 24293 5675 24327
rect 5675 24293 5684 24327
rect 5632 24284 5684 24293
rect 11428 24352 11480 24404
rect 12532 24395 12584 24404
rect 12532 24361 12541 24395
rect 12541 24361 12575 24395
rect 12575 24361 12584 24395
rect 12532 24352 12584 24361
rect 19248 24352 19300 24404
rect 23756 24395 23808 24404
rect 23756 24361 23765 24395
rect 23765 24361 23799 24395
rect 23799 24361 23808 24395
rect 23756 24352 23808 24361
rect 27896 24352 27948 24404
rect 4160 24148 4212 24200
rect 4344 24148 4396 24200
rect 4896 24191 4948 24200
rect 4896 24157 4905 24191
rect 4905 24157 4939 24191
rect 4939 24157 4948 24191
rect 4896 24148 4948 24157
rect 5080 24191 5132 24200
rect 5080 24157 5089 24191
rect 5089 24157 5123 24191
rect 5123 24157 5132 24191
rect 5080 24148 5132 24157
rect 5540 24191 5592 24200
rect 5540 24157 5549 24191
rect 5549 24157 5583 24191
rect 5583 24157 5592 24191
rect 5540 24148 5592 24157
rect 4620 24080 4672 24132
rect 8852 24148 8904 24200
rect 9036 24148 9088 24200
rect 12716 24216 12768 24268
rect 9312 24191 9364 24200
rect 9312 24157 9321 24191
rect 9321 24157 9355 24191
rect 9355 24157 9364 24191
rect 9312 24148 9364 24157
rect 10232 24148 10284 24200
rect 12992 24148 13044 24200
rect 14004 24148 14056 24200
rect 4252 24012 4304 24064
rect 6828 24012 6880 24064
rect 9956 24080 10008 24132
rect 10416 24080 10468 24132
rect 12532 24080 12584 24132
rect 13912 24080 13964 24132
rect 18328 24216 18380 24268
rect 22008 24216 22060 24268
rect 19064 24148 19116 24200
rect 19800 24148 19852 24200
rect 21824 24148 21876 24200
rect 22744 24191 22796 24200
rect 22744 24157 22748 24191
rect 22748 24157 22782 24191
rect 22782 24157 22796 24191
rect 22744 24148 22796 24157
rect 25412 24284 25464 24336
rect 23572 24216 23624 24268
rect 24952 24216 25004 24268
rect 25228 24259 25280 24268
rect 25228 24225 25237 24259
rect 25237 24225 25271 24259
rect 25271 24225 25280 24259
rect 25228 24216 25280 24225
rect 26240 24216 26292 24268
rect 23204 24191 23256 24200
rect 23204 24157 23213 24191
rect 23213 24157 23247 24191
rect 23247 24157 23256 24191
rect 23204 24148 23256 24157
rect 25320 24148 25372 24200
rect 25596 24148 25648 24200
rect 26148 24148 26200 24200
rect 8208 24012 8260 24064
rect 9588 24012 9640 24064
rect 10692 24012 10744 24064
rect 20904 24080 20956 24132
rect 15016 24012 15068 24064
rect 17224 24012 17276 24064
rect 19984 24012 20036 24064
rect 22100 24055 22152 24064
rect 22100 24021 22109 24055
rect 22109 24021 22143 24055
rect 22143 24021 22152 24055
rect 24584 24080 24636 24132
rect 24860 24080 24912 24132
rect 25136 24123 25188 24132
rect 25136 24089 25145 24123
rect 25145 24089 25179 24123
rect 25179 24089 25188 24123
rect 25136 24080 25188 24089
rect 22100 24012 22152 24021
rect 27804 24012 27856 24064
rect 28540 24012 28592 24064
rect 28724 24055 28776 24064
rect 28724 24021 28733 24055
rect 28733 24021 28767 24055
rect 28767 24021 28776 24055
rect 28724 24012 28776 24021
rect 8034 23910 8086 23962
rect 8098 23910 8150 23962
rect 8162 23910 8214 23962
rect 8226 23910 8278 23962
rect 8290 23910 8342 23962
rect 15118 23910 15170 23962
rect 15182 23910 15234 23962
rect 15246 23910 15298 23962
rect 15310 23910 15362 23962
rect 15374 23910 15426 23962
rect 22202 23910 22254 23962
rect 22266 23910 22318 23962
rect 22330 23910 22382 23962
rect 22394 23910 22446 23962
rect 22458 23910 22510 23962
rect 29286 23910 29338 23962
rect 29350 23910 29402 23962
rect 29414 23910 29466 23962
rect 29478 23910 29530 23962
rect 29542 23910 29594 23962
rect 4620 23851 4672 23860
rect 4620 23817 4629 23851
rect 4629 23817 4663 23851
rect 4663 23817 4672 23851
rect 4620 23808 4672 23817
rect 6552 23808 6604 23860
rect 9036 23851 9088 23860
rect 9036 23817 9045 23851
rect 9045 23817 9079 23851
rect 9079 23817 9088 23851
rect 9036 23808 9088 23817
rect 10232 23851 10284 23860
rect 10232 23817 10241 23851
rect 10241 23817 10275 23851
rect 10275 23817 10284 23851
rect 10232 23808 10284 23817
rect 10508 23808 10560 23860
rect 14464 23808 14516 23860
rect 14648 23851 14700 23860
rect 14648 23817 14657 23851
rect 14657 23817 14691 23851
rect 14691 23817 14700 23851
rect 14648 23808 14700 23817
rect 18328 23808 18380 23860
rect 19156 23808 19208 23860
rect 19616 23808 19668 23860
rect 20812 23808 20864 23860
rect 21824 23851 21876 23860
rect 21824 23817 21833 23851
rect 21833 23817 21867 23851
rect 21867 23817 21876 23851
rect 21824 23808 21876 23817
rect 23204 23808 23256 23860
rect 25228 23808 25280 23860
rect 8116 23740 8168 23792
rect 9312 23740 9364 23792
rect 6184 23672 6236 23724
rect 6460 23672 6512 23724
rect 6828 23715 6880 23724
rect 6828 23681 6837 23715
rect 6837 23681 6871 23715
rect 6871 23681 6880 23715
rect 6828 23672 6880 23681
rect 6276 23604 6328 23656
rect 4344 23536 4396 23588
rect 3976 23468 4028 23520
rect 8852 23672 8904 23724
rect 9496 23672 9548 23724
rect 9864 23715 9916 23724
rect 9864 23681 9873 23715
rect 9873 23681 9907 23715
rect 9907 23681 9916 23715
rect 9864 23672 9916 23681
rect 15844 23740 15896 23792
rect 13544 23672 13596 23724
rect 14372 23672 14424 23724
rect 12716 23604 12768 23656
rect 17224 23672 17276 23724
rect 21732 23740 21784 23792
rect 22008 23740 22060 23792
rect 22100 23740 22152 23792
rect 22560 23740 22612 23792
rect 13452 23536 13504 23588
rect 14188 23536 14240 23588
rect 15752 23579 15804 23588
rect 15752 23545 15761 23579
rect 15761 23545 15795 23579
rect 15795 23545 15804 23579
rect 15752 23536 15804 23545
rect 8852 23468 8904 23520
rect 10784 23511 10836 23520
rect 10784 23477 10793 23511
rect 10793 23477 10827 23511
rect 10827 23477 10836 23511
rect 10784 23468 10836 23477
rect 14832 23511 14884 23520
rect 14832 23477 14841 23511
rect 14841 23477 14875 23511
rect 14875 23477 14884 23511
rect 14832 23468 14884 23477
rect 16764 23468 16816 23520
rect 17040 23536 17092 23588
rect 19432 23672 19484 23724
rect 22928 23672 22980 23724
rect 19800 23604 19852 23656
rect 23940 23647 23992 23656
rect 20720 23536 20772 23588
rect 23940 23613 23949 23647
rect 23949 23613 23983 23647
rect 23983 23613 23992 23647
rect 23940 23604 23992 23613
rect 25320 23672 25372 23724
rect 26148 23672 26200 23724
rect 28264 23672 28316 23724
rect 24860 23604 24912 23656
rect 25504 23604 25556 23656
rect 17500 23468 17552 23520
rect 19340 23468 19392 23520
rect 19892 23468 19944 23520
rect 21180 23468 21232 23520
rect 26884 23536 26936 23588
rect 22928 23468 22980 23520
rect 25136 23511 25188 23520
rect 25136 23477 25145 23511
rect 25145 23477 25179 23511
rect 25179 23477 25188 23511
rect 25136 23468 25188 23477
rect 27528 23468 27580 23520
rect 28632 23511 28684 23520
rect 28632 23477 28641 23511
rect 28641 23477 28675 23511
rect 28675 23477 28684 23511
rect 28632 23468 28684 23477
rect 4492 23366 4544 23418
rect 4556 23366 4608 23418
rect 4620 23366 4672 23418
rect 4684 23366 4736 23418
rect 4748 23366 4800 23418
rect 11576 23366 11628 23418
rect 11640 23366 11692 23418
rect 11704 23366 11756 23418
rect 11768 23366 11820 23418
rect 11832 23366 11884 23418
rect 18660 23366 18712 23418
rect 18724 23366 18776 23418
rect 18788 23366 18840 23418
rect 18852 23366 18904 23418
rect 18916 23366 18968 23418
rect 25744 23366 25796 23418
rect 25808 23366 25860 23418
rect 25872 23366 25924 23418
rect 25936 23366 25988 23418
rect 26000 23366 26052 23418
rect 4344 23307 4396 23316
rect 4344 23273 4353 23307
rect 4353 23273 4387 23307
rect 4387 23273 4396 23307
rect 4344 23264 4396 23273
rect 6184 23307 6236 23316
rect 6184 23273 6193 23307
rect 6193 23273 6227 23307
rect 6227 23273 6236 23307
rect 6184 23264 6236 23273
rect 10968 23264 11020 23316
rect 14188 23307 14240 23316
rect 7748 23128 7800 23180
rect 4160 23060 4212 23112
rect 4344 23103 4396 23112
rect 4344 23069 4353 23103
rect 4353 23069 4387 23103
rect 4387 23069 4396 23103
rect 4344 23060 4396 23069
rect 4988 23060 5040 23112
rect 6552 23060 6604 23112
rect 7380 23060 7432 23112
rect 8116 23103 8168 23112
rect 8116 23069 8125 23103
rect 8125 23069 8159 23103
rect 8159 23069 8168 23103
rect 8116 23060 8168 23069
rect 9588 23060 9640 23112
rect 10324 23060 10376 23112
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 14188 23273 14197 23307
rect 14197 23273 14231 23307
rect 14231 23273 14240 23307
rect 14188 23264 14240 23273
rect 14372 23264 14424 23316
rect 15844 23307 15896 23316
rect 13176 23239 13228 23248
rect 13176 23205 13185 23239
rect 13185 23205 13219 23239
rect 13219 23205 13228 23239
rect 15844 23273 15853 23307
rect 15853 23273 15887 23307
rect 15887 23273 15896 23307
rect 15844 23264 15896 23273
rect 17040 23307 17092 23316
rect 17040 23273 17049 23307
rect 17049 23273 17083 23307
rect 17083 23273 17092 23307
rect 17040 23264 17092 23273
rect 19156 23264 19208 23316
rect 13176 23196 13228 23205
rect 13268 23128 13320 23180
rect 19340 23196 19392 23248
rect 15108 23128 15160 23180
rect 16948 23128 17000 23180
rect 12532 23103 12584 23112
rect 6276 23035 6328 23044
rect 6276 23001 6285 23035
rect 6285 23001 6319 23035
rect 6319 23001 6328 23035
rect 6276 22992 6328 23001
rect 6460 23035 6512 23044
rect 6460 23001 6469 23035
rect 6469 23001 6503 23035
rect 6503 23001 6512 23035
rect 6460 22992 6512 23001
rect 10048 23035 10100 23044
rect 1584 22924 1636 22976
rect 3792 22924 3844 22976
rect 7012 22967 7064 22976
rect 7012 22933 7021 22967
rect 7021 22933 7055 22967
rect 7055 22933 7064 22967
rect 7012 22924 7064 22933
rect 7472 22967 7524 22976
rect 7472 22933 7481 22967
rect 7481 22933 7515 22967
rect 7515 22933 7524 22967
rect 7472 22924 7524 22933
rect 10048 23001 10057 23035
rect 10057 23001 10091 23035
rect 10091 23001 10100 23035
rect 10048 22992 10100 23001
rect 10784 22992 10836 23044
rect 12532 23069 12541 23103
rect 12541 23069 12575 23103
rect 12575 23069 12584 23103
rect 12532 23060 12584 23069
rect 13544 23060 13596 23112
rect 14372 23103 14424 23112
rect 14372 23069 14381 23103
rect 14381 23069 14415 23103
rect 14415 23069 14424 23103
rect 14372 23060 14424 23069
rect 15016 23060 15068 23112
rect 15384 23103 15436 23112
rect 15384 23069 15391 23103
rect 15391 23069 15436 23103
rect 15384 23060 15436 23069
rect 16304 23060 16356 23112
rect 16488 23103 16540 23112
rect 16488 23069 16497 23103
rect 16497 23069 16531 23103
rect 16531 23069 16540 23103
rect 16488 23060 16540 23069
rect 18972 23060 19024 23112
rect 19432 23060 19484 23112
rect 19597 23103 19649 23112
rect 19597 23069 19622 23103
rect 19622 23069 19649 23103
rect 19597 23060 19649 23069
rect 19892 23264 19944 23316
rect 20812 23264 20864 23316
rect 22744 23307 22796 23316
rect 22744 23273 22753 23307
rect 22753 23273 22787 23307
rect 22787 23273 22796 23307
rect 22744 23264 22796 23273
rect 21088 23128 21140 23180
rect 25228 23128 25280 23180
rect 26240 23128 26292 23180
rect 26976 23128 27028 23180
rect 27804 23171 27856 23180
rect 27804 23137 27813 23171
rect 27813 23137 27847 23171
rect 27847 23137 27856 23171
rect 27804 23128 27856 23137
rect 28080 23171 28132 23180
rect 28080 23137 28089 23171
rect 28089 23137 28123 23171
rect 28123 23137 28132 23171
rect 28080 23128 28132 23137
rect 28448 23128 28500 23180
rect 19984 23060 20036 23112
rect 20904 23103 20956 23112
rect 20904 23069 20913 23103
rect 20913 23069 20947 23103
rect 20947 23069 20956 23103
rect 20904 23060 20956 23069
rect 21180 23103 21232 23112
rect 21180 23069 21189 23103
rect 21189 23069 21223 23103
rect 21223 23069 21232 23103
rect 21180 23060 21232 23069
rect 21824 23060 21876 23112
rect 14096 22992 14148 23044
rect 10416 22924 10468 22976
rect 16672 22992 16724 23044
rect 21272 22992 21324 23044
rect 24216 23060 24268 23112
rect 24768 23103 24820 23112
rect 24768 23069 24777 23103
rect 24777 23069 24811 23103
rect 24811 23069 24820 23103
rect 24768 23060 24820 23069
rect 25320 23060 25372 23112
rect 27712 23103 27764 23112
rect 27712 23069 27730 23103
rect 27730 23069 27764 23103
rect 27712 23060 27764 23069
rect 28540 23103 28592 23112
rect 28540 23069 28549 23103
rect 28549 23069 28583 23103
rect 28583 23069 28592 23103
rect 28540 23060 28592 23069
rect 15660 22924 15712 22976
rect 19340 22924 19392 22976
rect 19708 22924 19760 22976
rect 21088 22967 21140 22976
rect 21088 22933 21097 22967
rect 21097 22933 21131 22967
rect 21131 22933 21140 22967
rect 21088 22924 21140 22933
rect 22008 22924 22060 22976
rect 25964 22967 26016 22976
rect 25964 22933 25973 22967
rect 25973 22933 26007 22967
rect 26007 22933 26016 22967
rect 25964 22924 26016 22933
rect 8034 22822 8086 22874
rect 8098 22822 8150 22874
rect 8162 22822 8214 22874
rect 8226 22822 8278 22874
rect 8290 22822 8342 22874
rect 15118 22822 15170 22874
rect 15182 22822 15234 22874
rect 15246 22822 15298 22874
rect 15310 22822 15362 22874
rect 15374 22822 15426 22874
rect 22202 22822 22254 22874
rect 22266 22822 22318 22874
rect 22330 22822 22382 22874
rect 22394 22822 22446 22874
rect 22458 22822 22510 22874
rect 29286 22822 29338 22874
rect 29350 22822 29402 22874
rect 29414 22822 29466 22874
rect 29478 22822 29530 22874
rect 29542 22822 29594 22874
rect 4988 22720 5040 22772
rect 6552 22720 6604 22772
rect 9680 22763 9732 22772
rect 9680 22729 9689 22763
rect 9689 22729 9723 22763
rect 9723 22729 9732 22763
rect 9680 22720 9732 22729
rect 10324 22720 10376 22772
rect 10416 22720 10468 22772
rect 12992 22763 13044 22772
rect 12992 22729 13001 22763
rect 13001 22729 13035 22763
rect 13035 22729 13044 22763
rect 12992 22720 13044 22729
rect 14832 22720 14884 22772
rect 16672 22763 16724 22772
rect 16672 22729 16681 22763
rect 16681 22729 16715 22763
rect 16715 22729 16724 22763
rect 16672 22720 16724 22729
rect 18144 22720 18196 22772
rect 18328 22720 18380 22772
rect 19340 22763 19392 22772
rect 19340 22729 19349 22763
rect 19349 22729 19383 22763
rect 19383 22729 19392 22763
rect 19340 22720 19392 22729
rect 20812 22720 20864 22772
rect 24768 22720 24820 22772
rect 25964 22720 26016 22772
rect 3332 22695 3384 22704
rect 3332 22661 3341 22695
rect 3341 22661 3375 22695
rect 3375 22661 3384 22695
rect 3332 22652 3384 22661
rect 6460 22652 6512 22704
rect 8852 22695 8904 22704
rect 8852 22661 8861 22695
rect 8861 22661 8895 22695
rect 8895 22661 8904 22695
rect 8852 22652 8904 22661
rect 10048 22652 10100 22704
rect 11980 22695 12032 22704
rect 11980 22661 11989 22695
rect 11989 22661 12023 22695
rect 12023 22661 12032 22695
rect 11980 22652 12032 22661
rect 1584 22627 1636 22636
rect 1584 22593 1593 22627
rect 1593 22593 1627 22627
rect 1627 22593 1636 22627
rect 1584 22584 1636 22593
rect 2228 22584 2280 22636
rect 3056 22584 3108 22636
rect 3976 22627 4028 22636
rect 3976 22593 3985 22627
rect 3985 22593 4019 22627
rect 4019 22593 4028 22627
rect 3976 22584 4028 22593
rect 4252 22627 4304 22636
rect 4252 22593 4261 22627
rect 4261 22593 4295 22627
rect 4295 22593 4304 22627
rect 4252 22584 4304 22593
rect 1768 22491 1820 22500
rect 1768 22457 1777 22491
rect 1777 22457 1811 22491
rect 1811 22457 1820 22491
rect 1768 22448 1820 22457
rect 7288 22584 7340 22636
rect 7564 22627 7616 22636
rect 7564 22593 7573 22627
rect 7573 22593 7607 22627
rect 7607 22593 7616 22627
rect 7564 22584 7616 22593
rect 13544 22652 13596 22704
rect 15752 22652 15804 22704
rect 21088 22652 21140 22704
rect 15016 22627 15068 22636
rect 15016 22593 15025 22627
rect 15025 22593 15059 22627
rect 15059 22593 15068 22627
rect 15016 22584 15068 22593
rect 16856 22627 16908 22636
rect 8852 22448 8904 22500
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 16948 22627 17000 22636
rect 16948 22593 16957 22627
rect 16957 22593 16991 22627
rect 16991 22593 17000 22627
rect 16948 22584 17000 22593
rect 19248 22584 19300 22636
rect 21548 22584 21600 22636
rect 21824 22627 21876 22636
rect 21824 22593 21833 22627
rect 21833 22593 21867 22627
rect 21867 22593 21876 22627
rect 21824 22584 21876 22593
rect 22560 22627 22612 22636
rect 22560 22593 22569 22627
rect 22569 22593 22603 22627
rect 22603 22593 22612 22627
rect 22560 22584 22612 22593
rect 23112 22652 23164 22704
rect 24216 22652 24268 22704
rect 22836 22627 22888 22636
rect 22836 22593 22845 22627
rect 22845 22593 22879 22627
rect 22879 22593 22888 22627
rect 22836 22584 22888 22593
rect 16396 22516 16448 22568
rect 17868 22448 17920 22500
rect 19616 22448 19668 22500
rect 21916 22448 21968 22500
rect 22744 22448 22796 22500
rect 25136 22584 25188 22636
rect 28080 22584 28132 22636
rect 25320 22516 25372 22568
rect 24032 22448 24084 22500
rect 3516 22380 3568 22432
rect 8208 22423 8260 22432
rect 8208 22389 8217 22423
rect 8217 22389 8251 22423
rect 8251 22389 8260 22423
rect 8208 22380 8260 22389
rect 9956 22380 10008 22432
rect 19892 22380 19944 22432
rect 23388 22380 23440 22432
rect 25596 22423 25648 22432
rect 25596 22389 25605 22423
rect 25605 22389 25639 22423
rect 25639 22389 25648 22423
rect 25596 22380 25648 22389
rect 27896 22380 27948 22432
rect 4492 22278 4544 22330
rect 4556 22278 4608 22330
rect 4620 22278 4672 22330
rect 4684 22278 4736 22330
rect 4748 22278 4800 22330
rect 11576 22278 11628 22330
rect 11640 22278 11692 22330
rect 11704 22278 11756 22330
rect 11768 22278 11820 22330
rect 11832 22278 11884 22330
rect 18660 22278 18712 22330
rect 18724 22278 18776 22330
rect 18788 22278 18840 22330
rect 18852 22278 18904 22330
rect 18916 22278 18968 22330
rect 25744 22278 25796 22330
rect 25808 22278 25860 22330
rect 25872 22278 25924 22330
rect 25936 22278 25988 22330
rect 26000 22278 26052 22330
rect 2228 22219 2280 22228
rect 2228 22185 2237 22219
rect 2237 22185 2271 22219
rect 2271 22185 2280 22219
rect 2228 22176 2280 22185
rect 7564 22108 7616 22160
rect 2964 22040 3016 22092
rect 7012 22040 7064 22092
rect 1676 21972 1728 22024
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 6552 21972 6604 22024
rect 11980 22176 12032 22228
rect 13176 22040 13228 22092
rect 14924 22083 14976 22092
rect 7840 21972 7892 22024
rect 9864 21972 9916 22024
rect 14188 21972 14240 22024
rect 7380 21904 7432 21956
rect 8208 21904 8260 21956
rect 8668 21904 8720 21956
rect 9404 21904 9456 21956
rect 10600 21947 10652 21956
rect 10600 21913 10609 21947
rect 10609 21913 10643 21947
rect 10643 21913 10652 21947
rect 10600 21904 10652 21913
rect 14464 22015 14516 22024
rect 14464 21981 14473 22015
rect 14473 21981 14507 22015
rect 14507 21981 14516 22015
rect 14924 22049 14933 22083
rect 14933 22049 14967 22083
rect 14967 22049 14976 22083
rect 14924 22040 14976 22049
rect 14464 21972 14516 21981
rect 14740 22015 14792 22024
rect 14740 21981 14749 22015
rect 14749 21981 14783 22015
rect 14783 21981 14792 22015
rect 19064 22176 19116 22228
rect 22008 22176 22060 22228
rect 14740 21972 14792 21981
rect 18328 22015 18380 22024
rect 18328 21981 18337 22015
rect 18337 21981 18371 22015
rect 18371 21981 18380 22015
rect 18328 21972 18380 21981
rect 19248 22040 19300 22092
rect 19892 22083 19944 22092
rect 19892 22049 19901 22083
rect 19901 22049 19935 22083
rect 19935 22049 19944 22083
rect 19892 22040 19944 22049
rect 21364 22083 21416 22092
rect 21364 22049 21382 22083
rect 21382 22049 21416 22083
rect 21364 22040 21416 22049
rect 21640 22040 21692 22092
rect 21824 22108 21876 22160
rect 22008 22040 22060 22092
rect 18972 21972 19024 22024
rect 19616 22015 19668 22024
rect 19616 21981 19625 22015
rect 19625 21981 19659 22015
rect 19659 21981 19668 22015
rect 19616 21972 19668 21981
rect 21180 22015 21232 22024
rect 21180 21981 21189 22015
rect 21189 21981 21223 22015
rect 21223 21981 21232 22015
rect 26792 22040 26844 22092
rect 28080 22083 28132 22092
rect 28080 22049 28089 22083
rect 28089 22049 28123 22083
rect 28123 22049 28132 22083
rect 28080 22040 28132 22049
rect 21180 21972 21232 21981
rect 14556 21904 14608 21956
rect 16856 21904 16908 21956
rect 19156 21904 19208 21956
rect 19708 21947 19760 21956
rect 19708 21913 19717 21947
rect 19717 21913 19751 21947
rect 19751 21913 19760 21947
rect 19708 21904 19760 21913
rect 25596 21972 25648 22024
rect 22744 21904 22796 21956
rect 3884 21879 3936 21888
rect 3884 21845 3893 21879
rect 3893 21845 3927 21879
rect 3927 21845 3936 21879
rect 3884 21836 3936 21845
rect 9772 21879 9824 21888
rect 9772 21845 9781 21879
rect 9781 21845 9815 21879
rect 9815 21845 9824 21879
rect 10140 21879 10192 21888
rect 9772 21836 9824 21845
rect 10140 21845 10149 21879
rect 10149 21845 10183 21879
rect 10183 21845 10192 21879
rect 10140 21836 10192 21845
rect 13360 21836 13412 21888
rect 17500 21879 17552 21888
rect 17500 21845 17509 21879
rect 17509 21845 17543 21879
rect 17543 21845 17552 21879
rect 17500 21836 17552 21845
rect 17960 21879 18012 21888
rect 17960 21845 17969 21879
rect 17969 21845 18003 21879
rect 18003 21845 18012 21879
rect 17960 21836 18012 21845
rect 20904 21836 20956 21888
rect 24768 21904 24820 21956
rect 28448 21904 28500 21956
rect 24124 21836 24176 21888
rect 24584 21836 24636 21888
rect 26976 21836 27028 21888
rect 27252 21836 27304 21888
rect 27988 21879 28040 21888
rect 27988 21845 27997 21879
rect 27997 21845 28031 21879
rect 28031 21845 28040 21879
rect 27988 21836 28040 21845
rect 8034 21734 8086 21786
rect 8098 21734 8150 21786
rect 8162 21734 8214 21786
rect 8226 21734 8278 21786
rect 8290 21734 8342 21786
rect 15118 21734 15170 21786
rect 15182 21734 15234 21786
rect 15246 21734 15298 21786
rect 15310 21734 15362 21786
rect 15374 21734 15426 21786
rect 22202 21734 22254 21786
rect 22266 21734 22318 21786
rect 22330 21734 22382 21786
rect 22394 21734 22446 21786
rect 22458 21734 22510 21786
rect 29286 21734 29338 21786
rect 29350 21734 29402 21786
rect 29414 21734 29466 21786
rect 29478 21734 29530 21786
rect 29542 21734 29594 21786
rect 4344 21632 4396 21684
rect 8668 21675 8720 21684
rect 8668 21641 8677 21675
rect 8677 21641 8711 21675
rect 8711 21641 8720 21675
rect 8668 21632 8720 21641
rect 8944 21632 8996 21684
rect 9680 21632 9732 21684
rect 10508 21632 10560 21684
rect 12900 21632 12952 21684
rect 13912 21632 13964 21684
rect 14096 21675 14148 21684
rect 14096 21641 14105 21675
rect 14105 21641 14139 21675
rect 14139 21641 14148 21675
rect 14096 21632 14148 21641
rect 14280 21632 14332 21684
rect 14372 21632 14424 21684
rect 16948 21632 17000 21684
rect 4160 21496 4212 21548
rect 4344 21496 4396 21548
rect 10048 21564 10100 21616
rect 15384 21564 15436 21616
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 2964 21292 3016 21344
rect 3700 21335 3752 21344
rect 3700 21301 3709 21335
rect 3709 21301 3743 21335
rect 3743 21301 3752 21335
rect 3700 21292 3752 21301
rect 8668 21292 8720 21344
rect 9680 21539 9732 21548
rect 9680 21505 9725 21539
rect 9725 21505 9732 21539
rect 9680 21496 9732 21505
rect 12440 21496 12492 21548
rect 12900 21496 12952 21548
rect 9588 21360 9640 21412
rect 9772 21360 9824 21412
rect 12716 21428 12768 21480
rect 13176 21428 13228 21480
rect 13360 21496 13412 21548
rect 14004 21496 14056 21548
rect 13544 21428 13596 21480
rect 14372 21539 14424 21548
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 14924 21496 14976 21548
rect 17960 21564 18012 21616
rect 18696 21564 18748 21616
rect 19708 21632 19760 21684
rect 21364 21632 21416 21684
rect 24032 21632 24084 21684
rect 27988 21632 28040 21684
rect 28540 21675 28592 21684
rect 28540 21641 28549 21675
rect 28549 21641 28583 21675
rect 28583 21641 28592 21675
rect 28540 21632 28592 21641
rect 17040 21539 17092 21548
rect 17040 21505 17049 21539
rect 17049 21505 17083 21539
rect 17083 21505 17092 21539
rect 17040 21496 17092 21505
rect 16580 21428 16632 21480
rect 17132 21471 17184 21480
rect 17132 21437 17141 21471
rect 17141 21437 17175 21471
rect 17175 21437 17184 21471
rect 17132 21428 17184 21437
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 17776 21428 17828 21480
rect 20812 21539 20864 21548
rect 20812 21505 20821 21539
rect 20821 21505 20855 21539
rect 20855 21505 20864 21539
rect 20812 21496 20864 21505
rect 20904 21496 20956 21548
rect 21732 21496 21784 21548
rect 23112 21564 23164 21616
rect 27620 21564 27672 21616
rect 24032 21539 24084 21548
rect 10876 21292 10928 21344
rect 14372 21292 14424 21344
rect 16488 21360 16540 21412
rect 18696 21360 18748 21412
rect 19340 21360 19392 21412
rect 21640 21428 21692 21480
rect 23112 21428 23164 21480
rect 24032 21505 24041 21539
rect 24041 21505 24075 21539
rect 24075 21505 24084 21539
rect 24032 21496 24084 21505
rect 24124 21539 24176 21548
rect 24124 21505 24133 21539
rect 24133 21505 24167 21539
rect 24167 21505 24176 21539
rect 24124 21496 24176 21505
rect 24768 21496 24820 21548
rect 28724 21539 28776 21548
rect 28724 21505 28733 21539
rect 28733 21505 28767 21539
rect 28767 21505 28776 21539
rect 28724 21496 28776 21505
rect 23664 21428 23716 21480
rect 26424 21428 26476 21480
rect 26884 21428 26936 21480
rect 27528 21471 27580 21480
rect 27528 21437 27537 21471
rect 27537 21437 27571 21471
rect 27571 21437 27580 21471
rect 27528 21428 27580 21437
rect 19892 21360 19944 21412
rect 22560 21360 22612 21412
rect 24032 21360 24084 21412
rect 26516 21360 26568 21412
rect 17408 21292 17460 21344
rect 20904 21335 20956 21344
rect 20904 21301 20913 21335
rect 20913 21301 20947 21335
rect 20947 21301 20956 21335
rect 20904 21292 20956 21301
rect 21364 21292 21416 21344
rect 23572 21292 23624 21344
rect 26240 21292 26292 21344
rect 4492 21190 4544 21242
rect 4556 21190 4608 21242
rect 4620 21190 4672 21242
rect 4684 21190 4736 21242
rect 4748 21190 4800 21242
rect 11576 21190 11628 21242
rect 11640 21190 11692 21242
rect 11704 21190 11756 21242
rect 11768 21190 11820 21242
rect 11832 21190 11884 21242
rect 18660 21190 18712 21242
rect 18724 21190 18776 21242
rect 18788 21190 18840 21242
rect 18852 21190 18904 21242
rect 18916 21190 18968 21242
rect 25744 21190 25796 21242
rect 25808 21190 25860 21242
rect 25872 21190 25924 21242
rect 25936 21190 25988 21242
rect 26000 21190 26052 21242
rect 9680 21088 9732 21140
rect 10600 21088 10652 21140
rect 12440 21131 12492 21140
rect 12440 21097 12449 21131
rect 12449 21097 12483 21131
rect 12483 21097 12492 21131
rect 13544 21131 13596 21140
rect 12440 21088 12492 21097
rect 13544 21097 13553 21131
rect 13553 21097 13587 21131
rect 13587 21097 13596 21131
rect 13544 21088 13596 21097
rect 16580 21131 16632 21140
rect 16580 21097 16589 21131
rect 16589 21097 16623 21131
rect 16623 21097 16632 21131
rect 16580 21088 16632 21097
rect 17132 21088 17184 21140
rect 17316 21088 17368 21140
rect 18328 21088 18380 21140
rect 19340 21088 19392 21140
rect 26056 21088 26108 21140
rect 26240 21131 26292 21140
rect 26240 21097 26249 21131
rect 26249 21097 26283 21131
rect 26283 21097 26292 21131
rect 26240 21088 26292 21097
rect 27712 21088 27764 21140
rect 28172 21088 28224 21140
rect 9496 21020 9548 21072
rect 9496 20927 9548 20936
rect 9496 20893 9505 20927
rect 9505 20893 9539 20927
rect 9539 20893 9548 20927
rect 9496 20884 9548 20893
rect 10784 21020 10836 21072
rect 16948 21020 17000 21072
rect 6552 20791 6604 20800
rect 6552 20757 6561 20791
rect 6561 20757 6595 20791
rect 6595 20757 6604 20791
rect 6552 20748 6604 20757
rect 7932 20748 7984 20800
rect 10140 20884 10192 20936
rect 10508 20884 10560 20936
rect 11980 20884 12032 20936
rect 12624 20927 12676 20936
rect 10876 20859 10928 20868
rect 10876 20825 10885 20859
rect 10885 20825 10919 20859
rect 10919 20825 10928 20859
rect 10876 20816 10928 20825
rect 12624 20893 12633 20927
rect 12633 20893 12667 20927
rect 12667 20893 12676 20927
rect 12624 20884 12676 20893
rect 14096 20884 14148 20936
rect 14648 20927 14700 20936
rect 14648 20893 14656 20927
rect 14656 20893 14690 20927
rect 14690 20893 14700 20927
rect 14648 20884 14700 20893
rect 10600 20791 10652 20800
rect 10600 20757 10609 20791
rect 10609 20757 10643 20791
rect 10643 20757 10652 20791
rect 10600 20748 10652 20757
rect 14188 20816 14240 20868
rect 14372 20859 14424 20868
rect 14372 20825 14381 20859
rect 14381 20825 14415 20859
rect 14415 20825 14424 20859
rect 14372 20816 14424 20825
rect 14280 20748 14332 20800
rect 14556 20816 14608 20868
rect 16396 20927 16448 20936
rect 16396 20893 16405 20927
rect 16405 20893 16439 20927
rect 16439 20893 16448 20927
rect 16396 20884 16448 20893
rect 16856 20884 16908 20936
rect 17408 20884 17460 20936
rect 20812 20952 20864 21004
rect 26976 21020 27028 21072
rect 21088 20952 21140 21004
rect 24584 20952 24636 21004
rect 26424 20952 26476 21004
rect 26700 20952 26752 21004
rect 27712 20995 27764 21004
rect 27712 20961 27721 20995
rect 27721 20961 27755 20995
rect 27755 20961 27764 20995
rect 27712 20952 27764 20961
rect 28080 20952 28132 21004
rect 21640 20927 21692 20936
rect 21640 20893 21649 20927
rect 21649 20893 21683 20927
rect 21683 20893 21692 20927
rect 21640 20884 21692 20893
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 23388 20884 23440 20893
rect 23664 20884 23716 20936
rect 26516 20884 26568 20936
rect 27620 20927 27672 20936
rect 27620 20893 27638 20927
rect 27638 20893 27672 20927
rect 27620 20884 27672 20893
rect 28264 20884 28316 20936
rect 21364 20816 21416 20868
rect 24492 20816 24544 20868
rect 18696 20791 18748 20800
rect 18696 20757 18705 20791
rect 18705 20757 18739 20791
rect 18739 20757 18748 20791
rect 18696 20748 18748 20757
rect 19248 20791 19300 20800
rect 19248 20757 19257 20791
rect 19257 20757 19291 20791
rect 19291 20757 19300 20791
rect 19248 20748 19300 20757
rect 23480 20791 23532 20800
rect 23480 20757 23489 20791
rect 23489 20757 23523 20791
rect 23523 20757 23532 20791
rect 23480 20748 23532 20757
rect 23848 20748 23900 20800
rect 24768 20748 24820 20800
rect 26148 20748 26200 20800
rect 27528 20748 27580 20800
rect 27804 20748 27856 20800
rect 8034 20646 8086 20698
rect 8098 20646 8150 20698
rect 8162 20646 8214 20698
rect 8226 20646 8278 20698
rect 8290 20646 8342 20698
rect 15118 20646 15170 20698
rect 15182 20646 15234 20698
rect 15246 20646 15298 20698
rect 15310 20646 15362 20698
rect 15374 20646 15426 20698
rect 22202 20646 22254 20698
rect 22266 20646 22318 20698
rect 22330 20646 22382 20698
rect 22394 20646 22446 20698
rect 22458 20646 22510 20698
rect 29286 20646 29338 20698
rect 29350 20646 29402 20698
rect 29414 20646 29466 20698
rect 29478 20646 29530 20698
rect 29542 20646 29594 20698
rect 1860 20544 1912 20596
rect 8300 20544 8352 20596
rect 3148 20451 3200 20460
rect 3148 20417 3157 20451
rect 3157 20417 3191 20451
rect 3191 20417 3200 20451
rect 3148 20408 3200 20417
rect 3240 20408 3292 20460
rect 4344 20476 4396 20528
rect 9772 20544 9824 20596
rect 11980 20587 12032 20596
rect 11980 20553 11989 20587
rect 11989 20553 12023 20587
rect 12023 20553 12032 20587
rect 11980 20544 12032 20553
rect 12624 20587 12676 20596
rect 12624 20553 12633 20587
rect 12633 20553 12667 20587
rect 12667 20553 12676 20587
rect 12624 20544 12676 20553
rect 4252 20408 4304 20460
rect 5908 20408 5960 20460
rect 7104 20451 7156 20460
rect 7104 20417 7113 20451
rect 7113 20417 7147 20451
rect 7147 20417 7156 20451
rect 7104 20408 7156 20417
rect 7472 20408 7524 20460
rect 8300 20408 8352 20460
rect 9128 20408 9180 20460
rect 3884 20340 3936 20392
rect 7012 20340 7064 20392
rect 7288 20340 7340 20392
rect 7380 20340 7432 20392
rect 7932 20340 7984 20392
rect 10508 20408 10560 20460
rect 12808 20451 12860 20460
rect 12808 20417 12817 20451
rect 12817 20417 12851 20451
rect 12851 20417 12860 20451
rect 12808 20408 12860 20417
rect 13268 20408 13320 20460
rect 14280 20544 14332 20596
rect 16396 20544 16448 20596
rect 16580 20544 16632 20596
rect 17316 20544 17368 20596
rect 17684 20544 17736 20596
rect 25044 20587 25096 20596
rect 25044 20553 25053 20587
rect 25053 20553 25087 20587
rect 25087 20553 25096 20587
rect 25044 20544 25096 20553
rect 14096 20519 14148 20528
rect 14096 20485 14105 20519
rect 14105 20485 14139 20519
rect 14139 20485 14148 20519
rect 14096 20476 14148 20485
rect 14188 20451 14240 20460
rect 14188 20417 14197 20451
rect 14197 20417 14231 20451
rect 14231 20417 14240 20451
rect 14188 20408 14240 20417
rect 20904 20476 20956 20528
rect 23480 20476 23532 20528
rect 25596 20476 25648 20528
rect 26976 20519 27028 20528
rect 26976 20485 26985 20519
rect 26985 20485 27019 20519
rect 27019 20485 27028 20519
rect 26976 20476 27028 20485
rect 27620 20476 27672 20528
rect 18696 20408 18748 20460
rect 19064 20408 19116 20460
rect 19892 20408 19944 20460
rect 21640 20408 21692 20460
rect 23848 20408 23900 20460
rect 24492 20451 24544 20460
rect 24492 20417 24501 20451
rect 24501 20417 24535 20451
rect 24535 20417 24544 20451
rect 24492 20408 24544 20417
rect 26148 20408 26200 20460
rect 20812 20340 20864 20392
rect 24768 20340 24820 20392
rect 26240 20340 26292 20392
rect 1676 20272 1728 20324
rect 4160 20272 4212 20324
rect 3976 20204 4028 20256
rect 6460 20247 6512 20256
rect 6460 20213 6469 20247
rect 6469 20213 6503 20247
rect 6503 20213 6512 20247
rect 6460 20204 6512 20213
rect 6920 20247 6972 20256
rect 6920 20213 6929 20247
rect 6929 20213 6963 20247
rect 6963 20213 6972 20247
rect 6920 20204 6972 20213
rect 7932 20204 7984 20256
rect 8116 20204 8168 20256
rect 9956 20204 10008 20256
rect 21640 20272 21692 20324
rect 23112 20315 23164 20324
rect 23112 20281 23121 20315
rect 23121 20281 23155 20315
rect 23155 20281 23164 20315
rect 23112 20272 23164 20281
rect 28448 20272 28500 20324
rect 10784 20204 10836 20256
rect 13360 20204 13412 20256
rect 14556 20204 14608 20256
rect 17776 20204 17828 20256
rect 18052 20204 18104 20256
rect 19248 20204 19300 20256
rect 19892 20204 19944 20256
rect 20628 20204 20680 20256
rect 25504 20204 25556 20256
rect 27988 20204 28040 20256
rect 28172 20204 28224 20256
rect 4492 20102 4544 20154
rect 4556 20102 4608 20154
rect 4620 20102 4672 20154
rect 4684 20102 4736 20154
rect 4748 20102 4800 20154
rect 11576 20102 11628 20154
rect 11640 20102 11692 20154
rect 11704 20102 11756 20154
rect 11768 20102 11820 20154
rect 11832 20102 11884 20154
rect 18660 20102 18712 20154
rect 18724 20102 18776 20154
rect 18788 20102 18840 20154
rect 18852 20102 18904 20154
rect 18916 20102 18968 20154
rect 25744 20102 25796 20154
rect 25808 20102 25860 20154
rect 25872 20102 25924 20154
rect 25936 20102 25988 20154
rect 26000 20102 26052 20154
rect 3240 20043 3292 20052
rect 3240 20009 3249 20043
rect 3249 20009 3283 20043
rect 3283 20009 3292 20043
rect 3240 20000 3292 20009
rect 5908 20043 5960 20052
rect 5908 20009 5917 20043
rect 5917 20009 5951 20043
rect 5951 20009 5960 20043
rect 5908 20000 5960 20009
rect 4160 19932 4212 19984
rect 6552 20000 6604 20052
rect 7012 20000 7064 20052
rect 8300 20043 8352 20052
rect 6460 19932 6512 19984
rect 7840 19932 7892 19984
rect 8300 20009 8309 20043
rect 8309 20009 8343 20043
rect 8343 20009 8352 20043
rect 8300 20000 8352 20009
rect 9956 20043 10008 20052
rect 9956 20009 9965 20043
rect 9965 20009 9999 20043
rect 9999 20009 10008 20043
rect 9956 20000 10008 20009
rect 12900 20000 12952 20052
rect 13544 20000 13596 20052
rect 9588 19932 9640 19984
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 2228 19796 2280 19848
rect 2688 19796 2740 19848
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 4252 19839 4304 19848
rect 4252 19805 4261 19839
rect 4261 19805 4295 19839
rect 4295 19805 4304 19839
rect 4252 19796 4304 19805
rect 4436 19839 4488 19848
rect 4436 19805 4445 19839
rect 4445 19805 4479 19839
rect 4479 19805 4488 19839
rect 4436 19796 4488 19805
rect 5264 19839 5316 19848
rect 3700 19728 3752 19780
rect 3884 19728 3936 19780
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 4068 19660 4120 19712
rect 5264 19805 5273 19839
rect 5273 19805 5307 19839
rect 5307 19805 5316 19839
rect 5264 19796 5316 19805
rect 7104 19839 7156 19848
rect 7104 19805 7113 19839
rect 7113 19805 7147 19839
rect 7147 19805 7156 19839
rect 7104 19796 7156 19805
rect 9864 19864 9916 19916
rect 14648 19932 14700 19984
rect 13544 19864 13596 19916
rect 13912 19864 13964 19916
rect 14464 19864 14516 19916
rect 7012 19728 7064 19780
rect 7380 19796 7432 19848
rect 10600 19796 10652 19848
rect 7472 19728 7524 19780
rect 9864 19728 9916 19780
rect 10784 19771 10836 19780
rect 10784 19737 10793 19771
rect 10793 19737 10827 19771
rect 10827 19737 10836 19771
rect 10784 19728 10836 19737
rect 11520 19771 11572 19780
rect 11520 19737 11529 19771
rect 11529 19737 11563 19771
rect 11563 19737 11572 19771
rect 11520 19728 11572 19737
rect 4712 19660 4764 19712
rect 5724 19660 5776 19712
rect 7288 19660 7340 19712
rect 10876 19660 10928 19712
rect 12716 19660 12768 19712
rect 14556 19839 14608 19848
rect 12900 19728 12952 19780
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 17684 19932 17736 19984
rect 22744 20000 22796 20052
rect 25596 20000 25648 20052
rect 26240 20000 26292 20052
rect 25504 19932 25556 19984
rect 27804 19932 27856 19984
rect 17776 19864 17828 19916
rect 18144 19864 18196 19916
rect 19248 19907 19300 19916
rect 19248 19873 19257 19907
rect 19257 19873 19291 19907
rect 19291 19873 19300 19907
rect 19248 19864 19300 19873
rect 20720 19864 20772 19916
rect 17316 19728 17368 19780
rect 18604 19839 18656 19848
rect 18604 19805 18613 19839
rect 18613 19805 18647 19839
rect 18647 19805 18656 19839
rect 18604 19796 18656 19805
rect 20628 19796 20680 19848
rect 20996 19839 21048 19848
rect 20996 19805 21005 19839
rect 21005 19805 21039 19839
rect 21039 19805 21048 19839
rect 20996 19796 21048 19805
rect 20536 19728 20588 19780
rect 21824 19796 21876 19848
rect 23020 19864 23072 19916
rect 22744 19839 22796 19848
rect 22744 19805 22753 19839
rect 22753 19805 22787 19839
rect 22787 19805 22796 19839
rect 22744 19796 22796 19805
rect 23112 19796 23164 19848
rect 27988 19839 28040 19848
rect 24768 19728 24820 19780
rect 27988 19805 27997 19839
rect 27997 19805 28031 19839
rect 28031 19805 28040 19839
rect 27988 19796 28040 19805
rect 13360 19660 13412 19712
rect 13820 19660 13872 19712
rect 15568 19703 15620 19712
rect 15568 19669 15577 19703
rect 15577 19669 15611 19703
rect 15611 19669 15620 19703
rect 15568 19660 15620 19669
rect 16672 19660 16724 19712
rect 18144 19703 18196 19712
rect 18144 19669 18153 19703
rect 18153 19669 18187 19703
rect 18187 19669 18196 19703
rect 18144 19660 18196 19669
rect 20352 19660 20404 19712
rect 22836 19660 22888 19712
rect 28172 19703 28224 19712
rect 28172 19669 28181 19703
rect 28181 19669 28215 19703
rect 28215 19669 28224 19703
rect 28172 19660 28224 19669
rect 8034 19558 8086 19610
rect 8098 19558 8150 19610
rect 8162 19558 8214 19610
rect 8226 19558 8278 19610
rect 8290 19558 8342 19610
rect 15118 19558 15170 19610
rect 15182 19558 15234 19610
rect 15246 19558 15298 19610
rect 15310 19558 15362 19610
rect 15374 19558 15426 19610
rect 22202 19558 22254 19610
rect 22266 19558 22318 19610
rect 22330 19558 22382 19610
rect 22394 19558 22446 19610
rect 22458 19558 22510 19610
rect 29286 19558 29338 19610
rect 29350 19558 29402 19610
rect 29414 19558 29466 19610
rect 29478 19558 29530 19610
rect 29542 19558 29594 19610
rect 2780 19499 2832 19508
rect 2780 19465 2789 19499
rect 2789 19465 2823 19499
rect 2823 19465 2832 19499
rect 2780 19456 2832 19465
rect 3148 19456 3200 19508
rect 4436 19456 4488 19508
rect 4712 19499 4764 19508
rect 4712 19465 4721 19499
rect 4721 19465 4755 19499
rect 4755 19465 4764 19499
rect 4712 19456 4764 19465
rect 5264 19499 5316 19508
rect 5264 19465 5273 19499
rect 5273 19465 5307 19499
rect 5307 19465 5316 19499
rect 5264 19456 5316 19465
rect 6920 19456 6972 19508
rect 10048 19499 10100 19508
rect 10048 19465 10057 19499
rect 10057 19465 10091 19499
rect 10091 19465 10100 19499
rect 10048 19456 10100 19465
rect 12072 19456 12124 19508
rect 2412 19431 2464 19440
rect 2412 19397 2421 19431
rect 2421 19397 2455 19431
rect 2455 19397 2464 19431
rect 2412 19388 2464 19397
rect 4252 19388 4304 19440
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 2320 19363 2372 19372
rect 2320 19329 2329 19363
rect 2329 19329 2363 19363
rect 2363 19329 2372 19363
rect 2320 19320 2372 19329
rect 2504 19320 2556 19372
rect 3884 19363 3936 19372
rect 3884 19329 3893 19363
rect 3893 19329 3927 19363
rect 3927 19329 3936 19363
rect 3884 19320 3936 19329
rect 4068 19320 4120 19372
rect 5908 19320 5960 19372
rect 7656 19388 7708 19440
rect 9128 19431 9180 19440
rect 9128 19397 9137 19431
rect 9137 19397 9171 19431
rect 9171 19397 9180 19431
rect 9128 19388 9180 19397
rect 9404 19388 9456 19440
rect 9496 19320 9548 19372
rect 9864 19320 9916 19372
rect 16120 19456 16172 19508
rect 17040 19456 17092 19508
rect 17316 19499 17368 19508
rect 17316 19465 17325 19499
rect 17325 19465 17359 19499
rect 17359 19465 17368 19499
rect 17316 19456 17368 19465
rect 20352 19499 20404 19508
rect 13820 19363 13872 19372
rect 13820 19329 13829 19363
rect 13829 19329 13863 19363
rect 13863 19329 13872 19363
rect 13820 19320 13872 19329
rect 18144 19388 18196 19440
rect 14648 19320 14700 19372
rect 16672 19363 16724 19372
rect 7104 19252 7156 19304
rect 7380 19252 7432 19304
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 16856 19363 16908 19372
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 20352 19465 20361 19499
rect 20361 19465 20395 19499
rect 20395 19465 20404 19499
rect 20352 19456 20404 19465
rect 27804 19499 27856 19508
rect 27804 19465 27813 19499
rect 27813 19465 27847 19499
rect 27847 19465 27856 19499
rect 27804 19456 27856 19465
rect 20444 19388 20496 19440
rect 23480 19431 23532 19440
rect 23480 19397 23489 19431
rect 23489 19397 23523 19431
rect 23523 19397 23532 19431
rect 23480 19388 23532 19397
rect 19984 19320 20036 19372
rect 23112 19320 23164 19372
rect 23204 19320 23256 19372
rect 24584 19363 24636 19372
rect 18052 19252 18104 19304
rect 1952 19184 2004 19236
rect 2320 19116 2372 19168
rect 2412 19116 2464 19168
rect 6184 19116 6236 19168
rect 7288 19116 7340 19168
rect 10232 19184 10284 19236
rect 7656 19116 7708 19168
rect 7932 19116 7984 19168
rect 8208 19159 8260 19168
rect 8208 19125 8217 19159
rect 8217 19125 8251 19159
rect 8251 19125 8260 19159
rect 8208 19116 8260 19125
rect 13912 19159 13964 19168
rect 13912 19125 13921 19159
rect 13921 19125 13955 19159
rect 13955 19125 13964 19159
rect 13912 19116 13964 19125
rect 16028 19116 16080 19168
rect 16304 19116 16356 19168
rect 16580 19116 16632 19168
rect 16764 19116 16816 19168
rect 20536 19252 20588 19304
rect 24584 19329 24593 19363
rect 24593 19329 24627 19363
rect 24627 19329 24636 19363
rect 24584 19320 24636 19329
rect 21364 19116 21416 19168
rect 24768 19295 24820 19304
rect 24768 19261 24777 19295
rect 24777 19261 24811 19295
rect 24811 19261 24820 19295
rect 24768 19252 24820 19261
rect 26332 19295 26384 19304
rect 26332 19261 26341 19295
rect 26341 19261 26375 19295
rect 26375 19261 26384 19295
rect 26332 19252 26384 19261
rect 27712 19252 27764 19304
rect 28172 19320 28224 19372
rect 28080 19295 28132 19304
rect 28080 19261 28089 19295
rect 28089 19261 28123 19295
rect 28123 19261 28132 19295
rect 28080 19252 28132 19261
rect 23112 19159 23164 19168
rect 23112 19125 23121 19159
rect 23121 19125 23155 19159
rect 23155 19125 23164 19159
rect 23112 19116 23164 19125
rect 27436 19159 27488 19168
rect 27436 19125 27445 19159
rect 27445 19125 27479 19159
rect 27479 19125 27488 19159
rect 27436 19116 27488 19125
rect 28172 19116 28224 19168
rect 28448 19116 28500 19168
rect 4492 19014 4544 19066
rect 4556 19014 4608 19066
rect 4620 19014 4672 19066
rect 4684 19014 4736 19066
rect 4748 19014 4800 19066
rect 11576 19014 11628 19066
rect 11640 19014 11692 19066
rect 11704 19014 11756 19066
rect 11768 19014 11820 19066
rect 11832 19014 11884 19066
rect 18660 19014 18712 19066
rect 18724 19014 18776 19066
rect 18788 19014 18840 19066
rect 18852 19014 18904 19066
rect 18916 19014 18968 19066
rect 25744 19014 25796 19066
rect 25808 19014 25860 19066
rect 25872 19014 25924 19066
rect 25936 19014 25988 19066
rect 26000 19014 26052 19066
rect 2228 18955 2280 18964
rect 2228 18921 2237 18955
rect 2237 18921 2271 18955
rect 2271 18921 2280 18955
rect 2228 18912 2280 18921
rect 5356 18912 5408 18964
rect 7472 18912 7524 18964
rect 2412 18776 2464 18828
rect 1492 18572 1544 18624
rect 2320 18751 2372 18760
rect 2320 18717 2329 18751
rect 2329 18717 2363 18751
rect 2363 18717 2372 18751
rect 2320 18708 2372 18717
rect 2504 18683 2556 18692
rect 2504 18649 2513 18683
rect 2513 18649 2547 18683
rect 2547 18649 2556 18683
rect 2504 18640 2556 18649
rect 2596 18640 2648 18692
rect 5540 18844 5592 18896
rect 7748 18844 7800 18896
rect 5632 18776 5684 18828
rect 8392 18912 8444 18964
rect 9496 18955 9548 18964
rect 9496 18921 9505 18955
rect 9505 18921 9539 18955
rect 9539 18921 9548 18955
rect 9496 18912 9548 18921
rect 9772 18912 9824 18964
rect 15476 18955 15528 18964
rect 15476 18921 15485 18955
rect 15485 18921 15519 18955
rect 15519 18921 15528 18955
rect 15476 18912 15528 18921
rect 17868 18955 17920 18964
rect 17868 18921 17877 18955
rect 17877 18921 17911 18955
rect 17911 18921 17920 18955
rect 17868 18912 17920 18921
rect 20720 18912 20772 18964
rect 21732 18912 21784 18964
rect 23664 18912 23716 18964
rect 24676 18912 24728 18964
rect 27988 18912 28040 18964
rect 16304 18844 16356 18896
rect 5908 18751 5960 18760
rect 5908 18717 5917 18751
rect 5917 18717 5951 18751
rect 5951 18717 5960 18751
rect 5908 18708 5960 18717
rect 6184 18751 6236 18760
rect 6184 18717 6193 18751
rect 6193 18717 6227 18751
rect 6227 18717 6236 18751
rect 6184 18708 6236 18717
rect 7012 18708 7064 18760
rect 8576 18776 8628 18828
rect 15568 18776 15620 18828
rect 16764 18776 16816 18828
rect 21088 18844 21140 18896
rect 17776 18776 17828 18828
rect 18052 18776 18104 18828
rect 20720 18776 20772 18828
rect 23480 18776 23532 18828
rect 8208 18708 8260 18760
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 14188 18640 14240 18692
rect 15016 18640 15068 18692
rect 5540 18572 5592 18624
rect 5724 18615 5776 18624
rect 5724 18581 5733 18615
rect 5733 18581 5767 18615
rect 5767 18581 5776 18615
rect 5724 18572 5776 18581
rect 14096 18615 14148 18624
rect 14096 18581 14105 18615
rect 14105 18581 14139 18615
rect 14139 18581 14148 18615
rect 14096 18572 14148 18581
rect 17040 18708 17092 18760
rect 20812 18708 20864 18760
rect 19892 18683 19944 18692
rect 15568 18572 15620 18624
rect 15844 18615 15896 18624
rect 15844 18581 15853 18615
rect 15853 18581 15887 18615
rect 15887 18581 15896 18615
rect 15844 18572 15896 18581
rect 16856 18572 16908 18624
rect 19892 18649 19901 18683
rect 19901 18649 19935 18683
rect 19935 18649 19944 18683
rect 19892 18640 19944 18649
rect 21456 18708 21508 18760
rect 23204 18708 23256 18760
rect 26240 18776 26292 18828
rect 28080 18844 28132 18896
rect 26148 18708 26200 18760
rect 27712 18751 27764 18760
rect 27712 18717 27721 18751
rect 27721 18717 27755 18751
rect 27755 18717 27764 18751
rect 27712 18708 27764 18717
rect 28724 18751 28776 18760
rect 28724 18717 28733 18751
rect 28733 18717 28767 18751
rect 28767 18717 28776 18751
rect 28724 18708 28776 18717
rect 21364 18640 21416 18692
rect 18236 18615 18288 18624
rect 18236 18581 18245 18615
rect 18245 18581 18279 18615
rect 18279 18581 18288 18615
rect 18236 18572 18288 18581
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 19432 18572 19484 18624
rect 20352 18615 20404 18624
rect 20352 18581 20361 18615
rect 20361 18581 20395 18615
rect 20395 18581 20404 18615
rect 20352 18572 20404 18581
rect 20904 18572 20956 18624
rect 20996 18572 21048 18624
rect 21824 18572 21876 18624
rect 24676 18572 24728 18624
rect 24952 18572 25004 18624
rect 27068 18572 27120 18624
rect 27160 18572 27212 18624
rect 28172 18572 28224 18624
rect 8034 18470 8086 18522
rect 8098 18470 8150 18522
rect 8162 18470 8214 18522
rect 8226 18470 8278 18522
rect 8290 18470 8342 18522
rect 15118 18470 15170 18522
rect 15182 18470 15234 18522
rect 15246 18470 15298 18522
rect 15310 18470 15362 18522
rect 15374 18470 15426 18522
rect 22202 18470 22254 18522
rect 22266 18470 22318 18522
rect 22330 18470 22382 18522
rect 22394 18470 22446 18522
rect 22458 18470 22510 18522
rect 29286 18470 29338 18522
rect 29350 18470 29402 18522
rect 29414 18470 29466 18522
rect 29478 18470 29530 18522
rect 29542 18470 29594 18522
rect 2504 18368 2556 18420
rect 2596 18300 2648 18352
rect 1584 18232 1636 18284
rect 6920 18368 6972 18420
rect 8392 18368 8444 18420
rect 9496 18368 9548 18420
rect 9680 18368 9732 18420
rect 10416 18368 10468 18420
rect 4988 18343 5040 18352
rect 4988 18309 4997 18343
rect 4997 18309 5031 18343
rect 5031 18309 5040 18343
rect 4988 18300 5040 18309
rect 5172 18300 5224 18352
rect 7288 18300 7340 18352
rect 7472 18232 7524 18284
rect 7656 18275 7708 18284
rect 7656 18241 7665 18275
rect 7665 18241 7699 18275
rect 7699 18241 7708 18275
rect 7656 18232 7708 18241
rect 4988 18096 5040 18148
rect 8392 18232 8444 18284
rect 8576 18232 8628 18284
rect 11980 18300 12032 18352
rect 12072 18275 12124 18284
rect 12072 18241 12081 18275
rect 12081 18241 12115 18275
rect 12115 18241 12124 18275
rect 12072 18232 12124 18241
rect 12624 18164 12676 18216
rect 9220 18096 9272 18148
rect 4344 18028 4396 18080
rect 5264 18071 5316 18080
rect 5264 18037 5273 18071
rect 5273 18037 5307 18071
rect 5307 18037 5316 18071
rect 5264 18028 5316 18037
rect 7748 18071 7800 18080
rect 7748 18037 7757 18071
rect 7757 18037 7791 18071
rect 7791 18037 7800 18071
rect 7748 18028 7800 18037
rect 9956 18028 10008 18080
rect 10876 18028 10928 18080
rect 11060 18028 11112 18080
rect 15568 18368 15620 18420
rect 17776 18411 17828 18420
rect 17776 18377 17785 18411
rect 17785 18377 17819 18411
rect 17819 18377 17828 18411
rect 17776 18368 17828 18377
rect 18328 18368 18380 18420
rect 27712 18368 27764 18420
rect 13268 18300 13320 18352
rect 15476 18300 15528 18352
rect 14648 18275 14700 18284
rect 14648 18241 14657 18275
rect 14657 18241 14691 18275
rect 14691 18241 14700 18275
rect 14648 18232 14700 18241
rect 15016 18275 15068 18284
rect 15016 18241 15025 18275
rect 15025 18241 15059 18275
rect 15059 18241 15068 18275
rect 15016 18232 15068 18241
rect 16856 18275 16908 18284
rect 16856 18241 16865 18275
rect 16865 18241 16899 18275
rect 16899 18241 16908 18275
rect 16856 18232 16908 18241
rect 18144 18300 18196 18352
rect 19984 18300 20036 18352
rect 20352 18232 20404 18284
rect 20812 18300 20864 18352
rect 23112 18300 23164 18352
rect 24952 18300 25004 18352
rect 26516 18300 26568 18352
rect 20904 18232 20956 18284
rect 21456 18232 21508 18284
rect 27160 18275 27212 18284
rect 27160 18241 27169 18275
rect 27169 18241 27203 18275
rect 27203 18241 27212 18275
rect 27160 18232 27212 18241
rect 27528 18232 27580 18284
rect 14372 18164 14424 18216
rect 16580 18164 16632 18216
rect 16948 18207 17000 18216
rect 16948 18173 16957 18207
rect 16957 18173 16991 18207
rect 16991 18173 17000 18207
rect 16948 18164 17000 18173
rect 20812 18207 20864 18216
rect 20812 18173 20821 18207
rect 20821 18173 20855 18207
rect 20855 18173 20864 18207
rect 20812 18164 20864 18173
rect 23756 18207 23808 18216
rect 23756 18173 23765 18207
rect 23765 18173 23799 18207
rect 23799 18173 23808 18207
rect 23756 18164 23808 18173
rect 26700 18164 26752 18216
rect 14004 18071 14056 18080
rect 14004 18037 14013 18071
rect 14013 18037 14047 18071
rect 14047 18037 14056 18071
rect 14004 18028 14056 18037
rect 14280 18028 14332 18080
rect 16764 18028 16816 18080
rect 17316 18028 17368 18080
rect 19892 18028 19944 18080
rect 21088 18071 21140 18080
rect 21088 18037 21097 18071
rect 21097 18037 21131 18071
rect 21131 18037 21140 18071
rect 21088 18028 21140 18037
rect 27068 18071 27120 18080
rect 27068 18037 27077 18071
rect 27077 18037 27111 18071
rect 27111 18037 27120 18071
rect 27068 18028 27120 18037
rect 4492 17926 4544 17978
rect 4556 17926 4608 17978
rect 4620 17926 4672 17978
rect 4684 17926 4736 17978
rect 4748 17926 4800 17978
rect 11576 17926 11628 17978
rect 11640 17926 11692 17978
rect 11704 17926 11756 17978
rect 11768 17926 11820 17978
rect 11832 17926 11884 17978
rect 18660 17926 18712 17978
rect 18724 17926 18776 17978
rect 18788 17926 18840 17978
rect 18852 17926 18904 17978
rect 18916 17926 18968 17978
rect 25744 17926 25796 17978
rect 25808 17926 25860 17978
rect 25872 17926 25924 17978
rect 25936 17926 25988 17978
rect 26000 17926 26052 17978
rect 1584 17799 1636 17808
rect 1584 17765 1593 17799
rect 1593 17765 1627 17799
rect 1627 17765 1636 17799
rect 1584 17756 1636 17765
rect 4160 17799 4212 17808
rect 4160 17765 4169 17799
rect 4169 17765 4203 17799
rect 4203 17765 4212 17799
rect 4160 17756 4212 17765
rect 5264 17756 5316 17808
rect 6552 17756 6604 17808
rect 7012 17824 7064 17876
rect 11888 17824 11940 17876
rect 11980 17824 12032 17876
rect 13820 17824 13872 17876
rect 17776 17824 17828 17876
rect 18052 17824 18104 17876
rect 10600 17756 10652 17808
rect 13544 17756 13596 17808
rect 7288 17731 7340 17740
rect 7288 17697 7297 17731
rect 7297 17697 7331 17731
rect 7331 17697 7340 17731
rect 7288 17688 7340 17697
rect 7748 17688 7800 17740
rect 11060 17731 11112 17740
rect 4436 17620 4488 17672
rect 5724 17663 5776 17672
rect 5724 17629 5733 17663
rect 5733 17629 5767 17663
rect 5767 17629 5776 17663
rect 5724 17620 5776 17629
rect 6368 17663 6420 17672
rect 6368 17629 6377 17663
rect 6377 17629 6411 17663
rect 6411 17629 6420 17663
rect 6368 17620 6420 17629
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 7472 17620 7524 17672
rect 7656 17620 7708 17672
rect 9036 17620 9088 17672
rect 2228 17552 2280 17604
rect 5172 17552 5224 17604
rect 7104 17552 7156 17604
rect 8392 17595 8444 17604
rect 8392 17561 8401 17595
rect 8401 17561 8435 17595
rect 8435 17561 8444 17595
rect 8392 17552 8444 17561
rect 2872 17484 2924 17536
rect 7564 17527 7616 17536
rect 7564 17493 7573 17527
rect 7573 17493 7607 17527
rect 7607 17493 7616 17527
rect 7564 17484 7616 17493
rect 7932 17484 7984 17536
rect 9312 17527 9364 17536
rect 9312 17493 9321 17527
rect 9321 17493 9355 17527
rect 9355 17493 9364 17527
rect 9312 17484 9364 17493
rect 11060 17697 11069 17731
rect 11069 17697 11103 17731
rect 11103 17697 11112 17731
rect 11060 17688 11112 17697
rect 9956 17663 10008 17672
rect 9956 17629 9965 17663
rect 9965 17629 9999 17663
rect 9999 17629 10008 17663
rect 9956 17620 10008 17629
rect 9588 17595 9640 17604
rect 9588 17561 9597 17595
rect 9597 17561 9631 17595
rect 9631 17561 9640 17595
rect 9588 17552 9640 17561
rect 9680 17595 9732 17604
rect 9680 17561 9689 17595
rect 9689 17561 9723 17595
rect 9723 17561 9732 17595
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 12808 17620 12860 17672
rect 13268 17663 13320 17672
rect 13268 17629 13277 17663
rect 13277 17629 13311 17663
rect 13311 17629 13320 17663
rect 13268 17620 13320 17629
rect 14096 17620 14148 17672
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 16580 17688 16632 17740
rect 17132 17731 17184 17740
rect 17132 17697 17141 17731
rect 17141 17697 17175 17731
rect 17175 17697 17184 17731
rect 17132 17688 17184 17697
rect 14464 17595 14516 17604
rect 9680 17552 9732 17561
rect 9772 17484 9824 17536
rect 10692 17484 10744 17536
rect 14464 17561 14473 17595
rect 14473 17561 14507 17595
rect 14507 17561 14516 17595
rect 14464 17552 14516 17561
rect 16304 17552 16356 17604
rect 18696 17824 18748 17876
rect 23388 17824 23440 17876
rect 27804 17824 27856 17876
rect 28724 17867 28776 17876
rect 28724 17833 28733 17867
rect 28733 17833 28767 17867
rect 28767 17833 28776 17867
rect 28724 17824 28776 17833
rect 19248 17756 19300 17808
rect 19340 17663 19392 17672
rect 19340 17629 19349 17663
rect 19349 17629 19383 17663
rect 19383 17629 19392 17663
rect 19340 17620 19392 17629
rect 21732 17620 21784 17672
rect 21548 17552 21600 17604
rect 28356 17756 28408 17808
rect 24584 17620 24636 17672
rect 27896 17688 27948 17740
rect 24952 17663 25004 17672
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 27804 17620 27856 17672
rect 12164 17484 12216 17536
rect 12900 17527 12952 17536
rect 12900 17493 12909 17527
rect 12909 17493 12943 17527
rect 12943 17493 12952 17527
rect 12900 17484 12952 17493
rect 14096 17527 14148 17536
rect 14096 17493 14105 17527
rect 14105 17493 14139 17527
rect 14139 17493 14148 17527
rect 14096 17484 14148 17493
rect 15844 17484 15896 17536
rect 16580 17484 16632 17536
rect 21732 17527 21784 17536
rect 21732 17493 21741 17527
rect 21741 17493 21775 17527
rect 21775 17493 21784 17527
rect 21732 17484 21784 17493
rect 24492 17484 24544 17536
rect 26332 17527 26384 17536
rect 26332 17493 26341 17527
rect 26341 17493 26375 17527
rect 26375 17493 26384 17527
rect 26332 17484 26384 17493
rect 26976 17484 27028 17536
rect 28356 17484 28408 17536
rect 8034 17382 8086 17434
rect 8098 17382 8150 17434
rect 8162 17382 8214 17434
rect 8226 17382 8278 17434
rect 8290 17382 8342 17434
rect 15118 17382 15170 17434
rect 15182 17382 15234 17434
rect 15246 17382 15298 17434
rect 15310 17382 15362 17434
rect 15374 17382 15426 17434
rect 22202 17382 22254 17434
rect 22266 17382 22318 17434
rect 22330 17382 22382 17434
rect 22394 17382 22446 17434
rect 22458 17382 22510 17434
rect 29286 17382 29338 17434
rect 29350 17382 29402 17434
rect 29414 17382 29466 17434
rect 29478 17382 29530 17434
rect 29542 17382 29594 17434
rect 4988 17280 5040 17332
rect 6920 17280 6972 17332
rect 9312 17212 9364 17264
rect 9864 17255 9916 17264
rect 1768 17144 1820 17196
rect 7656 17144 7708 17196
rect 9496 17187 9548 17196
rect 5816 17076 5868 17128
rect 9496 17153 9505 17187
rect 9505 17153 9539 17187
rect 9539 17153 9548 17187
rect 9496 17144 9548 17153
rect 9864 17221 9873 17255
rect 9873 17221 9907 17255
rect 9907 17221 9916 17255
rect 9864 17212 9916 17221
rect 10048 17212 10100 17264
rect 11888 17187 11940 17196
rect 7932 17076 7984 17128
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 12900 17280 12952 17332
rect 14648 17280 14700 17332
rect 15200 17280 15252 17332
rect 17132 17280 17184 17332
rect 21272 17323 21324 17332
rect 21272 17289 21281 17323
rect 21281 17289 21315 17323
rect 21315 17289 21324 17323
rect 21272 17280 21324 17289
rect 22008 17280 22060 17332
rect 23388 17323 23440 17332
rect 23388 17289 23397 17323
rect 23397 17289 23431 17323
rect 23431 17289 23440 17323
rect 23388 17280 23440 17289
rect 27896 17280 27948 17332
rect 23756 17212 23808 17264
rect 12992 17144 13044 17196
rect 13912 17144 13964 17196
rect 19340 17187 19392 17196
rect 19340 17153 19349 17187
rect 19349 17153 19383 17187
rect 19383 17153 19392 17187
rect 19340 17144 19392 17153
rect 6552 17008 6604 17060
rect 8576 17008 8628 17060
rect 15476 17076 15528 17128
rect 18420 17076 18472 17128
rect 20720 17144 20772 17196
rect 21732 17144 21784 17196
rect 22008 17144 22060 17196
rect 22560 17144 22612 17196
rect 21180 17076 21232 17128
rect 23204 17187 23256 17196
rect 23204 17153 23213 17187
rect 23213 17153 23247 17187
rect 23247 17153 23256 17187
rect 27252 17187 27304 17196
rect 23204 17144 23256 17153
rect 27252 17153 27261 17187
rect 27261 17153 27295 17187
rect 27295 17153 27304 17187
rect 27252 17144 27304 17153
rect 27528 17144 27580 17196
rect 23572 17076 23624 17128
rect 13820 17008 13872 17060
rect 15568 17008 15620 17060
rect 17224 17008 17276 17060
rect 26332 17076 26384 17128
rect 27620 17076 27672 17128
rect 24308 17051 24360 17060
rect 24308 17017 24317 17051
rect 24317 17017 24351 17051
rect 24351 17017 24360 17051
rect 24308 17008 24360 17017
rect 1952 16940 2004 16992
rect 5816 16983 5868 16992
rect 5816 16949 5825 16983
rect 5825 16949 5859 16983
rect 5859 16949 5868 16983
rect 5816 16940 5868 16949
rect 6368 16940 6420 16992
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 9588 16940 9640 16992
rect 10692 16940 10744 16992
rect 11428 16940 11480 16992
rect 14096 16940 14148 16992
rect 14280 16940 14332 16992
rect 21640 16940 21692 16992
rect 22652 16940 22704 16992
rect 22928 16983 22980 16992
rect 22928 16949 22937 16983
rect 22937 16949 22971 16983
rect 22971 16949 22980 16983
rect 22928 16940 22980 16949
rect 26792 16940 26844 16992
rect 4492 16838 4544 16890
rect 4556 16838 4608 16890
rect 4620 16838 4672 16890
rect 4684 16838 4736 16890
rect 4748 16838 4800 16890
rect 11576 16838 11628 16890
rect 11640 16838 11692 16890
rect 11704 16838 11756 16890
rect 11768 16838 11820 16890
rect 11832 16838 11884 16890
rect 18660 16838 18712 16890
rect 18724 16838 18776 16890
rect 18788 16838 18840 16890
rect 18852 16838 18904 16890
rect 18916 16838 18968 16890
rect 25744 16838 25796 16890
rect 25808 16838 25860 16890
rect 25872 16838 25924 16890
rect 25936 16838 25988 16890
rect 26000 16838 26052 16890
rect 1768 16779 1820 16788
rect 1768 16745 1777 16779
rect 1777 16745 1811 16779
rect 1811 16745 1820 16779
rect 1768 16736 1820 16745
rect 2872 16779 2924 16788
rect 2872 16745 2881 16779
rect 2881 16745 2915 16779
rect 2915 16745 2924 16779
rect 2872 16736 2924 16745
rect 5172 16779 5224 16788
rect 5172 16745 5181 16779
rect 5181 16745 5215 16779
rect 5215 16745 5224 16779
rect 5172 16736 5224 16745
rect 7012 16736 7064 16788
rect 8392 16736 8444 16788
rect 9496 16779 9548 16788
rect 9496 16745 9505 16779
rect 9505 16745 9539 16779
rect 9539 16745 9548 16779
rect 9496 16736 9548 16745
rect 9864 16736 9916 16788
rect 10048 16736 10100 16788
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 13912 16736 13964 16788
rect 2228 16643 2280 16652
rect 2228 16609 2237 16643
rect 2237 16609 2271 16643
rect 2271 16609 2280 16643
rect 2228 16600 2280 16609
rect 8576 16600 8628 16652
rect 10600 16668 10652 16720
rect 17224 16668 17276 16720
rect 18144 16711 18196 16720
rect 18144 16677 18153 16711
rect 18153 16677 18187 16711
rect 18187 16677 18196 16711
rect 18144 16668 18196 16677
rect 19156 16668 19208 16720
rect 19340 16736 19392 16788
rect 20352 16736 20404 16788
rect 20720 16668 20772 16720
rect 13176 16600 13228 16652
rect 13544 16600 13596 16652
rect 2412 16532 2464 16584
rect 2872 16532 2924 16584
rect 11428 16532 11480 16584
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 12164 16532 12216 16584
rect 12624 16532 12676 16584
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 9864 16507 9916 16516
rect 9864 16473 9873 16507
rect 9873 16473 9907 16507
rect 9907 16473 9916 16507
rect 9864 16464 9916 16473
rect 13268 16532 13320 16584
rect 18236 16532 18288 16584
rect 19616 16532 19668 16584
rect 20904 16600 20956 16652
rect 20628 16532 20680 16584
rect 22928 16668 22980 16720
rect 26424 16736 26476 16788
rect 27436 16736 27488 16788
rect 23756 16600 23808 16652
rect 26792 16668 26844 16720
rect 26240 16600 26292 16652
rect 27252 16600 27304 16652
rect 27620 16643 27672 16652
rect 27620 16609 27629 16643
rect 27629 16609 27663 16643
rect 27663 16609 27672 16643
rect 27620 16600 27672 16609
rect 28080 16600 28132 16652
rect 21364 16575 21416 16584
rect 21364 16541 21373 16575
rect 21373 16541 21407 16575
rect 21407 16541 21416 16575
rect 21364 16532 21416 16541
rect 23388 16532 23440 16584
rect 23572 16532 23624 16584
rect 25320 16532 25372 16584
rect 16488 16464 16540 16516
rect 18604 16464 18656 16516
rect 19248 16464 19300 16516
rect 22560 16464 22612 16516
rect 10048 16396 10100 16448
rect 13820 16396 13872 16448
rect 14556 16396 14608 16448
rect 15200 16396 15252 16448
rect 16396 16396 16448 16448
rect 17316 16396 17368 16448
rect 22100 16396 22152 16448
rect 24768 16439 24820 16448
rect 24768 16405 24777 16439
rect 24777 16405 24811 16439
rect 24811 16405 24820 16439
rect 24768 16396 24820 16405
rect 26424 16439 26476 16448
rect 26424 16405 26433 16439
rect 26433 16405 26467 16439
rect 26467 16405 26476 16439
rect 26424 16396 26476 16405
rect 27436 16532 27488 16584
rect 28724 16575 28776 16584
rect 28724 16541 28733 16575
rect 28733 16541 28767 16575
rect 28767 16541 28776 16575
rect 28724 16532 28776 16541
rect 26792 16507 26844 16516
rect 26792 16473 26801 16507
rect 26801 16473 26835 16507
rect 26835 16473 26844 16507
rect 26792 16464 26844 16473
rect 27344 16464 27396 16516
rect 8034 16294 8086 16346
rect 8098 16294 8150 16346
rect 8162 16294 8214 16346
rect 8226 16294 8278 16346
rect 8290 16294 8342 16346
rect 15118 16294 15170 16346
rect 15182 16294 15234 16346
rect 15246 16294 15298 16346
rect 15310 16294 15362 16346
rect 15374 16294 15426 16346
rect 22202 16294 22254 16346
rect 22266 16294 22318 16346
rect 22330 16294 22382 16346
rect 22394 16294 22446 16346
rect 22458 16294 22510 16346
rect 29286 16294 29338 16346
rect 29350 16294 29402 16346
rect 29414 16294 29466 16346
rect 29478 16294 29530 16346
rect 29542 16294 29594 16346
rect 9036 16192 9088 16244
rect 9864 16192 9916 16244
rect 10048 16235 10100 16244
rect 10048 16201 10057 16235
rect 10057 16201 10091 16235
rect 10091 16201 10100 16235
rect 10048 16192 10100 16201
rect 10416 16192 10468 16244
rect 10968 16192 11020 16244
rect 12532 16192 12584 16244
rect 3792 16167 3844 16176
rect 3792 16133 3801 16167
rect 3801 16133 3835 16167
rect 3835 16133 3844 16167
rect 3792 16124 3844 16133
rect 3976 16167 4028 16176
rect 3976 16133 3985 16167
rect 3985 16133 4019 16167
rect 4019 16133 4028 16167
rect 3976 16124 4028 16133
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 4068 16099 4120 16108
rect 4068 16065 4077 16099
rect 4077 16065 4111 16099
rect 4111 16065 4120 16099
rect 6736 16099 6788 16108
rect 4068 16056 4120 16065
rect 6736 16065 6745 16099
rect 6745 16065 6779 16099
rect 6779 16065 6788 16099
rect 6736 16056 6788 16065
rect 6920 16056 6972 16108
rect 5540 15988 5592 16040
rect 7748 16056 7800 16108
rect 11980 16056 12032 16108
rect 12624 16056 12676 16108
rect 13176 16124 13228 16176
rect 14924 16192 14976 16244
rect 16212 16192 16264 16244
rect 16580 16192 16632 16244
rect 18236 16192 18288 16244
rect 22928 16192 22980 16244
rect 23664 16192 23716 16244
rect 24032 16192 24084 16244
rect 25044 16192 25096 16244
rect 27068 16192 27120 16244
rect 15016 16167 15068 16176
rect 15016 16133 15025 16167
rect 15025 16133 15059 16167
rect 15059 16133 15068 16167
rect 15016 16124 15068 16133
rect 17224 16124 17276 16176
rect 12900 15988 12952 16040
rect 7472 15920 7524 15972
rect 7656 15963 7708 15972
rect 7656 15929 7665 15963
rect 7665 15929 7699 15963
rect 7699 15929 7708 15963
rect 7656 15920 7708 15929
rect 7748 15920 7800 15972
rect 10784 15920 10836 15972
rect 12808 15920 12860 15972
rect 13268 16056 13320 16108
rect 13544 16056 13596 16108
rect 13912 16099 13964 16108
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 13912 16056 13964 16065
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 24768 16124 24820 16176
rect 19064 16056 19116 16108
rect 20352 16056 20404 16108
rect 21364 16056 21416 16108
rect 17316 16031 17368 16040
rect 17316 15997 17325 16031
rect 17325 15997 17359 16031
rect 17359 15997 17368 16031
rect 17316 15988 17368 15997
rect 18144 15988 18196 16040
rect 5264 15852 5316 15904
rect 6184 15852 6236 15904
rect 11980 15852 12032 15904
rect 12992 15895 13044 15904
rect 12992 15861 13001 15895
rect 13001 15861 13035 15895
rect 13035 15861 13044 15895
rect 12992 15852 13044 15861
rect 14464 15852 14516 15904
rect 14648 15895 14700 15904
rect 14648 15861 14657 15895
rect 14657 15861 14691 15895
rect 14691 15861 14700 15895
rect 14648 15852 14700 15861
rect 16212 15920 16264 15972
rect 19156 15988 19208 16040
rect 19616 15920 19668 15972
rect 23020 16056 23072 16108
rect 24308 16056 24360 16108
rect 20536 15920 20588 15972
rect 23664 15988 23716 16040
rect 27712 16056 27764 16108
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 27252 15988 27304 16040
rect 28080 15988 28132 16040
rect 28264 15988 28316 16040
rect 25412 15852 25464 15904
rect 4492 15750 4544 15802
rect 4556 15750 4608 15802
rect 4620 15750 4672 15802
rect 4684 15750 4736 15802
rect 4748 15750 4800 15802
rect 11576 15750 11628 15802
rect 11640 15750 11692 15802
rect 11704 15750 11756 15802
rect 11768 15750 11820 15802
rect 11832 15750 11884 15802
rect 18660 15750 18712 15802
rect 18724 15750 18776 15802
rect 18788 15750 18840 15802
rect 18852 15750 18904 15802
rect 18916 15750 18968 15802
rect 25744 15750 25796 15802
rect 25808 15750 25860 15802
rect 25872 15750 25924 15802
rect 25936 15750 25988 15802
rect 26000 15750 26052 15802
rect 4620 15648 4672 15700
rect 5172 15648 5224 15700
rect 5632 15691 5684 15700
rect 5632 15657 5641 15691
rect 5641 15657 5675 15691
rect 5675 15657 5684 15691
rect 5632 15648 5684 15657
rect 9680 15648 9732 15700
rect 16396 15691 16448 15700
rect 16396 15657 16405 15691
rect 16405 15657 16439 15691
rect 16439 15657 16448 15691
rect 16396 15648 16448 15657
rect 16488 15648 16540 15700
rect 19616 15648 19668 15700
rect 19892 15648 19944 15700
rect 20260 15648 20312 15700
rect 23020 15648 23072 15700
rect 23388 15648 23440 15700
rect 28724 15691 28776 15700
rect 28724 15657 28733 15691
rect 28733 15657 28767 15691
rect 28767 15657 28776 15691
rect 28724 15648 28776 15657
rect 15568 15580 15620 15632
rect 6184 15555 6236 15564
rect 6184 15521 6193 15555
rect 6193 15521 6227 15555
rect 6227 15521 6236 15555
rect 6184 15512 6236 15521
rect 14648 15512 14700 15564
rect 18052 15580 18104 15632
rect 24584 15580 24636 15632
rect 23388 15512 23440 15564
rect 23940 15512 23992 15564
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3792 15444 3844 15453
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 10692 15444 10744 15496
rect 15476 15487 15528 15496
rect 3976 15376 4028 15428
rect 5172 15376 5224 15428
rect 15476 15453 15485 15487
rect 15485 15453 15519 15487
rect 15519 15453 15528 15487
rect 15476 15444 15528 15453
rect 16672 15444 16724 15496
rect 17408 15444 17460 15496
rect 21364 15444 21416 15496
rect 25044 15444 25096 15496
rect 25412 15487 25464 15496
rect 25412 15453 25421 15487
rect 25421 15453 25455 15487
rect 25455 15453 25464 15487
rect 25412 15444 25464 15453
rect 27252 15487 27304 15496
rect 27252 15453 27261 15487
rect 27261 15453 27295 15487
rect 27295 15453 27304 15487
rect 27252 15444 27304 15453
rect 17960 15376 18012 15428
rect 18236 15419 18288 15428
rect 18236 15385 18245 15419
rect 18245 15385 18279 15419
rect 18279 15385 18288 15419
rect 18236 15376 18288 15385
rect 9312 15308 9364 15360
rect 12164 15351 12216 15360
rect 12164 15317 12173 15351
rect 12173 15317 12207 15351
rect 12207 15317 12216 15351
rect 12164 15308 12216 15317
rect 13912 15308 13964 15360
rect 15016 15308 15068 15360
rect 16764 15308 16816 15360
rect 17224 15308 17276 15360
rect 19064 15308 19116 15360
rect 23940 15308 23992 15360
rect 24584 15308 24636 15360
rect 24860 15308 24912 15360
rect 27528 15351 27580 15360
rect 27528 15317 27537 15351
rect 27537 15317 27571 15351
rect 27571 15317 27580 15351
rect 27528 15308 27580 15317
rect 8034 15206 8086 15258
rect 8098 15206 8150 15258
rect 8162 15206 8214 15258
rect 8226 15206 8278 15258
rect 8290 15206 8342 15258
rect 15118 15206 15170 15258
rect 15182 15206 15234 15258
rect 15246 15206 15298 15258
rect 15310 15206 15362 15258
rect 15374 15206 15426 15258
rect 22202 15206 22254 15258
rect 22266 15206 22318 15258
rect 22330 15206 22382 15258
rect 22394 15206 22446 15258
rect 22458 15206 22510 15258
rect 29286 15206 29338 15258
rect 29350 15206 29402 15258
rect 29414 15206 29466 15258
rect 29478 15206 29530 15258
rect 29542 15206 29594 15258
rect 4068 15104 4120 15156
rect 5172 15036 5224 15088
rect 5540 15104 5592 15156
rect 6736 15104 6788 15156
rect 9680 15104 9732 15156
rect 11980 15104 12032 15156
rect 13452 15104 13504 15156
rect 16764 15147 16816 15156
rect 5632 15036 5684 15088
rect 7472 15036 7524 15088
rect 9772 15036 9824 15088
rect 12900 15036 12952 15088
rect 4344 14968 4396 15020
rect 7104 14968 7156 15020
rect 9128 14968 9180 15020
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 4896 14900 4948 14952
rect 5356 14832 5408 14884
rect 7564 14832 7616 14884
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 5080 14764 5132 14816
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 9312 14764 9364 14816
rect 10600 14968 10652 15020
rect 10232 14900 10284 14952
rect 10876 14968 10928 15020
rect 11428 14968 11480 15020
rect 12992 14968 13044 15020
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 14004 15011 14056 15020
rect 14004 14977 14013 15011
rect 14013 14977 14047 15011
rect 14047 14977 14056 15011
rect 14004 14968 14056 14977
rect 16764 15113 16773 15147
rect 16773 15113 16807 15147
rect 16807 15113 16816 15147
rect 16764 15104 16816 15113
rect 18236 15104 18288 15156
rect 14648 14968 14700 15020
rect 12164 14900 12216 14952
rect 17592 15036 17644 15088
rect 21272 15104 21324 15156
rect 24768 15104 24820 15156
rect 27344 15147 27396 15156
rect 27344 15113 27353 15147
rect 27353 15113 27387 15147
rect 27387 15113 27396 15147
rect 27344 15104 27396 15113
rect 17408 14968 17460 15020
rect 17960 15011 18012 15020
rect 17960 14977 17969 15011
rect 17969 14977 18003 15011
rect 18003 14977 18012 15011
rect 17960 14968 18012 14977
rect 18420 14968 18472 15020
rect 20260 14968 20312 15020
rect 20812 15036 20864 15088
rect 21640 14968 21692 15020
rect 24308 14968 24360 15020
rect 17316 14943 17368 14952
rect 17316 14909 17325 14943
rect 17325 14909 17359 14943
rect 17359 14909 17368 14943
rect 17316 14900 17368 14909
rect 21088 14943 21140 14952
rect 10692 14832 10744 14884
rect 18052 14875 18104 14884
rect 18052 14841 18061 14875
rect 18061 14841 18095 14875
rect 18095 14841 18104 14875
rect 18052 14832 18104 14841
rect 20628 14832 20680 14884
rect 21088 14909 21097 14943
rect 21097 14909 21131 14943
rect 21131 14909 21140 14943
rect 21088 14900 21140 14909
rect 27344 14968 27396 15020
rect 10140 14764 10192 14816
rect 10968 14807 11020 14816
rect 10968 14773 10977 14807
rect 10977 14773 11011 14807
rect 11011 14773 11020 14807
rect 10968 14764 11020 14773
rect 11336 14764 11388 14816
rect 15660 14764 15712 14816
rect 16304 14764 16356 14816
rect 24308 14832 24360 14884
rect 25504 14900 25556 14952
rect 27436 14943 27488 14952
rect 27436 14909 27445 14943
rect 27445 14909 27479 14943
rect 27479 14909 27488 14943
rect 27436 14900 27488 14909
rect 27528 14943 27580 14952
rect 27528 14909 27537 14943
rect 27537 14909 27571 14943
rect 27571 14909 27580 14943
rect 27528 14900 27580 14909
rect 25228 14832 25280 14884
rect 23572 14764 23624 14816
rect 28264 14764 28316 14816
rect 4492 14662 4544 14714
rect 4556 14662 4608 14714
rect 4620 14662 4672 14714
rect 4684 14662 4736 14714
rect 4748 14662 4800 14714
rect 11576 14662 11628 14714
rect 11640 14662 11692 14714
rect 11704 14662 11756 14714
rect 11768 14662 11820 14714
rect 11832 14662 11884 14714
rect 18660 14662 18712 14714
rect 18724 14662 18776 14714
rect 18788 14662 18840 14714
rect 18852 14662 18904 14714
rect 18916 14662 18968 14714
rect 25744 14662 25796 14714
rect 25808 14662 25860 14714
rect 25872 14662 25924 14714
rect 25936 14662 25988 14714
rect 26000 14662 26052 14714
rect 4344 14560 4396 14612
rect 4988 14560 5040 14612
rect 6920 14560 6972 14612
rect 7564 14560 7616 14612
rect 9496 14603 9548 14612
rect 9496 14569 9505 14603
rect 9505 14569 9539 14603
rect 9539 14569 9548 14603
rect 9496 14560 9548 14569
rect 10232 14560 10284 14612
rect 10876 14560 10928 14612
rect 13544 14560 13596 14612
rect 18420 14603 18472 14612
rect 6828 14492 6880 14544
rect 18420 14569 18429 14603
rect 18429 14569 18463 14603
rect 18463 14569 18472 14603
rect 18420 14560 18472 14569
rect 19248 14560 19300 14612
rect 23940 14560 23992 14612
rect 24308 14560 24360 14612
rect 26148 14560 26200 14612
rect 27804 14560 27856 14612
rect 22744 14492 22796 14544
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 9588 14424 9640 14476
rect 2136 14356 2188 14365
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 4896 14356 4948 14408
rect 5264 14356 5316 14408
rect 6460 14399 6512 14408
rect 6460 14365 6469 14399
rect 6469 14365 6503 14399
rect 6503 14365 6512 14399
rect 6460 14356 6512 14365
rect 6644 14356 6696 14408
rect 7104 14399 7156 14408
rect 7104 14365 7113 14399
rect 7113 14365 7147 14399
rect 7147 14365 7156 14399
rect 7104 14356 7156 14365
rect 9680 14356 9732 14408
rect 10140 14399 10192 14408
rect 10140 14365 10149 14399
rect 10149 14365 10183 14399
rect 10183 14365 10192 14399
rect 10140 14356 10192 14365
rect 10968 14424 11020 14476
rect 19892 14467 19944 14476
rect 9312 14331 9364 14340
rect 1860 14220 1912 14272
rect 4252 14220 4304 14272
rect 6184 14263 6236 14272
rect 6184 14229 6193 14263
rect 6193 14229 6227 14263
rect 6227 14229 6236 14263
rect 6184 14220 6236 14229
rect 7840 14220 7892 14272
rect 9312 14297 9321 14331
rect 9321 14297 9355 14331
rect 9355 14297 9364 14331
rect 9312 14288 9364 14297
rect 10508 14399 10560 14408
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 11336 14399 11388 14408
rect 10508 14356 10560 14365
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 11612 14399 11664 14408
rect 11612 14365 11621 14399
rect 11621 14365 11655 14399
rect 11655 14365 11664 14399
rect 11612 14356 11664 14365
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 19892 14433 19901 14467
rect 19901 14433 19935 14467
rect 19935 14433 19944 14467
rect 19892 14424 19944 14433
rect 20628 14467 20680 14476
rect 20628 14433 20637 14467
rect 20637 14433 20671 14467
rect 20671 14433 20680 14467
rect 20628 14424 20680 14433
rect 21732 14424 21784 14476
rect 27344 14492 27396 14544
rect 15568 14399 15620 14408
rect 11980 14288 12032 14340
rect 15568 14365 15577 14399
rect 15577 14365 15611 14399
rect 15611 14365 15620 14399
rect 15568 14356 15620 14365
rect 14648 14288 14700 14340
rect 15476 14288 15528 14340
rect 17040 14356 17092 14408
rect 20904 14399 20956 14408
rect 17316 14288 17368 14340
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 24768 14424 24820 14476
rect 25044 14467 25096 14476
rect 25044 14433 25053 14467
rect 25053 14433 25087 14467
rect 25087 14433 25096 14467
rect 25044 14424 25096 14433
rect 20904 14356 20956 14365
rect 20812 14288 20864 14340
rect 21088 14288 21140 14340
rect 21732 14331 21784 14340
rect 21732 14297 21741 14331
rect 21741 14297 21775 14331
rect 21775 14297 21784 14331
rect 23940 14356 23992 14408
rect 24584 14399 24636 14408
rect 24584 14365 24601 14399
rect 24601 14365 24636 14399
rect 24584 14356 24636 14365
rect 24860 14399 24912 14408
rect 24860 14365 24869 14399
rect 24869 14365 24903 14399
rect 24903 14365 24912 14399
rect 24860 14356 24912 14365
rect 27896 14424 27948 14476
rect 21732 14288 21784 14297
rect 9588 14220 9640 14272
rect 10876 14220 10928 14272
rect 11612 14220 11664 14272
rect 12624 14220 12676 14272
rect 20076 14220 20128 14272
rect 21180 14220 21232 14272
rect 24308 14288 24360 14340
rect 25596 14288 25648 14340
rect 26332 14288 26384 14340
rect 22560 14220 22612 14272
rect 25320 14220 25372 14272
rect 27620 14220 27672 14272
rect 8034 14118 8086 14170
rect 8098 14118 8150 14170
rect 8162 14118 8214 14170
rect 8226 14118 8278 14170
rect 8290 14118 8342 14170
rect 15118 14118 15170 14170
rect 15182 14118 15234 14170
rect 15246 14118 15298 14170
rect 15310 14118 15362 14170
rect 15374 14118 15426 14170
rect 22202 14118 22254 14170
rect 22266 14118 22318 14170
rect 22330 14118 22382 14170
rect 22394 14118 22446 14170
rect 22458 14118 22510 14170
rect 29286 14118 29338 14170
rect 29350 14118 29402 14170
rect 29414 14118 29466 14170
rect 29478 14118 29530 14170
rect 29542 14118 29594 14170
rect 4620 14016 4672 14068
rect 4528 13948 4580 14000
rect 5264 14016 5316 14068
rect 9680 14016 9732 14068
rect 10600 14059 10652 14068
rect 10600 14025 10609 14059
rect 10609 14025 10643 14059
rect 10643 14025 10652 14059
rect 10600 14016 10652 14025
rect 11520 14016 11572 14068
rect 15384 14016 15436 14068
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 20628 14016 20680 14068
rect 20812 14016 20864 14068
rect 21088 14016 21140 14068
rect 6920 13991 6972 14000
rect 6920 13957 6929 13991
rect 6929 13957 6963 13991
rect 6963 13957 6972 13991
rect 7564 13991 7616 14000
rect 6920 13948 6972 13957
rect 7564 13957 7573 13991
rect 7573 13957 7607 13991
rect 7607 13957 7616 13991
rect 7564 13948 7616 13957
rect 10140 13948 10192 14000
rect 14004 13948 14056 14000
rect 23572 14016 23624 14068
rect 24308 14016 24360 14068
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 5816 13880 5868 13932
rect 6828 13923 6880 13932
rect 6828 13889 6837 13923
rect 6837 13889 6871 13923
rect 6871 13889 6880 13923
rect 6828 13880 6880 13889
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 9496 13880 9548 13932
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 8392 13812 8444 13864
rect 9312 13812 9364 13864
rect 9772 13812 9824 13864
rect 9956 13812 10008 13864
rect 10140 13855 10192 13864
rect 10140 13821 10149 13855
rect 10149 13821 10183 13855
rect 10183 13821 10192 13855
rect 10140 13812 10192 13821
rect 9588 13744 9640 13796
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 14280 13880 14332 13932
rect 15844 13880 15896 13932
rect 19892 13923 19944 13932
rect 19892 13889 19901 13923
rect 19901 13889 19935 13923
rect 19935 13889 19944 13923
rect 19892 13880 19944 13889
rect 20444 13880 20496 13932
rect 10416 13812 10468 13821
rect 12624 13812 12676 13864
rect 12808 13812 12860 13864
rect 19340 13812 19392 13864
rect 20260 13812 20312 13864
rect 21272 13880 21324 13932
rect 24032 13948 24084 14000
rect 24492 13991 24544 14000
rect 24492 13957 24501 13991
rect 24501 13957 24535 13991
rect 24535 13957 24544 13991
rect 24492 13948 24544 13957
rect 24768 14016 24820 14068
rect 28632 14059 28684 14068
rect 20812 13855 20864 13864
rect 20812 13821 20821 13855
rect 20821 13821 20855 13855
rect 20855 13821 20864 13855
rect 20812 13812 20864 13821
rect 11520 13787 11572 13796
rect 11520 13753 11529 13787
rect 11529 13753 11563 13787
rect 11563 13753 11572 13787
rect 11520 13744 11572 13753
rect 21272 13744 21324 13796
rect 21824 13744 21876 13796
rect 24676 13923 24728 13932
rect 28632 14025 28641 14059
rect 28641 14025 28675 14059
rect 28675 14025 28684 14059
rect 28632 14016 28684 14025
rect 27436 13991 27488 14000
rect 27436 13957 27445 13991
rect 27445 13957 27479 13991
rect 27479 13957 27488 13991
rect 27436 13948 27488 13957
rect 24676 13889 24711 13923
rect 24711 13889 24728 13923
rect 24676 13880 24728 13889
rect 27344 13880 27396 13932
rect 28264 13880 28316 13932
rect 28448 13923 28500 13932
rect 28448 13889 28457 13923
rect 28457 13889 28491 13923
rect 28491 13889 28500 13923
rect 28448 13880 28500 13889
rect 26516 13812 26568 13864
rect 28080 13812 28132 13864
rect 24584 13744 24636 13796
rect 27620 13787 27672 13796
rect 27620 13753 27629 13787
rect 27629 13753 27663 13787
rect 27663 13753 27672 13787
rect 27620 13744 27672 13753
rect 2136 13676 2188 13728
rect 10600 13676 10652 13728
rect 11612 13676 11664 13728
rect 14740 13676 14792 13728
rect 20444 13719 20496 13728
rect 20444 13685 20453 13719
rect 20453 13685 20487 13719
rect 20487 13685 20496 13719
rect 20444 13676 20496 13685
rect 23020 13719 23072 13728
rect 23020 13685 23029 13719
rect 23029 13685 23063 13719
rect 23063 13685 23072 13719
rect 23020 13676 23072 13685
rect 24216 13719 24268 13728
rect 24216 13685 24225 13719
rect 24225 13685 24259 13719
rect 24259 13685 24268 13719
rect 24216 13676 24268 13685
rect 4492 13574 4544 13626
rect 4556 13574 4608 13626
rect 4620 13574 4672 13626
rect 4684 13574 4736 13626
rect 4748 13574 4800 13626
rect 11576 13574 11628 13626
rect 11640 13574 11692 13626
rect 11704 13574 11756 13626
rect 11768 13574 11820 13626
rect 11832 13574 11884 13626
rect 18660 13574 18712 13626
rect 18724 13574 18776 13626
rect 18788 13574 18840 13626
rect 18852 13574 18904 13626
rect 18916 13574 18968 13626
rect 25744 13574 25796 13626
rect 25808 13574 25860 13626
rect 25872 13574 25924 13626
rect 25936 13574 25988 13626
rect 26000 13574 26052 13626
rect 10416 13472 10468 13524
rect 10508 13472 10560 13524
rect 10968 13472 11020 13524
rect 14372 13472 14424 13524
rect 24216 13472 24268 13524
rect 25596 13472 25648 13524
rect 26516 13515 26568 13524
rect 26516 13481 26525 13515
rect 26525 13481 26559 13515
rect 26559 13481 26568 13515
rect 26516 13472 26568 13481
rect 28448 13472 28500 13524
rect 12808 13404 12860 13456
rect 13176 13404 13228 13456
rect 19340 13447 19392 13456
rect 19340 13413 19349 13447
rect 19349 13413 19383 13447
rect 19383 13413 19392 13447
rect 19340 13404 19392 13413
rect 20260 13447 20312 13456
rect 20260 13413 20269 13447
rect 20269 13413 20303 13447
rect 20303 13413 20312 13447
rect 20260 13404 20312 13413
rect 22744 13447 22796 13456
rect 22744 13413 22753 13447
rect 22753 13413 22787 13447
rect 22787 13413 22796 13447
rect 22744 13404 22796 13413
rect 23940 13404 23992 13456
rect 24768 13404 24820 13456
rect 7012 13336 7064 13388
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 7472 13268 7524 13320
rect 8576 13336 8628 13388
rect 20444 13336 20496 13388
rect 10324 13268 10376 13320
rect 12716 13268 12768 13320
rect 13360 13268 13412 13320
rect 13452 13268 13504 13320
rect 18144 13268 18196 13320
rect 21180 13311 21232 13320
rect 21180 13277 21189 13311
rect 21189 13277 21223 13311
rect 21223 13277 21232 13311
rect 21180 13268 21232 13277
rect 21364 13311 21416 13320
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 22560 13268 22612 13320
rect 23020 13268 23072 13320
rect 8668 13200 8720 13252
rect 9588 13200 9640 13252
rect 24308 13268 24360 13320
rect 25504 13268 25556 13320
rect 26240 13268 26292 13320
rect 26608 13311 26660 13320
rect 26608 13277 26617 13311
rect 26617 13277 26651 13311
rect 26651 13277 26660 13311
rect 26608 13268 26660 13277
rect 2688 13132 2740 13184
rect 6828 13132 6880 13184
rect 8484 13132 8536 13184
rect 17316 13200 17368 13252
rect 23480 13200 23532 13252
rect 12624 13132 12676 13184
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 20536 13132 20588 13184
rect 23020 13175 23072 13184
rect 23020 13141 23029 13175
rect 23029 13141 23063 13175
rect 23063 13141 23072 13175
rect 23020 13132 23072 13141
rect 23204 13132 23256 13184
rect 24584 13132 24636 13184
rect 28172 13132 28224 13184
rect 8034 13030 8086 13082
rect 8098 13030 8150 13082
rect 8162 13030 8214 13082
rect 8226 13030 8278 13082
rect 8290 13030 8342 13082
rect 15118 13030 15170 13082
rect 15182 13030 15234 13082
rect 15246 13030 15298 13082
rect 15310 13030 15362 13082
rect 15374 13030 15426 13082
rect 22202 13030 22254 13082
rect 22266 13030 22318 13082
rect 22330 13030 22382 13082
rect 22394 13030 22446 13082
rect 22458 13030 22510 13082
rect 29286 13030 29338 13082
rect 29350 13030 29402 13082
rect 29414 13030 29466 13082
rect 29478 13030 29530 13082
rect 29542 13030 29594 13082
rect 7472 12971 7524 12980
rect 7472 12937 7481 12971
rect 7481 12937 7515 12971
rect 7515 12937 7524 12971
rect 7472 12928 7524 12937
rect 10324 12971 10376 12980
rect 6000 12860 6052 12912
rect 8392 12903 8444 12912
rect 8392 12869 8401 12903
rect 8401 12869 8435 12903
rect 8435 12869 8444 12903
rect 8392 12860 8444 12869
rect 6920 12792 6972 12844
rect 7288 12792 7340 12844
rect 8484 12792 8536 12844
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 9036 12835 9088 12844
rect 8852 12792 8904 12801
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 7012 12656 7064 12708
rect 5908 12588 5960 12640
rect 8668 12724 8720 12776
rect 10324 12937 10333 12971
rect 10333 12937 10367 12971
rect 10367 12937 10376 12971
rect 10324 12928 10376 12937
rect 14372 12928 14424 12980
rect 14464 12928 14516 12980
rect 14648 12971 14700 12980
rect 14648 12937 14657 12971
rect 14657 12937 14691 12971
rect 14691 12937 14700 12971
rect 14648 12928 14700 12937
rect 14740 12928 14792 12980
rect 17040 12928 17092 12980
rect 11980 12903 12032 12912
rect 10600 12835 10652 12844
rect 10600 12801 10609 12835
rect 10609 12801 10643 12835
rect 10643 12801 10652 12835
rect 10600 12792 10652 12801
rect 11980 12869 11989 12903
rect 11989 12869 12023 12903
rect 12023 12869 12032 12903
rect 11980 12860 12032 12869
rect 7840 12656 7892 12708
rect 8852 12656 8904 12708
rect 12072 12792 12124 12844
rect 13452 12835 13504 12844
rect 13452 12801 13461 12835
rect 13461 12801 13495 12835
rect 13495 12801 13504 12835
rect 13452 12792 13504 12801
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 16488 12792 16540 12844
rect 12808 12724 12860 12776
rect 15384 12767 15436 12776
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 19064 12928 19116 12980
rect 18328 12860 18380 12912
rect 20260 12928 20312 12980
rect 20812 12928 20864 12980
rect 23020 12928 23072 12980
rect 24768 12928 24820 12980
rect 26608 12928 26660 12980
rect 26884 12928 26936 12980
rect 27712 12928 27764 12980
rect 20904 12903 20956 12912
rect 18512 12792 18564 12844
rect 19248 12792 19300 12844
rect 20904 12869 20913 12903
rect 20913 12869 20947 12903
rect 20947 12869 20956 12903
rect 20904 12860 20956 12869
rect 22744 12860 22796 12912
rect 21088 12835 21140 12844
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 23480 12860 23532 12912
rect 23664 12860 23716 12912
rect 23572 12792 23624 12844
rect 25136 12835 25188 12844
rect 25136 12801 25145 12835
rect 25145 12801 25179 12835
rect 25179 12801 25188 12835
rect 25136 12792 25188 12801
rect 26240 12792 26292 12844
rect 27252 12792 27304 12844
rect 27528 12792 27580 12844
rect 23480 12767 23532 12776
rect 15016 12656 15068 12708
rect 18328 12656 18380 12708
rect 20904 12656 20956 12708
rect 9956 12588 10008 12640
rect 13544 12631 13596 12640
rect 13544 12597 13553 12631
rect 13553 12597 13587 12631
rect 13587 12597 13596 12631
rect 13544 12588 13596 12597
rect 15108 12588 15160 12640
rect 16028 12588 16080 12640
rect 18512 12631 18564 12640
rect 18512 12597 18521 12631
rect 18521 12597 18555 12631
rect 18555 12597 18564 12631
rect 18512 12588 18564 12597
rect 20076 12588 20128 12640
rect 20260 12588 20312 12640
rect 23480 12733 23489 12767
rect 23489 12733 23523 12767
rect 23523 12733 23532 12767
rect 23480 12724 23532 12733
rect 27712 12767 27764 12776
rect 27712 12733 27721 12767
rect 27721 12733 27755 12767
rect 27755 12733 27764 12767
rect 27712 12724 27764 12733
rect 27896 12792 27948 12844
rect 28172 12792 28224 12844
rect 28264 12724 28316 12776
rect 21364 12656 21416 12708
rect 24584 12588 24636 12640
rect 28632 12631 28684 12640
rect 28632 12597 28641 12631
rect 28641 12597 28675 12631
rect 28675 12597 28684 12631
rect 28632 12588 28684 12597
rect 4492 12486 4544 12538
rect 4556 12486 4608 12538
rect 4620 12486 4672 12538
rect 4684 12486 4736 12538
rect 4748 12486 4800 12538
rect 11576 12486 11628 12538
rect 11640 12486 11692 12538
rect 11704 12486 11756 12538
rect 11768 12486 11820 12538
rect 11832 12486 11884 12538
rect 18660 12486 18712 12538
rect 18724 12486 18776 12538
rect 18788 12486 18840 12538
rect 18852 12486 18904 12538
rect 18916 12486 18968 12538
rect 25744 12486 25796 12538
rect 25808 12486 25860 12538
rect 25872 12486 25924 12538
rect 25936 12486 25988 12538
rect 26000 12486 26052 12538
rect 7472 12427 7524 12436
rect 7472 12393 7481 12427
rect 7481 12393 7515 12427
rect 7515 12393 7524 12427
rect 7472 12384 7524 12393
rect 11704 12384 11756 12436
rect 12072 12427 12124 12436
rect 12072 12393 12081 12427
rect 12081 12393 12115 12427
rect 12115 12393 12124 12427
rect 12072 12384 12124 12393
rect 1768 12248 1820 12300
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 4712 12316 4764 12368
rect 4988 12248 5040 12300
rect 5264 12223 5316 12232
rect 5264 12189 5273 12223
rect 5273 12189 5307 12223
rect 5307 12189 5316 12223
rect 5264 12180 5316 12189
rect 5816 12223 5868 12232
rect 4252 12112 4304 12164
rect 5816 12189 5825 12223
rect 5825 12189 5859 12223
rect 5859 12189 5868 12223
rect 5816 12180 5868 12189
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 7380 12180 7432 12232
rect 9956 12316 10008 12368
rect 14464 12384 14516 12436
rect 2596 12044 2648 12096
rect 4344 12044 4396 12096
rect 7012 12112 7064 12164
rect 9772 12180 9824 12232
rect 10048 12180 10100 12232
rect 10692 12180 10744 12232
rect 10784 12180 10836 12232
rect 10968 12180 11020 12232
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11520 12223 11572 12232
rect 11336 12180 11388 12189
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 11704 12180 11756 12232
rect 15108 12359 15160 12368
rect 15108 12325 15117 12359
rect 15117 12325 15151 12359
rect 15151 12325 15160 12359
rect 15108 12316 15160 12325
rect 15844 12384 15896 12436
rect 16488 12384 16540 12436
rect 18512 12384 18564 12436
rect 19524 12384 19576 12436
rect 20076 12384 20128 12436
rect 20260 12384 20312 12436
rect 26148 12427 26200 12436
rect 26148 12393 26157 12427
rect 26157 12393 26191 12427
rect 26191 12393 26200 12427
rect 26148 12384 26200 12393
rect 10140 12155 10192 12164
rect 6736 12044 6788 12096
rect 7932 12044 7984 12096
rect 10140 12121 10149 12155
rect 10149 12121 10183 12155
rect 10183 12121 10192 12155
rect 10140 12112 10192 12121
rect 9680 12044 9732 12096
rect 11520 12044 11572 12096
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 12992 12180 13044 12232
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 13820 12180 13872 12232
rect 15384 12248 15436 12300
rect 14556 12112 14608 12164
rect 15568 12180 15620 12232
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 16396 12316 16448 12368
rect 22100 12316 22152 12368
rect 15384 12112 15436 12164
rect 16488 12180 16540 12232
rect 17868 12112 17920 12164
rect 19340 12180 19392 12232
rect 19524 12180 19576 12232
rect 20812 12112 20864 12164
rect 22100 12112 22152 12164
rect 22836 12112 22888 12164
rect 13636 12044 13688 12096
rect 14740 12044 14792 12096
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 17776 12087 17828 12096
rect 17776 12053 17785 12087
rect 17785 12053 17819 12087
rect 17819 12053 17828 12087
rect 17776 12044 17828 12053
rect 18512 12044 18564 12096
rect 19248 12087 19300 12096
rect 19248 12053 19257 12087
rect 19257 12053 19291 12087
rect 19291 12053 19300 12087
rect 19248 12044 19300 12053
rect 19340 12044 19392 12096
rect 24860 12248 24912 12300
rect 25504 12291 25556 12300
rect 25504 12257 25513 12291
rect 25513 12257 25547 12291
rect 25547 12257 25556 12291
rect 25504 12248 25556 12257
rect 28172 12316 28224 12368
rect 25228 12223 25280 12232
rect 25228 12189 25237 12223
rect 25237 12189 25271 12223
rect 25271 12189 25280 12223
rect 25228 12180 25280 12189
rect 26148 12180 26200 12232
rect 24676 12112 24728 12164
rect 26700 12155 26752 12164
rect 24032 12044 24084 12096
rect 26700 12121 26709 12155
rect 26709 12121 26743 12155
rect 26743 12121 26752 12155
rect 26700 12112 26752 12121
rect 28080 12248 28132 12300
rect 28356 12112 28408 12164
rect 26148 12044 26200 12096
rect 27620 12044 27672 12096
rect 8034 11942 8086 11994
rect 8098 11942 8150 11994
rect 8162 11942 8214 11994
rect 8226 11942 8278 11994
rect 8290 11942 8342 11994
rect 15118 11942 15170 11994
rect 15182 11942 15234 11994
rect 15246 11942 15298 11994
rect 15310 11942 15362 11994
rect 15374 11942 15426 11994
rect 22202 11942 22254 11994
rect 22266 11942 22318 11994
rect 22330 11942 22382 11994
rect 22394 11942 22446 11994
rect 22458 11942 22510 11994
rect 29286 11942 29338 11994
rect 29350 11942 29402 11994
rect 29414 11942 29466 11994
rect 29478 11942 29530 11994
rect 29542 11942 29594 11994
rect 3056 11840 3108 11892
rect 5264 11840 5316 11892
rect 5816 11840 5868 11892
rect 7012 11840 7064 11892
rect 8760 11840 8812 11892
rect 9772 11840 9824 11892
rect 10324 11840 10376 11892
rect 11520 11883 11572 11892
rect 11520 11849 11529 11883
rect 11529 11849 11563 11883
rect 11563 11849 11572 11883
rect 11520 11840 11572 11849
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 18420 11840 18472 11892
rect 19340 11840 19392 11892
rect 8484 11772 8536 11824
rect 10416 11815 10468 11824
rect 10416 11781 10425 11815
rect 10425 11781 10459 11815
rect 10459 11781 10468 11815
rect 10416 11772 10468 11781
rect 11060 11772 11112 11824
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 2596 11747 2648 11756
rect 2596 11713 2605 11747
rect 2605 11713 2639 11747
rect 2639 11713 2648 11747
rect 2596 11704 2648 11713
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 10048 11704 10100 11756
rect 10876 11704 10928 11756
rect 18512 11772 18564 11824
rect 12808 11747 12860 11756
rect 12808 11713 12817 11747
rect 12817 11713 12851 11747
rect 12851 11713 12860 11747
rect 12808 11704 12860 11713
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 13176 11704 13228 11756
rect 13728 11704 13780 11756
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 17316 11747 17368 11756
rect 17316 11713 17325 11747
rect 17325 11713 17359 11747
rect 17359 11713 17368 11747
rect 17316 11704 17368 11713
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 20444 11704 20496 11756
rect 20720 11840 20772 11892
rect 20812 11840 20864 11892
rect 22836 11840 22888 11892
rect 23296 11840 23348 11892
rect 23480 11840 23532 11892
rect 27252 11883 27304 11892
rect 27252 11849 27261 11883
rect 27261 11849 27295 11883
rect 27295 11849 27304 11883
rect 27252 11840 27304 11849
rect 27712 11840 27764 11892
rect 28080 11840 28132 11892
rect 23756 11772 23808 11824
rect 24584 11772 24636 11824
rect 20812 11747 20864 11756
rect 7932 11636 7984 11688
rect 19156 11679 19208 11688
rect 19156 11645 19165 11679
rect 19165 11645 19199 11679
rect 19199 11645 19208 11679
rect 19156 11636 19208 11645
rect 19892 11636 19944 11688
rect 20812 11713 20821 11747
rect 20821 11713 20855 11747
rect 20855 11713 20864 11747
rect 20812 11704 20864 11713
rect 20904 11747 20956 11756
rect 20904 11713 20913 11747
rect 20913 11713 20947 11747
rect 20947 11713 20956 11747
rect 23020 11747 23072 11756
rect 20904 11704 20956 11713
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 23664 11704 23716 11756
rect 23848 11747 23900 11756
rect 23848 11713 23857 11747
rect 23857 11713 23891 11747
rect 23891 11713 23900 11747
rect 23848 11704 23900 11713
rect 24032 11747 24084 11756
rect 24032 11713 24041 11747
rect 24041 11713 24075 11747
rect 24075 11713 24084 11747
rect 24032 11704 24084 11713
rect 24676 11747 24728 11756
rect 24676 11713 24685 11747
rect 24685 11713 24719 11747
rect 24719 11713 24728 11747
rect 24676 11704 24728 11713
rect 24768 11747 24820 11756
rect 24768 11713 24777 11747
rect 24777 11713 24811 11747
rect 24811 11713 24820 11747
rect 24952 11747 25004 11756
rect 24768 11704 24820 11713
rect 24952 11713 24961 11747
rect 24961 11713 24995 11747
rect 24995 11713 25004 11747
rect 24952 11704 25004 11713
rect 23296 11636 23348 11688
rect 26700 11636 26752 11688
rect 27712 11679 27764 11688
rect 27712 11645 27721 11679
rect 27721 11645 27755 11679
rect 27755 11645 27764 11679
rect 27712 11636 27764 11645
rect 28264 11636 28316 11688
rect 13912 11568 13964 11620
rect 17592 11568 17644 11620
rect 19248 11611 19300 11620
rect 19248 11577 19257 11611
rect 19257 11577 19291 11611
rect 19291 11577 19300 11611
rect 19248 11568 19300 11577
rect 4252 11500 4304 11552
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 6736 11500 6788 11552
rect 10140 11500 10192 11552
rect 10968 11500 11020 11552
rect 11336 11500 11388 11552
rect 12808 11500 12860 11552
rect 13728 11543 13780 11552
rect 13728 11509 13737 11543
rect 13737 11509 13771 11543
rect 13771 11509 13780 11543
rect 13728 11500 13780 11509
rect 20076 11543 20128 11552
rect 20076 11509 20085 11543
rect 20085 11509 20119 11543
rect 20119 11509 20128 11543
rect 20076 11500 20128 11509
rect 23940 11543 23992 11552
rect 23940 11509 23949 11543
rect 23949 11509 23983 11543
rect 23983 11509 23992 11543
rect 23940 11500 23992 11509
rect 4492 11398 4544 11450
rect 4556 11398 4608 11450
rect 4620 11398 4672 11450
rect 4684 11398 4736 11450
rect 4748 11398 4800 11450
rect 11576 11398 11628 11450
rect 11640 11398 11692 11450
rect 11704 11398 11756 11450
rect 11768 11398 11820 11450
rect 11832 11398 11884 11450
rect 18660 11398 18712 11450
rect 18724 11398 18776 11450
rect 18788 11398 18840 11450
rect 18852 11398 18904 11450
rect 18916 11398 18968 11450
rect 25744 11398 25796 11450
rect 25808 11398 25860 11450
rect 25872 11398 25924 11450
rect 25936 11398 25988 11450
rect 26000 11398 26052 11450
rect 1768 11339 1820 11348
rect 1768 11305 1777 11339
rect 1777 11305 1811 11339
rect 1811 11305 1820 11339
rect 1768 11296 1820 11305
rect 17224 11339 17276 11348
rect 17224 11305 17233 11339
rect 17233 11305 17267 11339
rect 17267 11305 17276 11339
rect 17224 11296 17276 11305
rect 5632 11228 5684 11280
rect 9864 11228 9916 11280
rect 17776 11296 17828 11348
rect 18512 11296 18564 11348
rect 19156 11228 19208 11280
rect 19892 11296 19944 11348
rect 20076 11296 20128 11348
rect 23756 11296 23808 11348
rect 24768 11296 24820 11348
rect 27620 11339 27672 11348
rect 27620 11305 27629 11339
rect 27629 11305 27663 11339
rect 27663 11305 27672 11339
rect 27620 11296 27672 11305
rect 27804 11296 27856 11348
rect 23388 11228 23440 11280
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 4896 11160 4948 11212
rect 7840 11160 7892 11212
rect 9036 11203 9088 11212
rect 9036 11169 9045 11203
rect 9045 11169 9079 11203
rect 9079 11169 9088 11203
rect 9036 11160 9088 11169
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 4804 11092 4856 11144
rect 5172 11092 5224 11144
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8392 11092 8444 11144
rect 8668 11092 8720 11144
rect 3332 11024 3384 11076
rect 4712 11024 4764 11076
rect 5080 11024 5132 11076
rect 6736 11024 6788 11076
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 11336 11160 11388 11212
rect 12900 11203 12952 11212
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 13544 11160 13596 11212
rect 15016 11160 15068 11212
rect 18512 11160 18564 11212
rect 21272 11160 21324 11212
rect 27160 11160 27212 11212
rect 28172 11160 28224 11212
rect 9128 11092 9180 11101
rect 8852 11024 8904 11076
rect 10692 11092 10744 11144
rect 9772 11024 9824 11076
rect 10784 11024 10836 11076
rect 7656 10956 7708 11008
rect 12716 10999 12768 11008
rect 12716 10965 12725 10999
rect 12725 10965 12759 10999
rect 12759 10965 12768 10999
rect 12716 10956 12768 10965
rect 12900 11024 12952 11076
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 14188 11135 14240 11144
rect 13176 11092 13228 11101
rect 14188 11101 14197 11135
rect 14197 11101 14231 11135
rect 14231 11101 14240 11135
rect 14188 11092 14240 11101
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 14648 11092 14700 11144
rect 17132 11135 17184 11144
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 17132 11092 17184 11101
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 16580 11067 16632 11076
rect 16580 11033 16589 11067
rect 16589 11033 16623 11067
rect 16623 11033 16632 11067
rect 16580 11024 16632 11033
rect 19156 11092 19208 11144
rect 20076 11092 20128 11144
rect 25504 11092 25556 11144
rect 27344 11092 27396 11144
rect 12992 10956 13044 11008
rect 14648 10999 14700 11008
rect 14648 10965 14657 10999
rect 14657 10965 14691 10999
rect 14691 10965 14700 10999
rect 14648 10956 14700 10965
rect 19892 11024 19944 11076
rect 27804 11024 27856 11076
rect 19340 10956 19392 11008
rect 8034 10854 8086 10906
rect 8098 10854 8150 10906
rect 8162 10854 8214 10906
rect 8226 10854 8278 10906
rect 8290 10854 8342 10906
rect 15118 10854 15170 10906
rect 15182 10854 15234 10906
rect 15246 10854 15298 10906
rect 15310 10854 15362 10906
rect 15374 10854 15426 10906
rect 22202 10854 22254 10906
rect 22266 10854 22318 10906
rect 22330 10854 22382 10906
rect 22394 10854 22446 10906
rect 22458 10854 22510 10906
rect 29286 10854 29338 10906
rect 29350 10854 29402 10906
rect 29414 10854 29466 10906
rect 29478 10854 29530 10906
rect 29542 10854 29594 10906
rect 1492 10795 1544 10804
rect 1492 10761 1501 10795
rect 1501 10761 1535 10795
rect 1535 10761 1544 10795
rect 1492 10752 1544 10761
rect 5632 10795 5684 10804
rect 5632 10761 5657 10795
rect 5657 10761 5684 10795
rect 5632 10752 5684 10761
rect 6000 10752 6052 10804
rect 10876 10752 10928 10804
rect 14188 10752 14240 10804
rect 17408 10752 17460 10804
rect 18236 10795 18288 10804
rect 18236 10761 18245 10795
rect 18245 10761 18279 10795
rect 18279 10761 18288 10795
rect 18236 10752 18288 10761
rect 20628 10795 20680 10804
rect 20628 10761 20637 10795
rect 20637 10761 20671 10795
rect 20671 10761 20680 10795
rect 20628 10752 20680 10761
rect 20812 10752 20864 10804
rect 21548 10752 21600 10804
rect 23388 10752 23440 10804
rect 5448 10727 5500 10736
rect 5448 10693 5457 10727
rect 5457 10693 5491 10727
rect 5491 10693 5500 10727
rect 5448 10684 5500 10693
rect 7840 10684 7892 10736
rect 2228 10616 2280 10668
rect 4896 10616 4948 10668
rect 7932 10659 7984 10668
rect 7932 10625 7941 10659
rect 7941 10625 7975 10659
rect 7975 10625 7984 10659
rect 7932 10616 7984 10625
rect 17132 10684 17184 10736
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8668 10616 8720 10625
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 12900 10616 12952 10668
rect 13452 10659 13504 10668
rect 13452 10625 13461 10659
rect 13461 10625 13495 10659
rect 13495 10625 13504 10659
rect 13452 10616 13504 10625
rect 13636 10659 13688 10668
rect 13636 10625 13645 10659
rect 13645 10625 13679 10659
rect 13679 10625 13688 10659
rect 13636 10616 13688 10625
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 19248 10684 19300 10736
rect 4252 10548 4304 10600
rect 4712 10591 4764 10600
rect 4712 10557 4721 10591
rect 4721 10557 4755 10591
rect 4755 10557 4764 10591
rect 4712 10548 4764 10557
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 5356 10548 5408 10600
rect 9404 10523 9456 10532
rect 9404 10489 9413 10523
rect 9413 10489 9447 10523
rect 9447 10489 9456 10523
rect 9404 10480 9456 10489
rect 11980 10480 12032 10532
rect 19432 10616 19484 10668
rect 21272 10616 21324 10668
rect 21456 10616 21508 10668
rect 21916 10659 21968 10668
rect 21916 10625 21925 10659
rect 21925 10625 21959 10659
rect 21959 10625 21968 10659
rect 21916 10616 21968 10625
rect 22284 10616 22336 10668
rect 23020 10684 23072 10736
rect 22744 10659 22796 10668
rect 22744 10625 22753 10659
rect 22753 10625 22787 10659
rect 22787 10625 22796 10659
rect 22744 10616 22796 10625
rect 23296 10659 23348 10668
rect 23296 10625 23305 10659
rect 23305 10625 23339 10659
rect 23339 10625 23348 10659
rect 23296 10616 23348 10625
rect 23388 10616 23440 10668
rect 2136 10412 2188 10464
rect 3148 10412 3200 10464
rect 4896 10412 4948 10464
rect 12900 10412 12952 10464
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 13728 10455 13780 10464
rect 13728 10421 13737 10455
rect 13737 10421 13771 10455
rect 13771 10421 13780 10455
rect 13728 10412 13780 10421
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 20720 10591 20772 10600
rect 19984 10548 20036 10557
rect 20720 10557 20729 10591
rect 20729 10557 20763 10591
rect 20763 10557 20772 10591
rect 20720 10548 20772 10557
rect 25136 10752 25188 10804
rect 27712 10752 27764 10804
rect 23848 10616 23900 10668
rect 24860 10659 24912 10668
rect 20352 10480 20404 10532
rect 23296 10480 23348 10532
rect 24216 10523 24268 10532
rect 24216 10489 24225 10523
rect 24225 10489 24259 10523
rect 24259 10489 24268 10523
rect 24216 10480 24268 10489
rect 24860 10625 24869 10659
rect 24869 10625 24903 10659
rect 24903 10625 24912 10659
rect 24860 10616 24912 10625
rect 25320 10616 25372 10668
rect 28264 10684 28316 10736
rect 25688 10616 25740 10668
rect 27160 10659 27212 10668
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 25136 10591 25188 10600
rect 24860 10480 24912 10532
rect 25136 10557 25145 10591
rect 25145 10557 25179 10591
rect 25179 10557 25188 10591
rect 25136 10548 25188 10557
rect 27804 10616 27856 10668
rect 25596 10480 25648 10532
rect 28172 10480 28224 10532
rect 20812 10412 20864 10464
rect 20904 10412 20956 10464
rect 22560 10455 22612 10464
rect 22560 10421 22569 10455
rect 22569 10421 22603 10455
rect 22603 10421 22612 10455
rect 22560 10412 22612 10421
rect 22744 10412 22796 10464
rect 25688 10412 25740 10464
rect 27804 10455 27856 10464
rect 27804 10421 27813 10455
rect 27813 10421 27847 10455
rect 27847 10421 27856 10455
rect 27804 10412 27856 10421
rect 4492 10310 4544 10362
rect 4556 10310 4608 10362
rect 4620 10310 4672 10362
rect 4684 10310 4736 10362
rect 4748 10310 4800 10362
rect 11576 10310 11628 10362
rect 11640 10310 11692 10362
rect 11704 10310 11756 10362
rect 11768 10310 11820 10362
rect 11832 10310 11884 10362
rect 18660 10310 18712 10362
rect 18724 10310 18776 10362
rect 18788 10310 18840 10362
rect 18852 10310 18904 10362
rect 18916 10310 18968 10362
rect 25744 10310 25796 10362
rect 25808 10310 25860 10362
rect 25872 10310 25924 10362
rect 25936 10310 25988 10362
rect 26000 10310 26052 10362
rect 9496 10208 9548 10260
rect 12716 10208 12768 10260
rect 13176 10208 13228 10260
rect 17316 10208 17368 10260
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 20720 10208 20772 10260
rect 13728 10140 13780 10192
rect 7656 10115 7708 10124
rect 7656 10081 7665 10115
rect 7665 10081 7699 10115
rect 7699 10081 7708 10115
rect 7656 10072 7708 10081
rect 13820 10072 13872 10124
rect 4160 10004 4212 10056
rect 8392 10004 8444 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 12348 10047 12400 10056
rect 12348 10013 12357 10047
rect 12357 10013 12391 10047
rect 12391 10013 12400 10047
rect 12348 10004 12400 10013
rect 12440 10047 12492 10056
rect 12440 10013 12450 10047
rect 12450 10013 12484 10047
rect 12484 10013 12492 10047
rect 12440 10004 12492 10013
rect 12992 10004 13044 10056
rect 15752 10004 15804 10056
rect 16764 10004 16816 10056
rect 12256 9936 12308 9988
rect 2412 9868 2464 9920
rect 7932 9911 7984 9920
rect 7932 9877 7941 9911
rect 7941 9877 7975 9911
rect 7975 9877 7984 9911
rect 7932 9868 7984 9877
rect 13084 9936 13136 9988
rect 13544 9936 13596 9988
rect 19340 10047 19392 10056
rect 19340 10013 19349 10047
rect 19349 10013 19383 10047
rect 19383 10013 19392 10047
rect 19340 10004 19392 10013
rect 20628 10004 20680 10056
rect 20720 9979 20772 9988
rect 20720 9945 20729 9979
rect 20729 9945 20763 9979
rect 20763 9945 20772 9979
rect 20720 9936 20772 9945
rect 21916 10208 21968 10260
rect 22284 10251 22336 10260
rect 22284 10217 22293 10251
rect 22293 10217 22327 10251
rect 22327 10217 22336 10251
rect 22284 10208 22336 10217
rect 23388 10208 23440 10260
rect 25136 10208 25188 10260
rect 22744 10072 22796 10124
rect 23112 10072 23164 10124
rect 21640 10047 21692 10056
rect 21640 10013 21649 10047
rect 21649 10013 21683 10047
rect 21683 10013 21692 10047
rect 21640 10004 21692 10013
rect 25320 10072 25372 10124
rect 25596 10072 25648 10124
rect 28172 10115 28224 10124
rect 28172 10081 28181 10115
rect 28181 10081 28215 10115
rect 28215 10081 28224 10115
rect 28172 10072 28224 10081
rect 28264 10115 28316 10124
rect 28264 10081 28273 10115
rect 28273 10081 28307 10115
rect 28307 10081 28316 10115
rect 28264 10072 28316 10081
rect 20904 9936 20956 9988
rect 22192 9936 22244 9988
rect 13912 9868 13964 9920
rect 16764 9868 16816 9920
rect 17776 9911 17828 9920
rect 17776 9877 17785 9911
rect 17785 9877 17819 9911
rect 17819 9877 17828 9911
rect 17776 9868 17828 9877
rect 18696 9911 18748 9920
rect 18696 9877 18705 9911
rect 18705 9877 18739 9911
rect 18739 9877 18748 9911
rect 18696 9868 18748 9877
rect 19432 9868 19484 9920
rect 25504 10047 25556 10056
rect 22744 9936 22796 9988
rect 23296 9936 23348 9988
rect 25504 10013 25513 10047
rect 25513 10013 25547 10047
rect 25547 10013 25556 10047
rect 25504 10004 25556 10013
rect 26884 10047 26936 10056
rect 26884 10013 26893 10047
rect 26893 10013 26927 10047
rect 26927 10013 26936 10047
rect 26884 10004 26936 10013
rect 27712 10004 27764 10056
rect 27620 9936 27672 9988
rect 22928 9868 22980 9920
rect 25412 9868 25464 9920
rect 26516 9911 26568 9920
rect 26516 9877 26525 9911
rect 26525 9877 26559 9911
rect 26559 9877 26568 9911
rect 26516 9868 26568 9877
rect 8034 9766 8086 9818
rect 8098 9766 8150 9818
rect 8162 9766 8214 9818
rect 8226 9766 8278 9818
rect 8290 9766 8342 9818
rect 15118 9766 15170 9818
rect 15182 9766 15234 9818
rect 15246 9766 15298 9818
rect 15310 9766 15362 9818
rect 15374 9766 15426 9818
rect 22202 9766 22254 9818
rect 22266 9766 22318 9818
rect 22330 9766 22382 9818
rect 22394 9766 22446 9818
rect 22458 9766 22510 9818
rect 29286 9766 29338 9818
rect 29350 9766 29402 9818
rect 29414 9766 29466 9818
rect 29478 9766 29530 9818
rect 29542 9766 29594 9818
rect 2228 9596 2280 9648
rect 3148 9639 3200 9648
rect 3148 9605 3157 9639
rect 3157 9605 3191 9639
rect 3191 9605 3200 9639
rect 3148 9596 3200 9605
rect 3884 9596 3936 9648
rect 7288 9639 7340 9648
rect 7288 9605 7297 9639
rect 7297 9605 7331 9639
rect 7331 9605 7340 9639
rect 7288 9596 7340 9605
rect 8300 9596 8352 9648
rect 8576 9596 8628 9648
rect 2412 9528 2464 9580
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 4344 9571 4396 9580
rect 3332 9528 3384 9537
rect 4344 9537 4353 9571
rect 4353 9537 4387 9571
rect 4387 9537 4396 9571
rect 4344 9528 4396 9537
rect 7012 9528 7064 9580
rect 7932 9571 7984 9580
rect 7932 9537 7941 9571
rect 7941 9537 7975 9571
rect 7975 9537 7984 9571
rect 7932 9528 7984 9537
rect 8392 9528 8444 9580
rect 9220 9596 9272 9648
rect 9680 9596 9732 9648
rect 10508 9664 10560 9716
rect 12348 9707 12400 9716
rect 12348 9673 12357 9707
rect 12357 9673 12391 9707
rect 12391 9673 12400 9707
rect 12348 9664 12400 9673
rect 17408 9707 17460 9716
rect 17408 9673 17417 9707
rect 17417 9673 17451 9707
rect 17451 9673 17460 9707
rect 17408 9664 17460 9673
rect 20720 9664 20772 9716
rect 22468 9664 22520 9716
rect 22928 9707 22980 9716
rect 22928 9673 22937 9707
rect 22937 9673 22971 9707
rect 22971 9673 22980 9707
rect 22928 9664 22980 9673
rect 27804 9707 27856 9716
rect 27804 9673 27813 9707
rect 27813 9673 27847 9707
rect 27847 9673 27856 9707
rect 27804 9664 27856 9673
rect 10968 9528 11020 9580
rect 13728 9596 13780 9648
rect 12808 9528 12860 9580
rect 14096 9528 14148 9580
rect 14924 9528 14976 9580
rect 17592 9596 17644 9648
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 17040 9528 17092 9580
rect 18696 9639 18748 9648
rect 7932 9392 7984 9444
rect 11060 9460 11112 9512
rect 12256 9460 12308 9512
rect 12532 9460 12584 9512
rect 13084 9460 13136 9512
rect 13912 9460 13964 9512
rect 14556 9460 14608 9512
rect 18696 9605 18705 9639
rect 18705 9605 18739 9639
rect 18739 9605 18748 9639
rect 18696 9596 18748 9605
rect 19616 9596 19668 9648
rect 23296 9596 23348 9648
rect 24952 9639 25004 9648
rect 24952 9605 24961 9639
rect 24961 9605 24995 9639
rect 24995 9605 25004 9639
rect 24952 9596 25004 9605
rect 25136 9596 25188 9648
rect 20812 9528 20864 9580
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 22468 9528 22520 9580
rect 23848 9571 23900 9580
rect 23848 9537 23857 9571
rect 23857 9537 23891 9571
rect 23891 9537 23900 9571
rect 23848 9528 23900 9537
rect 25228 9571 25280 9580
rect 25228 9537 25237 9571
rect 25237 9537 25271 9571
rect 25271 9537 25280 9571
rect 25228 9528 25280 9537
rect 25412 9571 25464 9580
rect 25412 9537 25421 9571
rect 25421 9537 25455 9571
rect 25455 9537 25464 9571
rect 25596 9571 25648 9580
rect 25412 9528 25464 9537
rect 25596 9537 25605 9571
rect 25605 9537 25639 9571
rect 25639 9537 25648 9571
rect 25596 9528 25648 9537
rect 14648 9392 14700 9444
rect 2504 9367 2556 9376
rect 2504 9333 2513 9367
rect 2513 9333 2547 9367
rect 2547 9333 2556 9367
rect 2504 9324 2556 9333
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 4344 9324 4396 9376
rect 7564 9324 7616 9376
rect 10968 9324 11020 9376
rect 12532 9367 12584 9376
rect 12532 9333 12541 9367
rect 12541 9333 12575 9367
rect 12575 9333 12584 9367
rect 12532 9324 12584 9333
rect 12624 9324 12676 9376
rect 14188 9324 14240 9376
rect 14924 9324 14976 9376
rect 17040 9324 17092 9376
rect 23480 9503 23532 9512
rect 23480 9469 23489 9503
rect 23489 9469 23523 9503
rect 23523 9469 23532 9503
rect 28724 9571 28776 9580
rect 28724 9537 28733 9571
rect 28733 9537 28767 9571
rect 28767 9537 28776 9571
rect 28724 9528 28776 9537
rect 23480 9460 23532 9469
rect 28080 9460 28132 9512
rect 20628 9324 20680 9376
rect 20904 9324 20956 9376
rect 27620 9392 27672 9444
rect 22744 9324 22796 9376
rect 22928 9324 22980 9376
rect 23664 9324 23716 9376
rect 28816 9392 28868 9444
rect 28540 9367 28592 9376
rect 28540 9333 28549 9367
rect 28549 9333 28583 9367
rect 28583 9333 28592 9367
rect 28540 9324 28592 9333
rect 4492 9222 4544 9274
rect 4556 9222 4608 9274
rect 4620 9222 4672 9274
rect 4684 9222 4736 9274
rect 4748 9222 4800 9274
rect 11576 9222 11628 9274
rect 11640 9222 11692 9274
rect 11704 9222 11756 9274
rect 11768 9222 11820 9274
rect 11832 9222 11884 9274
rect 18660 9222 18712 9274
rect 18724 9222 18776 9274
rect 18788 9222 18840 9274
rect 18852 9222 18904 9274
rect 18916 9222 18968 9274
rect 25744 9222 25796 9274
rect 25808 9222 25860 9274
rect 25872 9222 25924 9274
rect 25936 9222 25988 9274
rect 26000 9222 26052 9274
rect 2320 9120 2372 9172
rect 3884 9163 3936 9172
rect 3884 9129 3893 9163
rect 3893 9129 3927 9163
rect 3927 9129 3936 9163
rect 3884 9120 3936 9129
rect 5080 9120 5132 9172
rect 7012 9163 7064 9172
rect 7012 9129 7021 9163
rect 7021 9129 7055 9163
rect 7055 9129 7064 9163
rect 7012 9120 7064 9129
rect 8300 9163 8352 9172
rect 8300 9129 8309 9163
rect 8309 9129 8343 9163
rect 8343 9129 8352 9163
rect 8300 9120 8352 9129
rect 8760 9120 8812 9172
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 10784 9120 10836 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 8576 9052 8628 9104
rect 14096 9052 14148 9104
rect 2780 8984 2832 9036
rect 4896 9027 4948 9036
rect 4896 8993 4905 9027
rect 4905 8993 4939 9027
rect 4939 8993 4948 9027
rect 4896 8984 4948 8993
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 4344 8916 4396 8968
rect 4804 8916 4856 8968
rect 5632 8916 5684 8968
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 8300 8984 8352 9036
rect 4620 8823 4672 8832
rect 4620 8789 4629 8823
rect 4629 8789 4663 8823
rect 4663 8789 4672 8823
rect 4620 8780 4672 8789
rect 5448 8848 5500 8900
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 9036 8916 9088 8968
rect 13452 8984 13504 9036
rect 13820 8984 13872 9036
rect 23296 9120 23348 9172
rect 24860 9120 24912 9172
rect 27620 9120 27672 9172
rect 28080 9120 28132 9172
rect 28356 9120 28408 9172
rect 28724 9163 28776 9172
rect 28724 9129 28733 9163
rect 28733 9129 28767 9163
rect 28767 9129 28776 9163
rect 28724 9120 28776 9129
rect 14464 9052 14516 9104
rect 20628 9052 20680 9104
rect 28172 9052 28224 9104
rect 28540 9052 28592 9104
rect 9588 8916 9640 8968
rect 14464 8916 14516 8968
rect 14832 8984 14884 9036
rect 4988 8780 5040 8832
rect 6552 8780 6604 8832
rect 13636 8848 13688 8900
rect 13728 8848 13780 8900
rect 15108 8984 15160 9036
rect 17776 8984 17828 9036
rect 23848 8984 23900 9036
rect 25596 9027 25648 9036
rect 25596 8993 25605 9027
rect 25605 8993 25639 9027
rect 25639 8993 25648 9027
rect 25596 8984 25648 8993
rect 8300 8780 8352 8832
rect 8484 8780 8536 8832
rect 9588 8780 9640 8832
rect 12624 8780 12676 8832
rect 12900 8780 12952 8832
rect 16028 8916 16080 8968
rect 17592 8916 17644 8968
rect 26424 8916 26476 8968
rect 25228 8848 25280 8900
rect 15476 8780 15528 8832
rect 17592 8780 17644 8832
rect 23848 8780 23900 8832
rect 24216 8780 24268 8832
rect 25412 8823 25464 8832
rect 25412 8789 25421 8823
rect 25421 8789 25455 8823
rect 25455 8789 25464 8823
rect 25412 8780 25464 8789
rect 8034 8678 8086 8730
rect 8098 8678 8150 8730
rect 8162 8678 8214 8730
rect 8226 8678 8278 8730
rect 8290 8678 8342 8730
rect 15118 8678 15170 8730
rect 15182 8678 15234 8730
rect 15246 8678 15298 8730
rect 15310 8678 15362 8730
rect 15374 8678 15426 8730
rect 22202 8678 22254 8730
rect 22266 8678 22318 8730
rect 22330 8678 22382 8730
rect 22394 8678 22446 8730
rect 22458 8678 22510 8730
rect 29286 8678 29338 8730
rect 29350 8678 29402 8730
rect 29414 8678 29466 8730
rect 29478 8678 29530 8730
rect 29542 8678 29594 8730
rect 4988 8576 5040 8628
rect 5448 8576 5500 8628
rect 7196 8576 7248 8628
rect 1584 8551 1636 8560
rect 1584 8517 1593 8551
rect 1593 8517 1627 8551
rect 1627 8517 1636 8551
rect 1584 8508 1636 8517
rect 2320 8440 2372 8492
rect 4160 8508 4212 8560
rect 4896 8508 4948 8560
rect 5724 8551 5776 8560
rect 5724 8517 5733 8551
rect 5733 8517 5767 8551
rect 5767 8517 5776 8551
rect 5724 8508 5776 8517
rect 6552 8508 6604 8560
rect 7932 8508 7984 8560
rect 8760 8576 8812 8628
rect 9772 8508 9824 8560
rect 11060 8576 11112 8628
rect 14832 8576 14884 8628
rect 15476 8576 15528 8628
rect 17224 8576 17276 8628
rect 12256 8508 12308 8560
rect 14924 8551 14976 8560
rect 14924 8517 14933 8551
rect 14933 8517 14967 8551
rect 14967 8517 14976 8551
rect 14924 8508 14976 8517
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 8944 8440 8996 8492
rect 13912 8440 13964 8492
rect 14096 8440 14148 8492
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 16672 8508 16724 8560
rect 20076 8551 20128 8560
rect 14740 8440 14792 8449
rect 15476 8483 15528 8492
rect 15476 8449 15485 8483
rect 15485 8449 15519 8483
rect 15519 8449 15528 8483
rect 15660 8483 15712 8492
rect 15476 8440 15528 8449
rect 15660 8449 15669 8483
rect 15669 8449 15703 8483
rect 15703 8449 15712 8483
rect 15660 8440 15712 8449
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 20076 8517 20085 8551
rect 20085 8517 20119 8551
rect 20119 8517 20128 8551
rect 20076 8508 20128 8517
rect 22100 8576 22152 8628
rect 22376 8576 22428 8628
rect 23020 8619 23072 8628
rect 23020 8585 23029 8619
rect 23029 8585 23063 8619
rect 23063 8585 23072 8619
rect 23020 8576 23072 8585
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 25228 8619 25280 8628
rect 25228 8585 25237 8619
rect 25237 8585 25271 8619
rect 25271 8585 25280 8619
rect 25228 8576 25280 8585
rect 25412 8576 25464 8628
rect 27436 8576 27488 8628
rect 17592 8483 17644 8492
rect 1860 8372 1912 8424
rect 4804 8415 4856 8424
rect 4804 8381 4813 8415
rect 4813 8381 4847 8415
rect 4847 8381 4856 8415
rect 4804 8372 4856 8381
rect 5264 8372 5316 8424
rect 5632 8372 5684 8424
rect 8576 8372 8628 8424
rect 13084 8415 13136 8424
rect 13084 8381 13093 8415
rect 13093 8381 13127 8415
rect 13127 8381 13136 8415
rect 13084 8372 13136 8381
rect 13636 8372 13688 8424
rect 17592 8449 17601 8483
rect 17601 8449 17635 8483
rect 17635 8449 17644 8483
rect 17592 8440 17644 8449
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 22652 8508 22704 8560
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 20996 8440 21048 8492
rect 22100 8440 22152 8492
rect 25596 8440 25648 8492
rect 22560 8372 22612 8424
rect 27436 8415 27488 8424
rect 1860 8279 1912 8288
rect 1860 8245 1869 8279
rect 1869 8245 1903 8279
rect 1903 8245 1912 8279
rect 1860 8236 1912 8245
rect 1952 8236 2004 8288
rect 2780 8279 2832 8288
rect 2780 8245 2789 8279
rect 2789 8245 2823 8279
rect 2823 8245 2832 8279
rect 3424 8279 3476 8288
rect 2780 8236 2832 8245
rect 3424 8245 3433 8279
rect 3433 8245 3467 8279
rect 3467 8245 3476 8279
rect 3424 8236 3476 8245
rect 4620 8236 4672 8288
rect 5264 8236 5316 8288
rect 10692 8236 10744 8288
rect 15016 8236 15068 8288
rect 15568 8304 15620 8356
rect 17316 8304 17368 8356
rect 25596 8304 25648 8356
rect 27436 8381 27445 8415
rect 27445 8381 27479 8415
rect 27479 8381 27488 8415
rect 27436 8372 27488 8381
rect 27528 8415 27580 8424
rect 27528 8381 27537 8415
rect 27537 8381 27571 8415
rect 27571 8381 27580 8415
rect 27528 8372 27580 8381
rect 16764 8236 16816 8288
rect 16948 8279 17000 8288
rect 16948 8245 16957 8279
rect 16957 8245 16991 8279
rect 16991 8245 17000 8279
rect 16948 8236 17000 8245
rect 22468 8236 22520 8288
rect 22836 8236 22888 8288
rect 4492 8134 4544 8186
rect 4556 8134 4608 8186
rect 4620 8134 4672 8186
rect 4684 8134 4736 8186
rect 4748 8134 4800 8186
rect 11576 8134 11628 8186
rect 11640 8134 11692 8186
rect 11704 8134 11756 8186
rect 11768 8134 11820 8186
rect 11832 8134 11884 8186
rect 18660 8134 18712 8186
rect 18724 8134 18776 8186
rect 18788 8134 18840 8186
rect 18852 8134 18904 8186
rect 18916 8134 18968 8186
rect 25744 8134 25796 8186
rect 25808 8134 25860 8186
rect 25872 8134 25924 8186
rect 25936 8134 25988 8186
rect 26000 8134 26052 8186
rect 1584 8032 1636 8084
rect 2964 8032 3016 8084
rect 6184 8032 6236 8084
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 12440 8032 12492 8084
rect 13084 8032 13136 8084
rect 2504 7896 2556 7948
rect 4988 7964 5040 8016
rect 5172 7964 5224 8016
rect 5356 7964 5408 8016
rect 5724 7896 5776 7948
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 9864 7896 9916 7948
rect 14096 8007 14148 8016
rect 14096 7973 14105 8007
rect 14105 7973 14139 8007
rect 14139 7973 14148 8007
rect 14096 7964 14148 7973
rect 14464 7964 14516 8016
rect 14832 7964 14884 8016
rect 15660 8032 15712 8084
rect 15752 8032 15804 8084
rect 19616 8032 19668 8084
rect 20996 8075 21048 8084
rect 10876 7871 10928 7880
rect 7932 7760 7984 7812
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 11152 7760 11204 7812
rect 2044 7735 2096 7744
rect 2044 7701 2053 7735
rect 2053 7701 2087 7735
rect 2087 7701 2096 7735
rect 2044 7692 2096 7701
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 5080 7692 5132 7744
rect 10140 7735 10192 7744
rect 10140 7701 10149 7735
rect 10149 7701 10183 7735
rect 10183 7701 10192 7735
rect 10140 7692 10192 7701
rect 10324 7692 10376 7744
rect 15476 7828 15528 7880
rect 15660 7871 15712 7880
rect 15660 7837 15664 7871
rect 15664 7837 15698 7871
rect 15698 7837 15712 7871
rect 15660 7828 15712 7837
rect 13912 7760 13964 7812
rect 15936 7871 15988 7880
rect 19984 7896 20036 7948
rect 20996 8041 21005 8075
rect 21005 8041 21039 8075
rect 21039 8041 21048 8075
rect 20996 8032 21048 8041
rect 22468 8075 22520 8084
rect 22468 8041 22477 8075
rect 22477 8041 22511 8075
rect 22511 8041 22520 8075
rect 22468 8032 22520 8041
rect 25596 8032 25648 8084
rect 26148 8032 26200 8084
rect 27528 7964 27580 8016
rect 15936 7837 15981 7871
rect 15981 7837 15988 7871
rect 15936 7828 15988 7837
rect 19432 7871 19484 7880
rect 15844 7803 15896 7812
rect 15844 7769 15853 7803
rect 15853 7769 15887 7803
rect 15887 7769 15896 7803
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 23664 7896 23716 7948
rect 15844 7760 15896 7769
rect 20352 7760 20404 7812
rect 21916 7760 21968 7812
rect 12992 7735 13044 7744
rect 12992 7701 13001 7735
rect 13001 7701 13035 7735
rect 13035 7701 13044 7735
rect 12992 7692 13044 7701
rect 14280 7692 14332 7744
rect 15752 7692 15804 7744
rect 16028 7692 16080 7744
rect 18236 7692 18288 7744
rect 19432 7692 19484 7744
rect 19984 7735 20036 7744
rect 19984 7701 19993 7735
rect 19993 7701 20027 7735
rect 20027 7701 20036 7735
rect 19984 7692 20036 7701
rect 21180 7735 21232 7744
rect 21180 7701 21189 7735
rect 21189 7701 21223 7735
rect 21223 7701 21232 7735
rect 21180 7692 21232 7701
rect 22652 7828 22704 7880
rect 23848 7828 23900 7880
rect 27436 7828 27488 7880
rect 27712 7760 27764 7812
rect 28448 7803 28500 7812
rect 28448 7769 28457 7803
rect 28457 7769 28491 7803
rect 28491 7769 28500 7803
rect 28448 7760 28500 7769
rect 28724 7760 28776 7812
rect 22744 7692 22796 7744
rect 23756 7692 23808 7744
rect 25964 7692 26016 7744
rect 8034 7590 8086 7642
rect 8098 7590 8150 7642
rect 8162 7590 8214 7642
rect 8226 7590 8278 7642
rect 8290 7590 8342 7642
rect 15118 7590 15170 7642
rect 15182 7590 15234 7642
rect 15246 7590 15298 7642
rect 15310 7590 15362 7642
rect 15374 7590 15426 7642
rect 22202 7590 22254 7642
rect 22266 7590 22318 7642
rect 22330 7590 22382 7642
rect 22394 7590 22446 7642
rect 22458 7590 22510 7642
rect 29286 7590 29338 7642
rect 29350 7590 29402 7642
rect 29414 7590 29466 7642
rect 29478 7590 29530 7642
rect 29542 7590 29594 7642
rect 5356 7531 5408 7540
rect 5356 7497 5365 7531
rect 5365 7497 5399 7531
rect 5399 7497 5408 7531
rect 5356 7488 5408 7497
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 8852 7488 8904 7540
rect 9128 7488 9180 7540
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 4620 7284 4672 7336
rect 5080 7327 5132 7336
rect 5080 7293 5089 7327
rect 5089 7293 5123 7327
rect 5123 7293 5132 7327
rect 5080 7284 5132 7293
rect 5172 7327 5224 7336
rect 5172 7293 5181 7327
rect 5181 7293 5215 7327
rect 5215 7293 5224 7327
rect 5172 7284 5224 7293
rect 7196 7284 7248 7336
rect 8760 7395 8812 7404
rect 8760 7361 8769 7395
rect 8769 7361 8803 7395
rect 8803 7361 8812 7395
rect 8760 7352 8812 7361
rect 9220 7352 9272 7404
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 11060 7488 11112 7540
rect 11336 7488 11388 7540
rect 12532 7488 12584 7540
rect 10692 7463 10744 7472
rect 10692 7429 10701 7463
rect 10701 7429 10735 7463
rect 10735 7429 10744 7463
rect 10692 7420 10744 7429
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 4988 7216 5040 7268
rect 9404 7284 9456 7336
rect 9772 7284 9824 7336
rect 10968 7352 11020 7404
rect 12992 7420 13044 7472
rect 9312 7216 9364 7268
rect 10876 7216 10928 7268
rect 12716 7395 12768 7404
rect 12716 7361 12761 7395
rect 12761 7361 12768 7395
rect 12716 7352 12768 7361
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 14188 7463 14240 7472
rect 14188 7429 14197 7463
rect 14197 7429 14231 7463
rect 14231 7429 14240 7463
rect 14188 7420 14240 7429
rect 14372 7463 14424 7472
rect 14372 7429 14397 7463
rect 14397 7429 14424 7463
rect 14648 7488 14700 7540
rect 17868 7488 17920 7540
rect 14372 7420 14424 7429
rect 14740 7420 14792 7472
rect 19524 7488 19576 7540
rect 20076 7488 20128 7540
rect 21916 7531 21968 7540
rect 21916 7497 21925 7531
rect 21925 7497 21959 7531
rect 21959 7497 21968 7531
rect 21916 7488 21968 7497
rect 25136 7488 25188 7540
rect 25964 7531 26016 7540
rect 25964 7497 25973 7531
rect 25973 7497 26007 7531
rect 26007 7497 26016 7531
rect 25964 7488 26016 7497
rect 27436 7488 27488 7540
rect 27712 7531 27764 7540
rect 27712 7497 27721 7531
rect 27721 7497 27755 7531
rect 27755 7497 27764 7531
rect 27712 7488 27764 7497
rect 16948 7395 17000 7404
rect 12900 7352 12952 7361
rect 13176 7284 13228 7336
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 17224 7395 17276 7404
rect 17224 7361 17233 7395
rect 17233 7361 17267 7395
rect 17267 7361 17276 7395
rect 17224 7352 17276 7361
rect 17776 7395 17828 7404
rect 17776 7361 17785 7395
rect 17785 7361 17819 7395
rect 17819 7361 17828 7395
rect 17776 7352 17828 7361
rect 20444 7420 20496 7472
rect 18604 7352 18656 7404
rect 19432 7352 19484 7404
rect 19616 7395 19668 7404
rect 19616 7361 19620 7395
rect 19620 7361 19654 7395
rect 19654 7361 19668 7395
rect 19616 7352 19668 7361
rect 17132 7284 17184 7336
rect 20352 7352 20404 7404
rect 22100 7420 22152 7472
rect 28724 7463 28776 7472
rect 28724 7429 28733 7463
rect 28733 7429 28767 7463
rect 28767 7429 28776 7463
rect 28724 7420 28776 7429
rect 22836 7395 22888 7404
rect 22836 7361 22845 7395
rect 22845 7361 22879 7395
rect 22879 7361 22888 7395
rect 22836 7352 22888 7361
rect 12624 7216 12676 7268
rect 1860 7148 1912 7200
rect 10140 7148 10192 7200
rect 10692 7148 10744 7200
rect 11244 7148 11296 7200
rect 11336 7148 11388 7200
rect 12348 7148 12400 7200
rect 15936 7216 15988 7268
rect 22652 7284 22704 7336
rect 23204 7284 23256 7336
rect 20812 7216 20864 7268
rect 23572 7395 23624 7404
rect 23572 7361 23581 7395
rect 23581 7361 23615 7395
rect 23615 7361 23624 7395
rect 23572 7352 23624 7361
rect 25504 7352 25556 7404
rect 27160 7284 27212 7336
rect 14096 7148 14148 7200
rect 15752 7148 15804 7200
rect 17040 7148 17092 7200
rect 19340 7148 19392 7200
rect 21180 7148 21232 7200
rect 21824 7148 21876 7200
rect 25596 7148 25648 7200
rect 27068 7191 27120 7200
rect 27068 7157 27077 7191
rect 27077 7157 27111 7191
rect 27111 7157 27120 7191
rect 27068 7148 27120 7157
rect 27896 7191 27948 7200
rect 27896 7157 27905 7191
rect 27905 7157 27939 7191
rect 27939 7157 27948 7191
rect 27896 7148 27948 7157
rect 4492 7046 4544 7098
rect 4556 7046 4608 7098
rect 4620 7046 4672 7098
rect 4684 7046 4736 7098
rect 4748 7046 4800 7098
rect 11576 7046 11628 7098
rect 11640 7046 11692 7098
rect 11704 7046 11756 7098
rect 11768 7046 11820 7098
rect 11832 7046 11884 7098
rect 18660 7046 18712 7098
rect 18724 7046 18776 7098
rect 18788 7046 18840 7098
rect 18852 7046 18904 7098
rect 18916 7046 18968 7098
rect 25744 7046 25796 7098
rect 25808 7046 25860 7098
rect 25872 7046 25924 7098
rect 25936 7046 25988 7098
rect 26000 7046 26052 7098
rect 4896 6987 4948 6996
rect 4896 6953 4905 6987
rect 4905 6953 4939 6987
rect 4939 6953 4948 6987
rect 4896 6944 4948 6953
rect 9220 6944 9272 6996
rect 9588 6944 9640 6996
rect 11428 6944 11480 6996
rect 12900 6944 12952 6996
rect 13912 6944 13964 6996
rect 9404 6919 9456 6928
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 4896 6740 4948 6792
rect 9404 6885 9413 6919
rect 9413 6885 9447 6919
rect 9447 6885 9456 6919
rect 9404 6876 9456 6885
rect 8392 6808 8444 6860
rect 9772 6876 9824 6928
rect 10600 6876 10652 6928
rect 14372 6944 14424 6996
rect 17224 6944 17276 6996
rect 18512 6944 18564 6996
rect 21180 6944 21232 6996
rect 5264 6740 5316 6792
rect 5908 6740 5960 6792
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 7196 6783 7248 6792
rect 7196 6749 7205 6783
rect 7205 6749 7239 6783
rect 7239 6749 7248 6783
rect 7196 6740 7248 6749
rect 9220 6740 9272 6792
rect 9680 6740 9732 6792
rect 8484 6672 8536 6724
rect 9864 6672 9916 6724
rect 10508 6740 10560 6792
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 11244 6783 11296 6792
rect 10784 6740 10836 6749
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 13268 6740 13320 6792
rect 14280 6808 14332 6860
rect 15844 6876 15896 6928
rect 17776 6876 17828 6928
rect 14188 6783 14240 6792
rect 14188 6749 14197 6783
rect 14197 6749 14231 6783
rect 14231 6749 14240 6783
rect 14188 6740 14240 6749
rect 15660 6740 15712 6792
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 5356 6604 5408 6656
rect 6184 6647 6236 6656
rect 6184 6613 6193 6647
rect 6193 6613 6227 6647
rect 6227 6613 6236 6647
rect 6184 6604 6236 6613
rect 9404 6604 9456 6656
rect 13820 6672 13872 6724
rect 17500 6808 17552 6860
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 18236 6783 18288 6792
rect 16764 6740 16816 6749
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 18512 6808 18564 6860
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 19524 6808 19576 6860
rect 20720 6851 20772 6860
rect 20720 6817 20729 6851
rect 20729 6817 20763 6851
rect 20763 6817 20772 6851
rect 20720 6808 20772 6817
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 19340 6783 19392 6792
rect 19340 6749 19350 6783
rect 19350 6749 19384 6783
rect 19384 6749 19392 6783
rect 19616 6783 19668 6792
rect 19340 6740 19392 6749
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 20444 6783 20496 6792
rect 17960 6672 18012 6724
rect 10140 6647 10192 6656
rect 10140 6613 10149 6647
rect 10149 6613 10183 6647
rect 10183 6613 10192 6647
rect 10140 6604 10192 6613
rect 12348 6604 12400 6656
rect 14740 6604 14792 6656
rect 17500 6647 17552 6656
rect 17500 6613 17509 6647
rect 17509 6613 17543 6647
rect 17543 6613 17552 6647
rect 17500 6604 17552 6613
rect 19524 6715 19576 6724
rect 19524 6681 19533 6715
rect 19533 6681 19567 6715
rect 19567 6681 19576 6715
rect 19524 6672 19576 6681
rect 20444 6749 20453 6783
rect 20453 6749 20487 6783
rect 20487 6749 20496 6783
rect 20444 6740 20496 6749
rect 20536 6783 20588 6792
rect 20536 6749 20545 6783
rect 20545 6749 20579 6783
rect 20579 6749 20588 6783
rect 20536 6740 20588 6749
rect 20904 6740 20956 6792
rect 22008 6783 22060 6792
rect 22008 6749 22017 6783
rect 22017 6749 22051 6783
rect 22051 6749 22060 6783
rect 22008 6740 22060 6749
rect 22744 6740 22796 6792
rect 23572 6944 23624 6996
rect 25596 6944 25648 6996
rect 27068 6944 27120 6996
rect 27896 6944 27948 6996
rect 27528 6808 27580 6860
rect 27620 6808 27672 6860
rect 28080 6808 28132 6860
rect 28356 6851 28408 6860
rect 28356 6817 28365 6851
rect 28365 6817 28399 6851
rect 28399 6817 28408 6851
rect 28356 6808 28408 6817
rect 21272 6672 21324 6724
rect 21364 6672 21416 6724
rect 28448 6740 28500 6792
rect 23664 6715 23716 6724
rect 23664 6681 23673 6715
rect 23673 6681 23707 6715
rect 23707 6681 23716 6715
rect 23664 6672 23716 6681
rect 23848 6715 23900 6724
rect 23848 6681 23857 6715
rect 23857 6681 23891 6715
rect 23891 6681 23900 6715
rect 23848 6672 23900 6681
rect 28172 6715 28224 6724
rect 20812 6604 20864 6656
rect 21088 6604 21140 6656
rect 22744 6604 22796 6656
rect 25228 6647 25280 6656
rect 25228 6613 25237 6647
rect 25237 6613 25271 6647
rect 25271 6613 25280 6647
rect 25228 6604 25280 6613
rect 26976 6647 27028 6656
rect 26976 6613 26985 6647
rect 26985 6613 27019 6647
rect 27019 6613 27028 6647
rect 28172 6681 28181 6715
rect 28181 6681 28215 6715
rect 28215 6681 28224 6715
rect 28172 6672 28224 6681
rect 26976 6604 27028 6613
rect 27712 6604 27764 6656
rect 28264 6604 28316 6656
rect 8034 6502 8086 6554
rect 8098 6502 8150 6554
rect 8162 6502 8214 6554
rect 8226 6502 8278 6554
rect 8290 6502 8342 6554
rect 15118 6502 15170 6554
rect 15182 6502 15234 6554
rect 15246 6502 15298 6554
rect 15310 6502 15362 6554
rect 15374 6502 15426 6554
rect 22202 6502 22254 6554
rect 22266 6502 22318 6554
rect 22330 6502 22382 6554
rect 22394 6502 22446 6554
rect 22458 6502 22510 6554
rect 29286 6502 29338 6554
rect 29350 6502 29402 6554
rect 29414 6502 29466 6554
rect 29478 6502 29530 6554
rect 29542 6502 29594 6554
rect 1676 6400 1728 6452
rect 5448 6400 5500 6452
rect 3976 6332 4028 6384
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5172 6264 5224 6273
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 5908 6400 5960 6452
rect 6552 6400 6604 6452
rect 9220 6400 9272 6452
rect 11336 6400 11388 6452
rect 12348 6400 12400 6452
rect 12716 6400 12768 6452
rect 13268 6443 13320 6452
rect 13268 6409 13277 6443
rect 13277 6409 13311 6443
rect 13311 6409 13320 6443
rect 13268 6400 13320 6409
rect 14096 6443 14148 6452
rect 14096 6409 14105 6443
rect 14105 6409 14139 6443
rect 14139 6409 14148 6443
rect 14096 6400 14148 6409
rect 14556 6443 14608 6452
rect 14556 6409 14565 6443
rect 14565 6409 14599 6443
rect 14599 6409 14608 6443
rect 14556 6400 14608 6409
rect 16764 6400 16816 6452
rect 18420 6443 18472 6452
rect 18420 6409 18429 6443
rect 18429 6409 18463 6443
rect 18463 6409 18472 6443
rect 18420 6400 18472 6409
rect 18604 6400 18656 6452
rect 19248 6400 19300 6452
rect 19892 6400 19944 6452
rect 20536 6400 20588 6452
rect 22008 6400 22060 6452
rect 23848 6400 23900 6452
rect 24216 6400 24268 6452
rect 26976 6400 27028 6452
rect 27712 6400 27764 6452
rect 28080 6443 28132 6452
rect 28080 6409 28089 6443
rect 28089 6409 28123 6443
rect 28123 6409 28132 6443
rect 28080 6400 28132 6409
rect 6184 6332 6236 6384
rect 6736 6332 6788 6384
rect 7012 6307 7064 6316
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 10968 6332 11020 6384
rect 8484 6264 8536 6316
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9312 6264 9364 6316
rect 10876 6264 10928 6316
rect 12440 6264 12492 6316
rect 13176 6307 13228 6316
rect 10600 6196 10652 6248
rect 10784 6196 10836 6248
rect 10968 6196 11020 6248
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 13268 6264 13320 6316
rect 14188 6264 14240 6316
rect 15476 6332 15528 6384
rect 16028 6332 16080 6384
rect 18052 6332 18104 6384
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 18328 6264 18380 6316
rect 19340 6332 19392 6384
rect 20720 6332 20772 6384
rect 20076 6264 20128 6316
rect 4344 6060 4396 6112
rect 6184 6060 6236 6112
rect 10140 6128 10192 6180
rect 14280 6196 14332 6248
rect 15844 6196 15896 6248
rect 19064 6196 19116 6248
rect 19984 6196 20036 6248
rect 20444 6264 20496 6316
rect 22836 6332 22888 6384
rect 23664 6332 23716 6384
rect 27620 6375 27672 6384
rect 27620 6341 27629 6375
rect 27629 6341 27663 6375
rect 27663 6341 27672 6375
rect 27620 6332 27672 6341
rect 28356 6332 28408 6384
rect 22744 6264 22796 6316
rect 11428 6060 11480 6112
rect 12716 6128 12768 6180
rect 17776 6128 17828 6180
rect 19892 6128 19944 6180
rect 20812 6196 20864 6248
rect 21364 6196 21416 6248
rect 13912 6103 13964 6112
rect 13912 6069 13921 6103
rect 13921 6069 13955 6103
rect 13955 6069 13964 6103
rect 13912 6060 13964 6069
rect 19248 6060 19300 6112
rect 20536 6128 20588 6180
rect 21088 6103 21140 6112
rect 21088 6069 21097 6103
rect 21097 6069 21131 6103
rect 21131 6069 21140 6103
rect 21088 6060 21140 6069
rect 21180 6060 21232 6112
rect 22468 6128 22520 6180
rect 22928 6128 22980 6180
rect 25228 6128 25280 6180
rect 4492 5958 4544 6010
rect 4556 5958 4608 6010
rect 4620 5958 4672 6010
rect 4684 5958 4736 6010
rect 4748 5958 4800 6010
rect 11576 5958 11628 6010
rect 11640 5958 11692 6010
rect 11704 5958 11756 6010
rect 11768 5958 11820 6010
rect 11832 5958 11884 6010
rect 18660 5958 18712 6010
rect 18724 5958 18776 6010
rect 18788 5958 18840 6010
rect 18852 5958 18904 6010
rect 18916 5958 18968 6010
rect 25744 5958 25796 6010
rect 25808 5958 25860 6010
rect 25872 5958 25924 6010
rect 25936 5958 25988 6010
rect 26000 5958 26052 6010
rect 1400 5899 1452 5908
rect 1400 5865 1409 5899
rect 1409 5865 1443 5899
rect 1443 5865 1452 5899
rect 1400 5856 1452 5865
rect 5172 5856 5224 5908
rect 6184 5856 6236 5908
rect 9036 5856 9088 5908
rect 10600 5899 10652 5908
rect 10600 5865 10609 5899
rect 10609 5865 10643 5899
rect 10643 5865 10652 5899
rect 10600 5856 10652 5865
rect 14188 5856 14240 5908
rect 14464 5856 14516 5908
rect 15108 5856 15160 5908
rect 15844 5856 15896 5908
rect 17132 5856 17184 5908
rect 19524 5856 19576 5908
rect 21272 5856 21324 5908
rect 22560 5899 22612 5908
rect 22560 5865 22569 5899
rect 22569 5865 22603 5899
rect 22603 5865 22612 5899
rect 22560 5856 22612 5865
rect 26792 5856 26844 5908
rect 4896 5788 4948 5840
rect 5908 5695 5960 5704
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 6644 5695 6696 5704
rect 6644 5661 6653 5695
rect 6653 5661 6687 5695
rect 6687 5661 6696 5695
rect 6644 5652 6696 5661
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 9036 5652 9088 5704
rect 13820 5788 13872 5840
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 15108 5720 15160 5772
rect 16856 5720 16908 5772
rect 17960 5788 18012 5840
rect 21916 5788 21968 5840
rect 28172 5788 28224 5840
rect 18512 5720 18564 5772
rect 13176 5584 13228 5636
rect 13820 5652 13872 5704
rect 17040 5652 17092 5704
rect 19340 5720 19392 5772
rect 19616 5720 19668 5772
rect 20536 5763 20588 5772
rect 20536 5729 20545 5763
rect 20545 5729 20579 5763
rect 20579 5729 20588 5763
rect 20536 5720 20588 5729
rect 22836 5720 22888 5772
rect 19432 5695 19484 5704
rect 19432 5661 19441 5695
rect 19441 5661 19475 5695
rect 19475 5661 19484 5695
rect 19432 5652 19484 5661
rect 15476 5584 15528 5636
rect 17500 5584 17552 5636
rect 28724 5695 28776 5704
rect 28724 5661 28733 5695
rect 28733 5661 28767 5695
rect 28767 5661 28776 5695
rect 28724 5652 28776 5661
rect 21180 5627 21232 5636
rect 21180 5593 21205 5627
rect 21205 5593 21232 5627
rect 21180 5584 21232 5593
rect 7840 5559 7892 5568
rect 7840 5525 7849 5559
rect 7849 5525 7883 5559
rect 7883 5525 7892 5559
rect 7840 5516 7892 5525
rect 17040 5516 17092 5568
rect 17776 5516 17828 5568
rect 22468 5516 22520 5568
rect 8034 5414 8086 5466
rect 8098 5414 8150 5466
rect 8162 5414 8214 5466
rect 8226 5414 8278 5466
rect 8290 5414 8342 5466
rect 15118 5414 15170 5466
rect 15182 5414 15234 5466
rect 15246 5414 15298 5466
rect 15310 5414 15362 5466
rect 15374 5414 15426 5466
rect 22202 5414 22254 5466
rect 22266 5414 22318 5466
rect 22330 5414 22382 5466
rect 22394 5414 22446 5466
rect 22458 5414 22510 5466
rect 29286 5414 29338 5466
rect 29350 5414 29402 5466
rect 29414 5414 29466 5466
rect 29478 5414 29530 5466
rect 29542 5414 29594 5466
rect 6644 5312 6696 5364
rect 7932 5312 7984 5364
rect 10048 5355 10100 5364
rect 10048 5321 10057 5355
rect 10057 5321 10091 5355
rect 10091 5321 10100 5355
rect 10048 5312 10100 5321
rect 10876 5355 10928 5364
rect 10876 5321 10885 5355
rect 10885 5321 10919 5355
rect 10919 5321 10928 5355
rect 10876 5312 10928 5321
rect 13820 5355 13872 5364
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 13820 5312 13872 5321
rect 14372 5312 14424 5364
rect 17040 5312 17092 5364
rect 18052 5312 18104 5364
rect 18328 5312 18380 5364
rect 22560 5312 22612 5364
rect 23020 5312 23072 5364
rect 28724 5355 28776 5364
rect 28724 5321 28733 5355
rect 28733 5321 28767 5355
rect 28767 5321 28776 5355
rect 28724 5312 28776 5321
rect 7196 5219 7248 5228
rect 7196 5185 7205 5219
rect 7205 5185 7239 5219
rect 7239 5185 7248 5219
rect 7196 5176 7248 5185
rect 21824 5219 21876 5228
rect 21824 5185 21833 5219
rect 21833 5185 21867 5219
rect 21867 5185 21876 5219
rect 21824 5176 21876 5185
rect 21916 5219 21968 5228
rect 21916 5185 21925 5219
rect 21925 5185 21959 5219
rect 21959 5185 21968 5219
rect 21916 5176 21968 5185
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 7840 5108 7892 5160
rect 15936 5108 15988 5160
rect 22192 5287 22244 5296
rect 22192 5253 22201 5287
rect 22201 5253 22235 5287
rect 22235 5253 22244 5287
rect 22192 5244 22244 5253
rect 22560 5176 22612 5228
rect 23388 5176 23440 5228
rect 23756 5176 23808 5228
rect 22468 5083 22520 5092
rect 22468 5049 22477 5083
rect 22477 5049 22511 5083
rect 22511 5049 22520 5083
rect 22468 5040 22520 5049
rect 23480 5040 23532 5092
rect 6736 4972 6788 5024
rect 8484 4972 8536 5024
rect 19156 5015 19208 5024
rect 19156 4981 19165 5015
rect 19165 4981 19199 5015
rect 19199 4981 19208 5015
rect 19156 4972 19208 4981
rect 19248 4972 19300 5024
rect 23112 4972 23164 5024
rect 4492 4870 4544 4922
rect 4556 4870 4608 4922
rect 4620 4870 4672 4922
rect 4684 4870 4736 4922
rect 4748 4870 4800 4922
rect 11576 4870 11628 4922
rect 11640 4870 11692 4922
rect 11704 4870 11756 4922
rect 11768 4870 11820 4922
rect 11832 4870 11884 4922
rect 18660 4870 18712 4922
rect 18724 4870 18776 4922
rect 18788 4870 18840 4922
rect 18852 4870 18904 4922
rect 18916 4870 18968 4922
rect 25744 4870 25796 4922
rect 25808 4870 25860 4922
rect 25872 4870 25924 4922
rect 25936 4870 25988 4922
rect 26000 4870 26052 4922
rect 4344 4768 4396 4820
rect 6460 4768 6512 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 10508 4811 10560 4820
rect 10508 4777 10517 4811
rect 10517 4777 10551 4811
rect 10551 4777 10560 4811
rect 10508 4768 10560 4777
rect 14372 4811 14424 4820
rect 14372 4777 14381 4811
rect 14381 4777 14415 4811
rect 14415 4777 14424 4811
rect 14372 4768 14424 4777
rect 15200 4768 15252 4820
rect 15476 4768 15528 4820
rect 19248 4768 19300 4820
rect 20260 4768 20312 4820
rect 23388 4811 23440 4820
rect 14464 4700 14516 4752
rect 17776 4743 17828 4752
rect 17776 4709 17785 4743
rect 17785 4709 17819 4743
rect 17819 4709 17828 4743
rect 17776 4700 17828 4709
rect 7196 4632 7248 4684
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 7104 4564 7156 4616
rect 9772 4632 9824 4684
rect 10508 4564 10560 4616
rect 1584 4496 1636 4548
rect 10048 4496 10100 4548
rect 10600 4496 10652 4548
rect 12624 4632 12676 4684
rect 19156 4632 19208 4684
rect 20536 4675 20588 4684
rect 20536 4641 20545 4675
rect 20545 4641 20579 4675
rect 20579 4641 20588 4675
rect 20536 4632 20588 4641
rect 14280 4564 14332 4616
rect 14556 4564 14608 4616
rect 15200 4607 15252 4616
rect 15200 4573 15209 4607
rect 15209 4573 15243 4607
rect 15243 4573 15252 4607
rect 20076 4607 20128 4616
rect 15200 4564 15252 4573
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 20628 4564 20680 4616
rect 23388 4777 23397 4811
rect 23397 4777 23431 4811
rect 23431 4777 23440 4811
rect 23388 4768 23440 4777
rect 22008 4743 22060 4752
rect 22008 4709 22017 4743
rect 22017 4709 22051 4743
rect 22051 4709 22060 4743
rect 22008 4700 22060 4709
rect 22468 4564 22520 4616
rect 23664 4700 23716 4752
rect 19340 4496 19392 4548
rect 14372 4428 14424 4480
rect 20720 4428 20772 4480
rect 23204 4428 23256 4480
rect 8034 4326 8086 4378
rect 8098 4326 8150 4378
rect 8162 4326 8214 4378
rect 8226 4326 8278 4378
rect 8290 4326 8342 4378
rect 15118 4326 15170 4378
rect 15182 4326 15234 4378
rect 15246 4326 15298 4378
rect 15310 4326 15362 4378
rect 15374 4326 15426 4378
rect 22202 4326 22254 4378
rect 22266 4326 22318 4378
rect 22330 4326 22382 4378
rect 22394 4326 22446 4378
rect 22458 4326 22510 4378
rect 29286 4326 29338 4378
rect 29350 4326 29402 4378
rect 29414 4326 29466 4378
rect 29478 4326 29530 4378
rect 29542 4326 29594 4378
rect 10600 4224 10652 4276
rect 15936 4267 15988 4276
rect 1584 4199 1636 4208
rect 1584 4165 1593 4199
rect 1593 4165 1627 4199
rect 1627 4165 1636 4199
rect 1584 4156 1636 4165
rect 9772 4088 9824 4140
rect 2964 4063 3016 4072
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 10968 4088 11020 4140
rect 11980 4088 12032 4140
rect 14924 4156 14976 4208
rect 15200 4199 15252 4208
rect 15200 4165 15227 4199
rect 15227 4165 15252 4199
rect 15200 4156 15252 4165
rect 15936 4233 15945 4267
rect 15945 4233 15979 4267
rect 15979 4233 15988 4267
rect 15936 4224 15988 4233
rect 20720 4224 20772 4276
rect 22560 4224 22612 4276
rect 16764 4156 16816 4208
rect 14280 4131 14332 4140
rect 13544 4020 13596 4072
rect 10048 3952 10100 4004
rect 11428 3952 11480 4004
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 17776 4156 17828 4208
rect 18052 4156 18104 4208
rect 17960 4088 18012 4140
rect 20904 4131 20956 4140
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 21824 4131 21876 4140
rect 21824 4097 21833 4131
rect 21833 4097 21867 4131
rect 21867 4097 21876 4131
rect 21824 4088 21876 4097
rect 21916 4131 21968 4140
rect 21916 4097 21925 4131
rect 21925 4097 21959 4131
rect 21959 4097 21968 4131
rect 21916 4088 21968 4097
rect 23204 4131 23256 4140
rect 14464 4063 14516 4072
rect 14464 4029 14473 4063
rect 14473 4029 14507 4063
rect 14507 4029 14516 4063
rect 14464 4020 14516 4029
rect 15016 3995 15068 4004
rect 1676 3884 1728 3936
rect 10968 3884 11020 3936
rect 15016 3961 15025 3995
rect 15025 3961 15059 3995
rect 15059 3961 15068 3995
rect 15016 3952 15068 3961
rect 17776 4020 17828 4072
rect 20812 4063 20864 4072
rect 19340 3952 19392 4004
rect 20812 4029 20821 4063
rect 20821 4029 20855 4063
rect 20855 4029 20864 4063
rect 20812 4020 20864 4029
rect 21456 4020 21508 4072
rect 23204 4097 23213 4131
rect 23213 4097 23247 4131
rect 23247 4097 23256 4131
rect 23204 4088 23256 4097
rect 23296 4131 23348 4140
rect 23296 4097 23305 4131
rect 23305 4097 23339 4131
rect 23339 4097 23348 4131
rect 23296 4088 23348 4097
rect 23664 4063 23716 4072
rect 23664 4029 23673 4063
rect 23673 4029 23707 4063
rect 23707 4029 23716 4063
rect 23664 4020 23716 4029
rect 23848 4088 23900 4140
rect 20996 3952 21048 4004
rect 22744 3952 22796 4004
rect 23020 3952 23072 4004
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 15292 3884 15344 3936
rect 15844 3884 15896 3936
rect 17224 3884 17276 3936
rect 17868 3884 17920 3936
rect 17960 3927 18012 3936
rect 17960 3893 17969 3927
rect 17969 3893 18003 3927
rect 18003 3893 18012 3927
rect 22928 3927 22980 3936
rect 17960 3884 18012 3893
rect 22928 3893 22937 3927
rect 22937 3893 22971 3927
rect 22971 3893 22980 3927
rect 22928 3884 22980 3893
rect 23480 3884 23532 3936
rect 28632 3927 28684 3936
rect 28632 3893 28641 3927
rect 28641 3893 28675 3927
rect 28675 3893 28684 3927
rect 28632 3884 28684 3893
rect 4492 3782 4544 3834
rect 4556 3782 4608 3834
rect 4620 3782 4672 3834
rect 4684 3782 4736 3834
rect 4748 3782 4800 3834
rect 11576 3782 11628 3834
rect 11640 3782 11692 3834
rect 11704 3782 11756 3834
rect 11768 3782 11820 3834
rect 11832 3782 11884 3834
rect 18660 3782 18712 3834
rect 18724 3782 18776 3834
rect 18788 3782 18840 3834
rect 18852 3782 18904 3834
rect 18916 3782 18968 3834
rect 25744 3782 25796 3834
rect 25808 3782 25860 3834
rect 25872 3782 25924 3834
rect 25936 3782 25988 3834
rect 26000 3782 26052 3834
rect 13544 3723 13596 3732
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 10968 3544 11020 3596
rect 11428 3544 11480 3596
rect 13544 3689 13553 3723
rect 13553 3689 13587 3723
rect 13587 3689 13596 3723
rect 13544 3680 13596 3689
rect 13636 3680 13688 3732
rect 15200 3680 15252 3732
rect 16580 3680 16632 3732
rect 20076 3723 20128 3732
rect 10600 3451 10652 3460
rect 10600 3417 10609 3451
rect 10609 3417 10643 3451
rect 10643 3417 10652 3451
rect 10600 3408 10652 3417
rect 11980 3476 12032 3528
rect 12624 3519 12676 3528
rect 12624 3485 12633 3519
rect 12633 3485 12667 3519
rect 12667 3485 12676 3519
rect 12624 3476 12676 3485
rect 11520 3408 11572 3460
rect 13360 3476 13412 3528
rect 15844 3655 15896 3664
rect 15844 3621 15853 3655
rect 15853 3621 15887 3655
rect 15887 3621 15896 3655
rect 15844 3612 15896 3621
rect 17316 3655 17368 3664
rect 17316 3621 17325 3655
rect 17325 3621 17359 3655
rect 17359 3621 17368 3655
rect 17316 3612 17368 3621
rect 18144 3612 18196 3664
rect 16580 3587 16632 3596
rect 16580 3553 16589 3587
rect 16589 3553 16623 3587
rect 16623 3553 16632 3587
rect 16580 3544 16632 3553
rect 17224 3544 17276 3596
rect 13912 3476 13964 3528
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 17684 3519 17736 3528
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 12532 3383 12584 3392
rect 12532 3349 12541 3383
rect 12541 3349 12575 3383
rect 12575 3349 12584 3383
rect 12532 3340 12584 3349
rect 15292 3340 15344 3392
rect 15568 3340 15620 3392
rect 17684 3485 17693 3519
rect 17693 3485 17727 3519
rect 17727 3485 17736 3519
rect 17684 3476 17736 3485
rect 20076 3689 20085 3723
rect 20085 3689 20119 3723
rect 20119 3689 20128 3723
rect 20076 3680 20128 3689
rect 20812 3723 20864 3732
rect 20812 3689 20821 3723
rect 20821 3689 20855 3723
rect 20855 3689 20864 3723
rect 20812 3680 20864 3689
rect 22100 3680 22152 3732
rect 23296 3723 23348 3732
rect 23296 3689 23305 3723
rect 23305 3689 23339 3723
rect 23339 3689 23348 3723
rect 23296 3680 23348 3689
rect 23664 3680 23716 3732
rect 23112 3612 23164 3664
rect 17868 3476 17920 3528
rect 18972 3476 19024 3528
rect 17960 3408 18012 3460
rect 20904 3519 20956 3528
rect 18052 3340 18104 3392
rect 20536 3340 20588 3392
rect 20904 3485 20913 3519
rect 20913 3485 20947 3519
rect 20947 3485 20956 3519
rect 20904 3476 20956 3485
rect 20996 3519 21048 3528
rect 20996 3485 21005 3519
rect 21005 3485 21039 3519
rect 21039 3485 21048 3519
rect 21456 3519 21508 3528
rect 20996 3476 21048 3485
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 21456 3476 21508 3485
rect 21824 3544 21876 3596
rect 21916 3476 21968 3528
rect 23480 3544 23532 3596
rect 22744 3476 22796 3528
rect 23848 3476 23900 3528
rect 23020 3408 23072 3460
rect 27436 3340 27488 3392
rect 8034 3238 8086 3290
rect 8098 3238 8150 3290
rect 8162 3238 8214 3290
rect 8226 3238 8278 3290
rect 8290 3238 8342 3290
rect 15118 3238 15170 3290
rect 15182 3238 15234 3290
rect 15246 3238 15298 3290
rect 15310 3238 15362 3290
rect 15374 3238 15426 3290
rect 22202 3238 22254 3290
rect 22266 3238 22318 3290
rect 22330 3238 22382 3290
rect 22394 3238 22446 3290
rect 22458 3238 22510 3290
rect 29286 3238 29338 3290
rect 29350 3238 29402 3290
rect 29414 3238 29466 3290
rect 29478 3238 29530 3290
rect 29542 3238 29594 3290
rect 10048 3136 10100 3188
rect 2412 3068 2464 3120
rect 10600 3136 10652 3188
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 12624 3136 12676 3188
rect 13912 3179 13964 3188
rect 13912 3145 13921 3179
rect 13921 3145 13955 3179
rect 13955 3145 13964 3179
rect 13912 3136 13964 3145
rect 14464 3136 14516 3188
rect 17684 3136 17736 3188
rect 2044 3000 2096 3052
rect 10876 3000 10928 3052
rect 14096 3068 14148 3120
rect 18972 3111 19024 3120
rect 12532 3000 12584 3052
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14924 3000 14976 3052
rect 18972 3077 18981 3111
rect 18981 3077 19015 3111
rect 19015 3077 19024 3111
rect 18972 3068 19024 3077
rect 21456 3136 21508 3188
rect 23020 3136 23072 3188
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 18236 3000 18288 3052
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 20720 3043 20772 3052
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 20996 3068 21048 3120
rect 28632 3043 28684 3052
rect 28632 3009 28641 3043
rect 28641 3009 28675 3043
rect 28675 3009 28684 3043
rect 28632 3000 28684 3009
rect 21824 2975 21876 2984
rect 21824 2941 21833 2975
rect 21833 2941 21867 2975
rect 21867 2941 21876 2975
rect 21824 2932 21876 2941
rect 15568 2864 15620 2916
rect 29644 2864 29696 2916
rect 20 2796 72 2848
rect 14096 2839 14148 2848
rect 14096 2805 14105 2839
rect 14105 2805 14139 2839
rect 14139 2805 14148 2839
rect 14096 2796 14148 2805
rect 16764 2796 16816 2848
rect 19248 2796 19300 2848
rect 4492 2694 4544 2746
rect 4556 2694 4608 2746
rect 4620 2694 4672 2746
rect 4684 2694 4736 2746
rect 4748 2694 4800 2746
rect 11576 2694 11628 2746
rect 11640 2694 11692 2746
rect 11704 2694 11756 2746
rect 11768 2694 11820 2746
rect 11832 2694 11884 2746
rect 18660 2694 18712 2746
rect 18724 2694 18776 2746
rect 18788 2694 18840 2746
rect 18852 2694 18904 2746
rect 18916 2694 18968 2746
rect 25744 2694 25796 2746
rect 25808 2694 25860 2746
rect 25872 2694 25924 2746
rect 25936 2694 25988 2746
rect 26000 2694 26052 2746
rect 6736 2592 6788 2644
rect 14004 2592 14056 2644
rect 14924 2592 14976 2644
rect 19616 2592 19668 2644
rect 20904 2635 20956 2644
rect 20904 2601 20913 2635
rect 20913 2601 20947 2635
rect 20947 2601 20956 2635
rect 20904 2592 20956 2601
rect 27988 2635 28040 2644
rect 27988 2601 27997 2635
rect 27997 2601 28031 2635
rect 28031 2601 28040 2635
rect 27988 2592 28040 2601
rect 4252 2431 4304 2440
rect 4252 2397 4261 2431
rect 4261 2397 4295 2431
rect 4295 2397 4304 2431
rect 4252 2388 4304 2397
rect 1952 2320 2004 2372
rect 8576 2388 8628 2440
rect 3884 2252 3936 2304
rect 5816 2295 5868 2304
rect 5816 2261 5825 2295
rect 5825 2261 5859 2295
rect 5859 2261 5868 2295
rect 5816 2252 5868 2261
rect 8392 2252 8444 2304
rect 10324 2252 10376 2304
rect 22928 2524 22980 2576
rect 24032 2524 24084 2576
rect 18236 2499 18288 2508
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 12256 2320 12308 2372
rect 16580 2320 16632 2372
rect 16764 2320 16816 2372
rect 18236 2465 18245 2499
rect 18245 2465 18279 2499
rect 18279 2465 18288 2499
rect 18236 2456 18288 2465
rect 19156 2456 19208 2508
rect 18696 2388 18748 2440
rect 19248 2431 19300 2440
rect 19248 2397 19257 2431
rect 19257 2397 19291 2431
rect 19291 2397 19300 2431
rect 19248 2388 19300 2397
rect 19800 2456 19852 2508
rect 20996 2431 21048 2440
rect 20996 2397 21005 2431
rect 21005 2397 21039 2431
rect 21039 2397 21048 2431
rect 20996 2388 21048 2397
rect 21824 2431 21876 2440
rect 21824 2397 21833 2431
rect 21833 2397 21867 2431
rect 21867 2397 21876 2431
rect 21824 2388 21876 2397
rect 19892 2320 19944 2372
rect 23204 2320 23256 2372
rect 25136 2320 25188 2372
rect 27712 2320 27764 2372
rect 14832 2252 14884 2304
rect 21272 2252 21324 2304
rect 8034 2150 8086 2202
rect 8098 2150 8150 2202
rect 8162 2150 8214 2202
rect 8226 2150 8278 2202
rect 8290 2150 8342 2202
rect 15118 2150 15170 2202
rect 15182 2150 15234 2202
rect 15246 2150 15298 2202
rect 15310 2150 15362 2202
rect 15374 2150 15426 2202
rect 22202 2150 22254 2202
rect 22266 2150 22318 2202
rect 22330 2150 22382 2202
rect 22394 2150 22446 2202
rect 22458 2150 22510 2202
rect 29286 2150 29338 2202
rect 29350 2150 29402 2202
rect 29414 2150 29466 2202
rect 29478 2150 29530 2202
rect 29542 2150 29594 2202
<< metal2 >>
rect 662 31965 718 32765
rect 2594 31965 2650 32765
rect 5170 31965 5226 32765
rect 7102 31965 7158 32765
rect 9034 31965 9090 32765
rect 11610 31965 11666 32765
rect 13542 31965 13598 32765
rect 15474 31965 15530 32765
rect 18050 31965 18106 32765
rect 19982 31965 20038 32765
rect 21914 31965 21970 32765
rect 24490 31965 24546 32765
rect 26422 31965 26478 32765
rect 28354 31965 28410 32765
rect 30286 31965 30342 32765
rect 676 30326 704 31965
rect 1858 31376 1914 31385
rect 1858 31311 1914 31320
rect 664 30320 716 30326
rect 664 30262 716 30268
rect 1308 30320 1360 30326
rect 1308 30262 1360 30268
rect 1320 29782 1348 30262
rect 1308 29776 1360 29782
rect 1308 29718 1360 29724
rect 1492 29504 1544 29510
rect 1492 29446 1544 29452
rect 1504 29345 1532 29446
rect 1490 29336 1546 29345
rect 1490 29271 1546 29280
rect 1872 29238 1900 31311
rect 2608 30326 2636 31965
rect 2596 30320 2648 30326
rect 2596 30262 2648 30268
rect 2044 30116 2096 30122
rect 2044 30058 2096 30064
rect 1860 29232 1912 29238
rect 1860 29174 1912 29180
rect 1872 28762 1900 29174
rect 1860 28756 1912 28762
rect 1860 28698 1912 28704
rect 1584 26988 1636 26994
rect 1584 26930 1636 26936
rect 1596 26625 1624 26930
rect 1860 26784 1912 26790
rect 1860 26726 1912 26732
rect 1582 26616 1638 26625
rect 1582 26551 1584 26560
rect 1636 26551 1638 26560
rect 1584 26522 1636 26528
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1412 24585 1440 24754
rect 1584 24608 1636 24614
rect 1398 24576 1454 24585
rect 1584 24550 1636 24556
rect 1398 24511 1454 24520
rect 1412 24410 1440 24511
rect 1596 24410 1624 24550
rect 1400 24404 1452 24410
rect 1400 24346 1452 24352
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1596 22642 1624 22918
rect 1584 22636 1636 22642
rect 1584 22578 1636 22584
rect 1596 22545 1624 22578
rect 1582 22536 1638 22545
rect 1582 22471 1638 22480
rect 1766 22536 1822 22545
rect 1766 22471 1768 22480
rect 1820 22471 1822 22480
rect 1768 22442 1820 22448
rect 1676 22024 1728 22030
rect 1676 21966 1728 21972
rect 1688 20330 1716 21966
rect 1872 20602 1900 26726
rect 2056 22794 2084 30058
rect 2608 29850 2636 30262
rect 5184 30122 5212 31965
rect 7116 30258 7144 31965
rect 8034 30492 8342 30501
rect 8034 30490 8040 30492
rect 8096 30490 8120 30492
rect 8176 30490 8200 30492
rect 8256 30490 8280 30492
rect 8336 30490 8342 30492
rect 8096 30438 8098 30490
rect 8278 30438 8280 30490
rect 8034 30436 8040 30438
rect 8096 30436 8120 30438
rect 8176 30436 8200 30438
rect 8256 30436 8280 30438
rect 8336 30436 8342 30438
rect 8034 30427 8342 30436
rect 5540 30252 5592 30258
rect 5540 30194 5592 30200
rect 7104 30252 7156 30258
rect 7104 30194 7156 30200
rect 7840 30252 7892 30258
rect 7840 30194 7892 30200
rect 5172 30116 5224 30122
rect 5172 30058 5224 30064
rect 4492 29948 4800 29957
rect 4492 29946 4498 29948
rect 4554 29946 4578 29948
rect 4634 29946 4658 29948
rect 4714 29946 4738 29948
rect 4794 29946 4800 29948
rect 4554 29894 4556 29946
rect 4736 29894 4738 29946
rect 4492 29892 4498 29894
rect 4554 29892 4578 29894
rect 4634 29892 4658 29894
rect 4714 29892 4738 29894
rect 4794 29892 4800 29894
rect 4492 29883 4800 29892
rect 2596 29844 2648 29850
rect 2596 29786 2648 29792
rect 2136 29640 2188 29646
rect 2136 29582 2188 29588
rect 2148 29102 2176 29582
rect 2136 29096 2188 29102
rect 2136 29038 2188 29044
rect 1964 22766 2084 22794
rect 1860 20596 1912 20602
rect 1860 20538 1912 20544
rect 1676 20324 1728 20330
rect 1676 20266 1728 20272
rect 1688 19854 1716 20266
rect 1676 19848 1728 19854
rect 1490 19816 1546 19825
rect 1676 19790 1728 19796
rect 1490 19751 1546 19760
rect 1504 19718 1532 19751
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 15745 1440 16050
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1504 13274 1532 18566
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17814 1624 18226
rect 1584 17808 1636 17814
rect 1582 17776 1584 17785
rect 1636 17776 1638 17785
rect 1582 17711 1638 17720
rect 1688 16574 1716 19790
rect 1872 19378 1900 20538
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1964 19242 1992 22766
rect 1952 19236 2004 19242
rect 1952 19178 2004 19184
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1780 16794 1808 17138
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1688 16546 1808 16574
rect 1504 13246 1716 13274
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1504 13025 1532 13126
rect 1490 13016 1546 13025
rect 1490 12951 1546 12960
rect 1490 10976 1546 10985
rect 1490 10911 1546 10920
rect 1504 10810 1532 10911
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1596 8566 1624 8871
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1596 8090 1624 8502
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1688 6458 1716 13246
rect 1780 12458 1808 16546
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1872 13870 1900 14214
rect 1964 13938 1992 16934
rect 2148 14414 2176 29038
rect 4988 29028 5040 29034
rect 4988 28970 5040 28976
rect 4492 28860 4800 28869
rect 4492 28858 4498 28860
rect 4554 28858 4578 28860
rect 4634 28858 4658 28860
rect 4714 28858 4738 28860
rect 4794 28858 4800 28860
rect 4554 28806 4556 28858
rect 4736 28806 4738 28858
rect 4492 28804 4498 28806
rect 4554 28804 4578 28806
rect 4634 28804 4658 28806
rect 4714 28804 4738 28806
rect 4794 28804 4800 28806
rect 4492 28795 4800 28804
rect 4492 27772 4800 27781
rect 4492 27770 4498 27772
rect 4554 27770 4578 27772
rect 4634 27770 4658 27772
rect 4714 27770 4738 27772
rect 4794 27770 4800 27772
rect 4554 27718 4556 27770
rect 4736 27718 4738 27770
rect 4492 27716 4498 27718
rect 4554 27716 4578 27718
rect 4634 27716 4658 27718
rect 4714 27716 4738 27718
rect 4794 27716 4800 27718
rect 4492 27707 4800 27716
rect 4492 26684 4800 26693
rect 4492 26682 4498 26684
rect 4554 26682 4578 26684
rect 4634 26682 4658 26684
rect 4714 26682 4738 26684
rect 4794 26682 4800 26684
rect 4554 26630 4556 26682
rect 4736 26630 4738 26682
rect 4492 26628 4498 26630
rect 4554 26628 4578 26630
rect 4634 26628 4658 26630
rect 4714 26628 4738 26630
rect 4794 26628 4800 26630
rect 4492 26619 4800 26628
rect 4344 25900 4396 25906
rect 4344 25842 4396 25848
rect 4252 25832 4304 25838
rect 4252 25774 4304 25780
rect 4264 25498 4292 25774
rect 4252 25492 4304 25498
rect 4252 25434 4304 25440
rect 4356 24206 4384 25842
rect 4492 25596 4800 25605
rect 4492 25594 4498 25596
rect 4554 25594 4578 25596
rect 4634 25594 4658 25596
rect 4714 25594 4738 25596
rect 4794 25594 4800 25596
rect 4554 25542 4556 25594
rect 4736 25542 4738 25594
rect 4492 25540 4498 25542
rect 4554 25540 4578 25542
rect 4634 25540 4658 25542
rect 4714 25540 4738 25542
rect 4794 25540 4800 25542
rect 4492 25531 4800 25540
rect 4620 25288 4672 25294
rect 4620 25230 4672 25236
rect 4632 24750 4660 25230
rect 5000 24954 5028 28970
rect 5552 28558 5580 30194
rect 6736 29164 6788 29170
rect 6736 29106 6788 29112
rect 5816 29028 5868 29034
rect 5816 28970 5868 28976
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 5356 26784 5408 26790
rect 5356 26726 5408 26732
rect 5368 26489 5396 26726
rect 5552 26586 5580 26930
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5724 26512 5776 26518
rect 5354 26480 5410 26489
rect 5724 26454 5776 26460
rect 5354 26415 5410 26424
rect 5080 26376 5132 26382
rect 5080 26318 5132 26324
rect 5092 26042 5120 26318
rect 5368 26314 5396 26415
rect 5736 26382 5764 26454
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5724 26376 5776 26382
rect 5724 26318 5776 26324
rect 5356 26308 5408 26314
rect 5356 26250 5408 26256
rect 5080 26036 5132 26042
rect 5080 25978 5132 25984
rect 5080 25900 5132 25906
rect 5080 25842 5132 25848
rect 5264 25900 5316 25906
rect 5264 25842 5316 25848
rect 5092 25294 5120 25842
rect 5276 25498 5304 25842
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 5264 25288 5316 25294
rect 5264 25230 5316 25236
rect 5092 25158 5120 25230
rect 5080 25152 5132 25158
rect 5080 25094 5132 25100
rect 4988 24948 5040 24954
rect 4988 24890 5040 24896
rect 5092 24834 5120 25094
rect 5172 24948 5224 24954
rect 5172 24890 5224 24896
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 5000 24806 5120 24834
rect 4620 24744 4672 24750
rect 4620 24686 4672 24692
rect 4492 24508 4800 24517
rect 4492 24506 4498 24508
rect 4554 24506 4578 24508
rect 4634 24506 4658 24508
rect 4714 24506 4738 24508
rect 4794 24506 4800 24508
rect 4554 24454 4556 24506
rect 4736 24454 4738 24506
rect 4492 24452 4498 24454
rect 4554 24452 4578 24454
rect 4634 24452 4658 24454
rect 4714 24452 4738 24454
rect 4794 24452 4800 24454
rect 4492 24443 4800 24452
rect 4908 24206 4936 24754
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4344 24200 4396 24206
rect 4344 24142 4396 24148
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 3976 23520 4028 23526
rect 3976 23462 4028 23468
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3332 22704 3384 22710
rect 3330 22672 3332 22681
rect 3384 22672 3386 22681
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 3056 22636 3108 22642
rect 3330 22607 3386 22616
rect 3056 22578 3108 22584
rect 2240 22234 2268 22578
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2964 22092 3016 22098
rect 2964 22034 3016 22040
rect 2976 21350 3004 22034
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2688 19848 2740 19854
rect 2740 19808 2820 19836
rect 2688 19790 2740 19796
rect 2240 18970 2268 19790
rect 2792 19514 2820 19808
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2412 19440 2464 19446
rect 2412 19382 2464 19388
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2332 19174 2360 19314
rect 2424 19174 2452 19382
rect 2504 19372 2556 19378
rect 2504 19314 2556 19320
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2332 18766 2360 19110
rect 2424 18834 2452 19110
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2516 18698 2544 19314
rect 2504 18692 2556 18698
rect 2504 18634 2556 18640
rect 2596 18692 2648 18698
rect 2596 18634 2648 18640
rect 2516 18426 2544 18634
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2608 18358 2636 18634
rect 2596 18352 2648 18358
rect 2596 18294 2648 18300
rect 2228 17604 2280 17610
rect 2228 17546 2280 17552
rect 2240 16658 2268 17546
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2884 16794 2912 17478
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 2136 13728 2188 13734
rect 2136 13670 2188 13676
rect 1780 12430 1900 12458
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 1780 11354 1808 12242
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1872 8430 1900 12430
rect 2148 12238 2176 13670
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2148 10470 2176 11086
rect 2240 10674 2268 16594
rect 2884 16590 2912 16730
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2240 9654 2268 10610
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2332 9178 2360 11698
rect 2424 9926 2452 16526
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 11762 2636 12038
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2424 9586 2452 9862
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2332 8498 2360 8910
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1872 7206 1900 8230
rect 1964 7886 1992 8230
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 6225 1440 6258
rect 1688 6225 1716 6394
rect 1398 6216 1454 6225
rect 1398 6151 1454 6160
rect 1674 6216 1730 6225
rect 1674 6151 1730 6160
rect 1412 5914 1440 6151
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1584 4548 1636 4554
rect 1584 4490 1636 4496
rect 1596 4214 1624 4490
rect 1584 4208 1636 4214
rect 1582 4176 1584 4185
rect 1636 4176 1638 4185
rect 1582 4111 1638 4120
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1688 3534 1716 3878
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 32 800 60 2790
rect 1504 2145 1532 3334
rect 2056 3058 2084 7686
rect 2424 3126 2452 9522
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2516 7954 2544 9318
rect 2700 8537 2728 13126
rect 2976 12434 3004 21286
rect 2884 12406 3004 12434
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2686 8528 2742 8537
rect 2686 8463 2742 8472
rect 2792 8294 2820 8978
rect 2884 8498 2912 12406
rect 3068 11898 3096 22578
rect 3516 22432 3568 22438
rect 3516 22374 3568 22380
rect 3528 21486 3556 22374
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3160 19514 3188 20402
rect 3252 20058 3280 20402
rect 3240 20052 3292 20058
rect 3240 19994 3292 20000
rect 3712 19786 3740 21286
rect 3700 19780 3752 19786
rect 3700 19722 3752 19728
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3804 16182 3832 22918
rect 3988 22642 4016 23462
rect 4172 23118 4200 24142
rect 4252 24064 4304 24070
rect 4252 24006 4304 24012
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4264 22642 4292 24006
rect 4356 23594 4384 24142
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4632 23866 4660 24074
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4344 23588 4396 23594
rect 4344 23530 4396 23536
rect 4356 23322 4384 23530
rect 4492 23420 4800 23429
rect 4492 23418 4498 23420
rect 4554 23418 4578 23420
rect 4634 23418 4658 23420
rect 4714 23418 4738 23420
rect 4794 23418 4800 23420
rect 4554 23366 4556 23418
rect 4736 23366 4738 23418
rect 4492 23364 4498 23366
rect 4554 23364 4578 23366
rect 4634 23364 4658 23366
rect 4714 23364 4738 23366
rect 4794 23364 4800 23366
rect 4492 23355 4800 23364
rect 4344 23316 4396 23322
rect 4344 23258 4396 23264
rect 5000 23118 5028 24806
rect 5080 24744 5132 24750
rect 5080 24686 5132 24692
rect 5092 24206 5120 24686
rect 5080 24200 5132 24206
rect 5080 24142 5132 24148
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 3976 22636 4028 22642
rect 3976 22578 4028 22584
rect 4252 22636 4304 22642
rect 4252 22578 4304 22584
rect 3988 22030 4016 22578
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3884 21888 3936 21894
rect 3884 21830 3936 21836
rect 3896 20398 3924 21830
rect 4356 21690 4384 23054
rect 5000 22778 5028 23054
rect 4988 22772 5040 22778
rect 4988 22714 5040 22720
rect 4492 22332 4800 22341
rect 4492 22330 4498 22332
rect 4554 22330 4578 22332
rect 4634 22330 4658 22332
rect 4714 22330 4738 22332
rect 4794 22330 4800 22332
rect 4554 22278 4556 22330
rect 4736 22278 4738 22330
rect 4492 22276 4498 22278
rect 4554 22276 4578 22278
rect 4634 22276 4658 22278
rect 4714 22276 4738 22278
rect 4794 22276 4800 22278
rect 4492 22267 4800 22276
rect 4344 21684 4396 21690
rect 4344 21626 4396 21632
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 4172 20330 4200 21490
rect 4356 20534 4384 21490
rect 4492 21244 4800 21253
rect 4492 21242 4498 21244
rect 4554 21242 4578 21244
rect 4634 21242 4658 21244
rect 4714 21242 4738 21244
rect 4794 21242 4800 21244
rect 4554 21190 4556 21242
rect 4736 21190 4738 21242
rect 4492 21188 4498 21190
rect 4554 21188 4578 21190
rect 4634 21188 4658 21190
rect 4714 21188 4738 21190
rect 4794 21188 4800 21190
rect 4492 21179 4800 21188
rect 4344 20528 4396 20534
rect 4344 20470 4396 20476
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3884 19780 3936 19786
rect 3884 19722 3936 19728
rect 3896 19378 3924 19722
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3988 16182 4016 20198
rect 4172 20074 4200 20266
rect 4080 20046 4200 20074
rect 4080 19854 4108 20046
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 4080 19718 4108 19790
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4080 19378 4108 19654
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4172 17814 4200 19926
rect 4264 19854 4292 20402
rect 4492 20156 4800 20165
rect 4492 20154 4498 20156
rect 4554 20154 4578 20156
rect 4634 20154 4658 20156
rect 4714 20154 4738 20156
rect 4794 20154 4800 20156
rect 4554 20102 4556 20154
rect 4736 20102 4738 20154
rect 4492 20100 4498 20102
rect 4554 20100 4578 20102
rect 4634 20100 4658 20102
rect 4714 20100 4738 20102
rect 4794 20100 4800 20102
rect 4492 20091 4800 20100
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4264 19446 4292 19790
rect 4448 19514 4476 19790
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4724 19514 4752 19654
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4252 19440 4304 19446
rect 4252 19382 4304 19388
rect 4492 19068 4800 19077
rect 4492 19066 4498 19068
rect 4554 19066 4578 19068
rect 4634 19066 4658 19068
rect 4714 19066 4738 19068
rect 4794 19066 4800 19068
rect 4554 19014 4556 19066
rect 4736 19014 4738 19066
rect 4492 19012 4498 19014
rect 4554 19012 4578 19014
rect 4634 19012 4658 19014
rect 4714 19012 4738 19014
rect 4794 19012 4800 19014
rect 4492 19003 4800 19012
rect 5184 18358 5212 24890
rect 5276 24818 5304 25230
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5276 19514 5304 19790
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5368 18970 5396 26250
rect 5552 25770 5580 26318
rect 5632 25900 5684 25906
rect 5632 25842 5684 25848
rect 5540 25764 5592 25770
rect 5540 25706 5592 25712
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5552 24206 5580 24550
rect 5644 24342 5672 25842
rect 5632 24336 5684 24342
rect 5632 24278 5684 24284
rect 5540 24200 5592 24206
rect 5540 24142 5592 24148
rect 5736 19718 5764 26318
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5552 18630 5580 18838
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 4988 18352 5040 18358
rect 4988 18294 5040 18300
rect 5172 18352 5224 18358
rect 5172 18294 5224 18300
rect 5000 18154 5028 18294
rect 4988 18148 5040 18154
rect 4988 18090 5040 18096
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4356 17660 4384 18022
rect 4492 17980 4800 17989
rect 4492 17978 4498 17980
rect 4554 17978 4578 17980
rect 4634 17978 4658 17980
rect 4714 17978 4738 17980
rect 4794 17978 4800 17980
rect 4554 17926 4556 17978
rect 4736 17926 4738 17978
rect 4492 17924 4498 17926
rect 4554 17924 4578 17926
rect 4634 17924 4658 17926
rect 4714 17924 4738 17926
rect 4794 17924 4800 17926
rect 4492 17915 4800 17924
rect 4436 17672 4488 17678
rect 4356 17632 4436 17660
rect 4436 17614 4488 17620
rect 5000 17338 5028 18090
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5276 17814 5304 18022
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5172 17604 5224 17610
rect 5172 17546 5224 17552
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4492 16892 4800 16901
rect 4492 16890 4498 16892
rect 4554 16890 4578 16892
rect 4634 16890 4658 16892
rect 4714 16890 4738 16892
rect 4794 16890 4800 16892
rect 4554 16838 4556 16890
rect 4736 16838 4738 16890
rect 4492 16836 4498 16838
rect 4554 16836 4578 16838
rect 4634 16836 4658 16838
rect 4714 16836 4738 16838
rect 4794 16836 4800 16838
rect 4492 16827 4800 16836
rect 5184 16794 5212 17546
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3804 15502 3832 16118
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3988 15434 4016 16118
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4080 15502 4108 16050
rect 5276 15994 5304 17750
rect 5184 15966 5304 15994
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 4492 15804 4800 15813
rect 4492 15802 4498 15804
rect 4554 15802 4578 15804
rect 4634 15802 4658 15804
rect 4714 15802 4738 15804
rect 4794 15802 4800 15804
rect 4554 15750 4556 15802
rect 4736 15750 4738 15802
rect 4492 15748 4498 15750
rect 4554 15748 4578 15750
rect 4634 15748 4658 15750
rect 4714 15748 4738 15750
rect 4794 15748 4800 15750
rect 4492 15739 4800 15748
rect 5184 15706 5212 15966
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3976 15428 4028 15434
rect 3976 15370 4028 15376
rect 4080 15162 4108 15438
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4356 14618 4384 14962
rect 4632 14822 4660 15642
rect 5172 15428 5224 15434
rect 5172 15370 5224 15376
rect 5184 15094 5212 15370
rect 5172 15088 5224 15094
rect 5172 15030 5224 15036
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4492 14716 4800 14725
rect 4492 14714 4498 14716
rect 4554 14714 4578 14716
rect 4634 14714 4658 14716
rect 4714 14714 4738 14716
rect 4794 14714 4800 14716
rect 4554 14662 4556 14714
rect 4736 14662 4738 14714
rect 4492 14660 4498 14662
rect 4554 14660 4578 14662
rect 4634 14660 4658 14662
rect 4714 14660 4738 14662
rect 4794 14660 4800 14662
rect 4492 14651 4800 14660
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4908 14414 4936 14894
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4264 12170 4292 14214
rect 4540 14006 4568 14350
rect 4632 14074 4660 14350
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4492 13628 4800 13637
rect 4492 13626 4498 13628
rect 4554 13626 4578 13628
rect 4634 13626 4658 13628
rect 4714 13626 4738 13628
rect 4794 13626 4800 13628
rect 4554 13574 4556 13626
rect 4736 13574 4738 13626
rect 4492 13572 4498 13574
rect 4554 13572 4578 13574
rect 4634 13572 4658 13574
rect 4714 13572 4738 13574
rect 4794 13572 4800 13574
rect 4492 13563 4800 13572
rect 4492 12540 4800 12549
rect 4492 12538 4498 12540
rect 4554 12538 4578 12540
rect 4634 12538 4658 12540
rect 4714 12538 4738 12540
rect 4794 12538 4800 12540
rect 4554 12486 4556 12538
rect 4736 12486 4738 12538
rect 4492 12484 4498 12486
rect 4554 12484 4578 12486
rect 4634 12484 4658 12486
rect 4714 12484 4738 12486
rect 4794 12484 4800 12486
rect 4492 12475 4800 12484
rect 5000 12434 5028 14554
rect 4908 12406 5028 12434
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4264 11150 4292 11494
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3160 9654 3188 10406
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3344 9586 3372 11018
rect 4264 10606 4292 11086
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2884 7834 2912 8434
rect 2976 8090 3004 9318
rect 3896 9178 3924 9590
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 4172 8566 4200 9998
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2884 7806 3004 7834
rect 2976 7750 3004 7806
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2976 4078 3004 7686
rect 3436 7313 3464 8230
rect 3422 7304 3478 7313
rect 3422 7239 3478 7248
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3988 6390 4016 6598
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 2964 4072 3016 4078
rect 2962 4040 2964 4049
rect 3016 4040 3018 4049
rect 2962 3975 3018 3984
rect 2412 3120 2464 3126
rect 2412 3062 2464 3068
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 4172 2774 4200 8502
rect 4264 6866 4292 10542
rect 4356 9586 4384 12038
rect 4724 11558 4752 12310
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4492 11452 4800 11461
rect 4492 11450 4498 11452
rect 4554 11450 4578 11452
rect 4634 11450 4658 11452
rect 4714 11450 4738 11452
rect 4794 11450 4800 11452
rect 4554 11398 4556 11450
rect 4736 11398 4738 11450
rect 4492 11396 4498 11398
rect 4554 11396 4578 11398
rect 4634 11396 4658 11398
rect 4714 11396 4738 11398
rect 4794 11396 4800 11398
rect 4492 11387 4800 11396
rect 4908 11218 4936 12406
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5000 11762 5028 12242
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4724 10606 4752 11018
rect 4816 10606 4844 11086
rect 4908 10674 4936 11154
rect 5092 11082 5120 14758
rect 5184 11150 5212 15030
rect 5276 14822 5304 15846
rect 5552 15162 5580 15982
rect 5644 15706 5672 18770
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5736 17678 5764 18566
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5828 17134 5856 28970
rect 6748 28762 6776 29106
rect 7852 28762 7880 30194
rect 9048 30122 9076 31965
rect 11336 30252 11388 30258
rect 11336 30194 11388 30200
rect 9036 30116 9088 30122
rect 9036 30058 9088 30064
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 8760 29504 8812 29510
rect 8760 29446 8812 29452
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 8034 29404 8342 29413
rect 8034 29402 8040 29404
rect 8096 29402 8120 29404
rect 8176 29402 8200 29404
rect 8256 29402 8280 29404
rect 8336 29402 8342 29404
rect 8096 29350 8098 29402
rect 8278 29350 8280 29402
rect 8034 29348 8040 29350
rect 8096 29348 8120 29350
rect 8176 29348 8200 29350
rect 8256 29348 8280 29350
rect 8336 29348 8342 29350
rect 8034 29339 8342 29348
rect 8668 29232 8720 29238
rect 8668 29174 8720 29180
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 6736 28756 6788 28762
rect 6736 28698 6788 28704
rect 7840 28756 7892 28762
rect 7840 28698 7892 28704
rect 7104 28552 7156 28558
rect 7104 28494 7156 28500
rect 6644 28416 6696 28422
rect 6644 28358 6696 28364
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6472 23730 6500 25094
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 6184 23724 6236 23730
rect 6184 23666 6236 23672
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6196 23322 6224 23666
rect 6276 23656 6328 23662
rect 6276 23598 6328 23604
rect 6184 23316 6236 23322
rect 6184 23258 6236 23264
rect 6288 23050 6316 23598
rect 6472 23050 6500 23666
rect 6564 23118 6592 23802
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 6276 23044 6328 23050
rect 6276 22986 6328 22992
rect 6460 23044 6512 23050
rect 6460 22986 6512 22992
rect 6472 22710 6500 22986
rect 6564 22778 6592 23054
rect 6552 22772 6604 22778
rect 6552 22714 6604 22720
rect 6460 22704 6512 22710
rect 6460 22646 6512 22652
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6564 20806 6592 21966
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 5908 20460 5960 20466
rect 5908 20402 5960 20408
rect 5920 20058 5948 20402
rect 6460 20256 6512 20262
rect 6460 20198 6512 20204
rect 5908 20052 5960 20058
rect 5908 19994 5960 20000
rect 6472 19990 6500 20198
rect 6564 20058 6592 20742
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 6460 19984 6512 19990
rect 6460 19926 6512 19932
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 5920 18766 5948 19314
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6196 18766 6224 19110
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6564 17678 6592 17750
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 6380 16998 6408 17614
rect 6564 17066 6592 17614
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5644 15094 5672 15642
rect 5632 15088 5684 15094
rect 5460 15036 5632 15042
rect 5460 15030 5684 15036
rect 5460 15014 5672 15030
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5368 14498 5396 14826
rect 5276 14470 5396 14498
rect 5276 14414 5304 14470
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5276 14074 5304 14350
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5276 11898 5304 12174
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5460 10742 5488 15014
rect 5828 13938 5856 16934
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 15570 6224 15846
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6472 14414 6500 15438
rect 6656 14414 6684 28358
rect 7116 26586 7144 28494
rect 7852 28218 7880 28698
rect 8312 28490 8340 29106
rect 8392 29096 8444 29102
rect 8392 29038 8444 29044
rect 8404 28762 8432 29038
rect 8392 28756 8444 28762
rect 8392 28698 8444 28704
rect 8680 28694 8708 29174
rect 8772 29170 8800 29446
rect 8760 29164 8812 29170
rect 8760 29106 8812 29112
rect 9312 29028 9364 29034
rect 9312 28970 9364 28976
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 8668 28688 8720 28694
rect 8668 28630 8720 28636
rect 9140 28626 9168 28902
rect 9128 28620 9180 28626
rect 9128 28562 9180 28568
rect 9324 28558 9352 28970
rect 8944 28552 8996 28558
rect 8944 28494 8996 28500
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 8300 28484 8352 28490
rect 8300 28426 8352 28432
rect 8034 28316 8342 28325
rect 8034 28314 8040 28316
rect 8096 28314 8120 28316
rect 8176 28314 8200 28316
rect 8256 28314 8280 28316
rect 8336 28314 8342 28316
rect 8096 28262 8098 28314
rect 8278 28262 8280 28314
rect 8034 28260 8040 28262
rect 8096 28260 8120 28262
rect 8176 28260 8200 28262
rect 8256 28260 8280 28262
rect 8336 28260 8342 28262
rect 8034 28251 8342 28260
rect 8956 28218 8984 28494
rect 9220 28484 9272 28490
rect 9220 28426 9272 28432
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 8944 28212 8996 28218
rect 8944 28154 8996 28160
rect 7656 28076 7708 28082
rect 7656 28018 7708 28024
rect 7668 27130 7696 28018
rect 9232 28014 9260 28426
rect 9416 28404 9444 29446
rect 10140 29096 10192 29102
rect 10140 29038 10192 29044
rect 10152 28422 10180 29038
rect 10980 28994 11008 29990
rect 11348 29510 11376 30194
rect 11624 30122 11652 31965
rect 13556 30326 13584 31965
rect 15118 30492 15426 30501
rect 15118 30490 15124 30492
rect 15180 30490 15204 30492
rect 15260 30490 15284 30492
rect 15340 30490 15364 30492
rect 15420 30490 15426 30492
rect 15180 30438 15182 30490
rect 15362 30438 15364 30490
rect 15118 30436 15124 30438
rect 15180 30436 15204 30438
rect 15260 30436 15284 30438
rect 15340 30436 15364 30438
rect 15420 30436 15426 30438
rect 15118 30427 15426 30436
rect 15488 30326 15516 31965
rect 13544 30320 13596 30326
rect 13544 30262 13596 30268
rect 15476 30320 15528 30326
rect 15476 30262 15528 30268
rect 18064 30258 18092 31965
rect 19996 30258 20024 31965
rect 21928 30258 21956 31965
rect 22202 30492 22510 30501
rect 22202 30490 22208 30492
rect 22264 30490 22288 30492
rect 22344 30490 22368 30492
rect 22424 30490 22448 30492
rect 22504 30490 22510 30492
rect 22264 30438 22266 30490
rect 22446 30438 22448 30490
rect 22202 30436 22208 30438
rect 22264 30436 22288 30438
rect 22344 30436 22368 30438
rect 22424 30436 22448 30438
rect 22504 30436 22510 30438
rect 22202 30427 22510 30436
rect 24504 30258 24532 31965
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 19984 30252 20036 30258
rect 19984 30194 20036 30200
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 24492 30252 24544 30258
rect 24492 30194 24544 30200
rect 26332 30252 26384 30258
rect 26332 30194 26384 30200
rect 13912 30184 13964 30190
rect 13912 30126 13964 30132
rect 11612 30116 11664 30122
rect 11612 30058 11664 30064
rect 13084 30116 13136 30122
rect 13360 30116 13412 30122
rect 13136 30076 13360 30104
rect 13084 30058 13136 30064
rect 13360 30058 13412 30064
rect 11576 29948 11884 29957
rect 11576 29946 11582 29948
rect 11638 29946 11662 29948
rect 11718 29946 11742 29948
rect 11798 29946 11822 29948
rect 11878 29946 11884 29948
rect 11638 29894 11640 29946
rect 11820 29894 11822 29946
rect 11576 29892 11582 29894
rect 11638 29892 11662 29894
rect 11718 29892 11742 29894
rect 11798 29892 11822 29894
rect 11878 29892 11884 29894
rect 11576 29883 11884 29892
rect 13360 29776 13412 29782
rect 13360 29718 13412 29724
rect 12992 29708 13044 29714
rect 12992 29650 13044 29656
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 11336 29504 11388 29510
rect 11336 29446 11388 29452
rect 10980 28966 11100 28994
rect 10232 28960 10284 28966
rect 10232 28902 10284 28908
rect 10244 28762 10272 28902
rect 10232 28756 10284 28762
rect 10232 28698 10284 28704
rect 9324 28376 9444 28404
rect 10140 28416 10192 28422
rect 9324 28082 9352 28376
rect 10140 28358 10192 28364
rect 9312 28076 9364 28082
rect 9312 28018 9364 28024
rect 9220 28008 9272 28014
rect 9220 27950 9272 27956
rect 7748 27940 7800 27946
rect 7748 27882 7800 27888
rect 7656 27124 7708 27130
rect 7656 27066 7708 27072
rect 7760 27010 7788 27882
rect 8392 27328 8444 27334
rect 9324 27316 9352 28018
rect 10152 27878 10180 28358
rect 10244 28218 10272 28698
rect 10232 28212 10284 28218
rect 10232 28154 10284 28160
rect 10692 28008 10744 28014
rect 10692 27950 10744 27956
rect 10140 27872 10192 27878
rect 10140 27814 10192 27820
rect 10048 27532 10100 27538
rect 10048 27474 10100 27480
rect 9404 27328 9456 27334
rect 9324 27288 9404 27316
rect 8392 27270 8444 27276
rect 9404 27270 9456 27276
rect 8034 27228 8342 27237
rect 8034 27226 8040 27228
rect 8096 27226 8120 27228
rect 8176 27226 8200 27228
rect 8256 27226 8280 27228
rect 8336 27226 8342 27228
rect 8096 27174 8098 27226
rect 8278 27174 8280 27226
rect 8034 27172 8040 27174
rect 8096 27172 8120 27174
rect 8176 27172 8200 27174
rect 8256 27172 8280 27174
rect 8336 27172 8342 27174
rect 8034 27163 8342 27172
rect 7668 26982 7788 27010
rect 7196 26920 7248 26926
rect 7196 26862 7248 26868
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 7012 26376 7064 26382
rect 7012 26318 7064 26324
rect 7024 26042 7052 26318
rect 7208 26042 7236 26862
rect 7012 26036 7064 26042
rect 7012 25978 7064 25984
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 7196 25900 7248 25906
rect 7196 25842 7248 25848
rect 6736 25832 6788 25838
rect 6736 25774 6788 25780
rect 6748 25158 6776 25774
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 6840 25294 6868 25638
rect 7024 25498 7052 25842
rect 7012 25492 7064 25498
rect 7012 25434 7064 25440
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 7208 25226 7236 25842
rect 7196 25220 7248 25226
rect 7196 25162 7248 25168
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 7208 24614 7236 25162
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6840 23730 6868 24006
rect 6828 23724 6880 23730
rect 6828 23666 6880 23672
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 7024 22098 7052 22918
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6932 19514 6960 20198
rect 7024 20058 7052 20334
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 7024 19786 7052 19994
rect 7116 19854 7144 20402
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6932 17338 6960 18362
rect 7024 17882 7052 18702
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 7116 17762 7144 19246
rect 7024 17734 7144 17762
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7024 16794 7052 17734
rect 7208 17626 7236 24550
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 7300 20398 7328 22578
rect 7392 21962 7420 23054
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7380 21956 7432 21962
rect 7380 21898 7432 21904
rect 7484 20466 7512 22918
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7576 22166 7604 22578
rect 7564 22160 7616 22166
rect 7564 22102 7616 22108
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7392 19854 7420 20334
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 19174 7328 19654
rect 7392 19310 7420 19790
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7300 18358 7328 19110
rect 7484 18970 7512 19722
rect 7668 19446 7696 26982
rect 8300 26784 8352 26790
rect 8300 26726 8352 26732
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7760 25362 7788 26522
rect 8312 26450 8340 26726
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8404 26382 8432 27270
rect 8944 26988 8996 26994
rect 8944 26930 8996 26936
rect 8760 26852 8812 26858
rect 8760 26794 8812 26800
rect 8484 26444 8536 26450
rect 8484 26386 8536 26392
rect 8392 26376 8444 26382
rect 8298 26344 8354 26353
rect 8392 26318 8444 26324
rect 8298 26279 8354 26288
rect 8312 26246 8340 26279
rect 7840 26240 7892 26246
rect 7840 26182 7892 26188
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 7852 25906 7880 26182
rect 8034 26140 8342 26149
rect 8034 26138 8040 26140
rect 8096 26138 8120 26140
rect 8176 26138 8200 26140
rect 8256 26138 8280 26140
rect 8336 26138 8342 26140
rect 8096 26086 8098 26138
rect 8278 26086 8280 26138
rect 8034 26084 8040 26086
rect 8096 26084 8120 26086
rect 8176 26084 8200 26086
rect 8256 26084 8280 26086
rect 8336 26084 8342 26086
rect 8034 26075 8342 26084
rect 8404 25906 8432 26318
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 7748 25356 7800 25362
rect 7748 25298 7800 25304
rect 7760 24818 7788 25298
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 7852 24886 7880 25230
rect 7944 24954 7972 25842
rect 8208 25764 8260 25770
rect 8208 25706 8260 25712
rect 8220 25498 8248 25706
rect 8208 25492 8260 25498
rect 8208 25434 8260 25440
rect 8034 25052 8342 25061
rect 8034 25050 8040 25052
rect 8096 25050 8120 25052
rect 8176 25050 8200 25052
rect 8256 25050 8280 25052
rect 8336 25050 8342 25052
rect 8096 24998 8098 25050
rect 8278 24998 8280 25050
rect 8034 24996 8040 24998
rect 8096 24996 8120 24998
rect 8176 24996 8200 24998
rect 8256 24996 8280 24998
rect 8336 24996 8342 24998
rect 8034 24987 8342 24996
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 7840 24880 7892 24886
rect 7840 24822 7892 24828
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 7760 23186 7788 24754
rect 8220 24070 8248 24754
rect 8208 24064 8260 24070
rect 8208 24006 8260 24012
rect 8034 23964 8342 23973
rect 8034 23962 8040 23964
rect 8096 23962 8120 23964
rect 8176 23962 8200 23964
rect 8256 23962 8280 23964
rect 8336 23962 8342 23964
rect 8096 23910 8098 23962
rect 8278 23910 8280 23962
rect 8034 23908 8040 23910
rect 8096 23908 8120 23910
rect 8176 23908 8200 23910
rect 8256 23908 8280 23910
rect 8336 23908 8342 23910
rect 8034 23899 8342 23908
rect 8116 23792 8168 23798
rect 8116 23734 8168 23740
rect 7748 23180 7800 23186
rect 7748 23122 7800 23128
rect 8128 23118 8156 23734
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8034 22876 8342 22885
rect 8034 22874 8040 22876
rect 8096 22874 8120 22876
rect 8176 22874 8200 22876
rect 8256 22874 8280 22876
rect 8336 22874 8342 22876
rect 8096 22822 8098 22874
rect 8278 22822 8280 22874
rect 8034 22820 8040 22822
rect 8096 22820 8120 22822
rect 8176 22820 8200 22822
rect 8256 22820 8280 22822
rect 8336 22820 8342 22822
rect 8034 22811 8342 22820
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7852 21026 7880 21966
rect 8220 21962 8248 22374
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8034 21788 8342 21797
rect 8034 21786 8040 21788
rect 8096 21786 8120 21788
rect 8176 21786 8200 21788
rect 8256 21786 8280 21788
rect 8336 21786 8342 21788
rect 8096 21734 8098 21786
rect 8278 21734 8280 21786
rect 8034 21732 8040 21734
rect 8096 21732 8120 21734
rect 8176 21732 8200 21734
rect 8256 21732 8280 21734
rect 8336 21732 8342 21734
rect 8034 21723 8342 21732
rect 7852 20998 7972 21026
rect 7944 20806 7972 20998
rect 7932 20800 7984 20806
rect 7932 20742 7984 20748
rect 7944 20584 7972 20742
rect 8034 20700 8342 20709
rect 8034 20698 8040 20700
rect 8096 20698 8120 20700
rect 8176 20698 8200 20700
rect 8256 20698 8280 20700
rect 8336 20698 8342 20700
rect 8096 20646 8098 20698
rect 8278 20646 8280 20698
rect 8034 20644 8040 20646
rect 8096 20644 8120 20646
rect 8176 20644 8200 20646
rect 8256 20644 8280 20646
rect 8336 20644 8342 20646
rect 8034 20635 8342 20644
rect 8300 20596 8352 20602
rect 7760 20556 8156 20584
rect 7656 19440 7708 19446
rect 7656 19382 7708 19388
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7300 17746 7328 18294
rect 7484 18290 7512 18906
rect 7668 18290 7696 19110
rect 7760 18902 7788 20556
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7944 20262 7972 20334
rect 8128 20262 8156 20556
rect 8300 20538 8352 20544
rect 8312 20466 8340 20538
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 7748 18896 7800 18902
rect 7748 18838 7800 18844
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7484 17678 7512 18226
rect 7668 17678 7696 18226
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7760 17746 7788 18022
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7116 17610 7236 17626
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7104 17604 7236 17610
rect 7156 17598 7236 17604
rect 7104 17546 7156 17552
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6920 16108 6972 16114
rect 7024 16096 7052 16730
rect 6972 16068 7052 16096
rect 6920 16050 6972 16056
rect 6748 15162 6776 16050
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 6000 12912 6052 12918
rect 6000 12854 6052 12860
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12238 5948 12582
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5828 11898 5856 12174
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5644 10810 5672 11222
rect 6012 10810 6040 12854
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4492 10364 4800 10373
rect 4492 10362 4498 10364
rect 4554 10362 4578 10364
rect 4634 10362 4658 10364
rect 4714 10362 4738 10364
rect 4794 10362 4800 10364
rect 4554 10310 4556 10362
rect 4736 10310 4738 10362
rect 4492 10308 4498 10310
rect 4554 10308 4578 10310
rect 4634 10308 4658 10310
rect 4714 10308 4738 10310
rect 4794 10308 4800 10310
rect 4492 10299 4800 10308
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 8974 4384 9318
rect 4492 9276 4800 9285
rect 4492 9274 4498 9276
rect 4554 9274 4578 9276
rect 4634 9274 4658 9276
rect 4714 9274 4738 9276
rect 4794 9274 4800 9276
rect 4554 9222 4556 9274
rect 4736 9222 4738 9274
rect 4492 9220 4498 9222
rect 4554 9220 4578 9222
rect 4634 9220 4658 9222
rect 4714 9220 4738 9222
rect 4794 9220 4800 9222
rect 4492 9211 4800 9220
rect 4908 9042 4936 10406
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4632 8294 4660 8774
rect 4816 8430 4844 8910
rect 4908 8566 4936 8978
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 5000 8634 5028 8774
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4804 8424 4856 8430
rect 4856 8372 4936 8378
rect 4804 8366 4936 8372
rect 4816 8350 4936 8366
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4492 8188 4800 8197
rect 4492 8186 4498 8188
rect 4554 8186 4578 8188
rect 4634 8186 4658 8188
rect 4714 8186 4738 8188
rect 4794 8186 4800 8188
rect 4554 8134 4556 8186
rect 4736 8134 4738 8186
rect 4492 8132 4498 8134
rect 4554 8132 4578 8134
rect 4634 8132 4658 8134
rect 4714 8132 4738 8134
rect 4794 8132 4800 8134
rect 4492 8123 4800 8132
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4632 7342 4660 7822
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4492 7100 4800 7109
rect 4492 7098 4498 7100
rect 4554 7098 4578 7100
rect 4634 7098 4658 7100
rect 4714 7098 4738 7100
rect 4794 7098 4800 7100
rect 4554 7046 4556 7098
rect 4736 7046 4738 7098
rect 4492 7044 4498 7046
rect 4554 7044 4578 7046
rect 4634 7044 4658 7046
rect 4714 7044 4738 7046
rect 4794 7044 4800 7046
rect 4492 7035 4800 7044
rect 4908 7002 4936 8350
rect 5000 8022 5028 8570
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5000 7410 5028 7822
rect 5092 7750 5120 9114
rect 5368 8514 5396 10542
rect 5460 8906 5488 10678
rect 5644 8974 5672 10746
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5460 8634 5488 8842
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5368 8486 5488 8514
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5276 8294 5304 8366
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 5092 7342 5120 7686
rect 5184 7342 5212 7958
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4896 6792 4948 6798
rect 5000 6780 5028 7210
rect 5276 6798 5304 8230
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5368 7546 5396 7958
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 4948 6752 5028 6780
rect 5264 6792 5316 6798
rect 4896 6734 4948 6740
rect 5264 6734 5316 6740
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4356 4826 4384 6054
rect 4492 6012 4800 6021
rect 4492 6010 4498 6012
rect 4554 6010 4578 6012
rect 4634 6010 4658 6012
rect 4714 6010 4738 6012
rect 4794 6010 4800 6012
rect 4554 5958 4556 6010
rect 4736 5958 4738 6010
rect 4492 5956 4498 5958
rect 4554 5956 4578 5958
rect 4634 5956 4658 5958
rect 4714 5956 4738 5958
rect 4794 5956 4800 5958
rect 4492 5947 4800 5956
rect 4908 5846 4936 6734
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6322 5396 6598
rect 5460 6458 5488 8486
rect 5644 8430 5672 8910
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5736 7954 5764 8502
rect 6196 8090 6224 14214
rect 6840 13938 6868 14486
rect 6932 14006 6960 14554
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6840 13190 6868 13874
rect 7024 13394 7052 16068
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7484 15094 7512 15914
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7116 14414 7144 14962
rect 7484 14498 7512 15030
rect 7576 14890 7604 17478
rect 7760 17218 7788 17682
rect 7668 17202 7788 17218
rect 7656 17196 7788 17202
rect 7708 17190 7788 17196
rect 7656 17138 7708 17144
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7654 16008 7710 16017
rect 7760 15978 7788 16050
rect 7852 16017 7880 19926
rect 7944 19174 7972 20198
rect 8312 20058 8340 20402
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8312 19700 8340 19994
rect 8312 19672 8432 19700
rect 8034 19612 8342 19621
rect 8034 19610 8040 19612
rect 8096 19610 8120 19612
rect 8176 19610 8200 19612
rect 8256 19610 8280 19612
rect 8336 19610 8342 19612
rect 8096 19558 8098 19610
rect 8278 19558 8280 19610
rect 8034 19556 8040 19558
rect 8096 19556 8120 19558
rect 8176 19556 8200 19558
rect 8256 19556 8280 19558
rect 8336 19556 8342 19558
rect 8034 19547 8342 19556
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8220 18766 8248 19110
rect 8404 18970 8432 19672
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8034 18524 8342 18533
rect 8034 18522 8040 18524
rect 8096 18522 8120 18524
rect 8176 18522 8200 18524
rect 8256 18522 8280 18524
rect 8336 18522 8342 18524
rect 8096 18470 8098 18522
rect 8278 18470 8280 18522
rect 8034 18468 8040 18470
rect 8096 18468 8120 18470
rect 8176 18468 8200 18470
rect 8256 18468 8280 18470
rect 8336 18468 8342 18470
rect 8034 18459 8342 18468
rect 8404 18426 8432 18906
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8404 17610 8432 18226
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17134 7972 17478
rect 8034 17436 8342 17445
rect 8034 17434 8040 17436
rect 8096 17434 8120 17436
rect 8176 17434 8200 17436
rect 8256 17434 8280 17436
rect 8336 17434 8342 17436
rect 8096 17382 8098 17434
rect 8278 17382 8280 17434
rect 8034 17380 8040 17382
rect 8096 17380 8120 17382
rect 8176 17380 8200 17382
rect 8256 17380 8280 17382
rect 8336 17380 8342 17382
rect 8034 17371 8342 17380
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 8404 16794 8432 17546
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8034 16348 8342 16357
rect 8034 16346 8040 16348
rect 8096 16346 8120 16348
rect 8176 16346 8200 16348
rect 8256 16346 8280 16348
rect 8336 16346 8342 16348
rect 8096 16294 8098 16346
rect 8278 16294 8280 16346
rect 8034 16292 8040 16294
rect 8096 16292 8120 16294
rect 8176 16292 8200 16294
rect 8256 16292 8280 16294
rect 8336 16292 8342 16294
rect 8034 16283 8342 16292
rect 7838 16008 7894 16017
rect 7654 15943 7656 15952
rect 7708 15943 7710 15952
rect 7748 15972 7800 15978
rect 7656 15914 7708 15920
rect 7838 15943 7894 15952
rect 7748 15914 7800 15920
rect 8034 15260 8342 15269
rect 8034 15258 8040 15260
rect 8096 15258 8120 15260
rect 8176 15258 8200 15260
rect 8256 15258 8280 15260
rect 8336 15258 8342 15260
rect 8096 15206 8098 15258
rect 8278 15206 8280 15258
rect 8034 15204 8040 15206
rect 8096 15204 8120 15206
rect 8176 15204 8200 15206
rect 8256 15204 8280 15206
rect 8336 15204 8342 15206
rect 8034 15195 8342 15204
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7576 14618 7604 14826
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7392 14470 7512 14498
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6920 12844 6972 12850
rect 7288 12844 7340 12850
rect 6972 12804 7288 12832
rect 6920 12786 6972 12792
rect 7288 12786 7340 12792
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 7024 12170 7052 12650
rect 7392 12238 7420 14470
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7564 14000 7616 14006
rect 7562 13968 7564 13977
rect 7616 13968 7618 13977
rect 7562 13903 7618 13912
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7484 12986 7512 13262
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7852 12714 7880 14214
rect 8034 14172 8342 14181
rect 8034 14170 8040 14172
rect 8096 14170 8120 14172
rect 8176 14170 8200 14172
rect 8256 14170 8280 14172
rect 8336 14170 8342 14172
rect 8096 14118 8098 14170
rect 8278 14118 8280 14170
rect 8034 14116 8040 14118
rect 8096 14116 8120 14118
rect 8176 14116 8200 14118
rect 8256 14116 8280 14118
rect 8336 14116 8342 14118
rect 8034 14107 8342 14116
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8034 13084 8342 13093
rect 8034 13082 8040 13084
rect 8096 13082 8120 13084
rect 8176 13082 8200 13084
rect 8256 13082 8280 13084
rect 8336 13082 8342 13084
rect 8096 13030 8098 13082
rect 8278 13030 8280 13082
rect 8034 13028 8040 13030
rect 8096 13028 8120 13030
rect 8176 13028 8200 13030
rect 8256 13028 8280 13030
rect 8336 13028 8342 13030
rect 8034 13019 8342 13028
rect 8404 13002 8432 13806
rect 8496 13190 8524 26386
rect 8772 26042 8800 26794
rect 8760 26036 8812 26042
rect 8760 25978 8812 25984
rect 8668 25900 8720 25906
rect 8668 25842 8720 25848
rect 8680 25362 8708 25842
rect 8668 25356 8720 25362
rect 8668 25298 8720 25304
rect 8852 24608 8904 24614
rect 8852 24550 8904 24556
rect 8864 24206 8892 24550
rect 8852 24200 8904 24206
rect 8852 24142 8904 24148
rect 8864 23730 8892 24142
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8864 23526 8892 23666
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 8864 22710 8892 23462
rect 8852 22704 8904 22710
rect 8852 22646 8904 22652
rect 8864 22506 8892 22646
rect 8852 22500 8904 22506
rect 8852 22442 8904 22448
rect 8668 21956 8720 21962
rect 8668 21898 8720 21904
rect 8680 21690 8708 21898
rect 8956 21690 8984 26930
rect 9220 25900 9272 25906
rect 9220 25842 9272 25848
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 9048 23866 9076 24142
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 8668 21684 8720 21690
rect 8668 21626 8720 21632
rect 8944 21684 8996 21690
rect 8944 21626 8996 21632
rect 8680 21350 8708 21626
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9140 19446 9168 20402
rect 9128 19440 9180 19446
rect 9128 19382 9180 19388
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8588 18290 8616 18770
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 9232 18154 9260 25842
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 9324 24206 9352 25230
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9324 23798 9352 24142
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9416 22094 9444 27270
rect 10060 26518 10088 27474
rect 10048 26512 10100 26518
rect 10048 26454 10100 26460
rect 9864 26308 9916 26314
rect 9864 26250 9916 26256
rect 9876 26042 9904 26250
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 9496 24676 9548 24682
rect 9496 24618 9548 24624
rect 9508 23730 9536 24618
rect 10048 24608 10100 24614
rect 10048 24550 10100 24556
rect 10060 24410 10088 24550
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 9956 24132 10008 24138
rect 9956 24074 10008 24080
rect 9588 24064 9640 24070
rect 9588 24006 9640 24012
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 9324 22066 9444 22094
rect 9324 18680 9352 22066
rect 9404 21956 9456 21962
rect 9404 21898 9456 21904
rect 9416 20924 9444 21898
rect 9508 21078 9536 23666
rect 9600 23118 9628 24006
rect 9864 23724 9916 23730
rect 9968 23712 9996 24074
rect 9916 23684 9996 23712
rect 9864 23666 9916 23672
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9692 21690 9720 22714
rect 9968 22438 9996 23684
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 10060 22710 10088 22986
rect 10048 22704 10100 22710
rect 10048 22646 10100 22652
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9968 22094 9996 22374
rect 9784 22066 9996 22094
rect 10152 22094 10180 27814
rect 10704 27606 10732 27950
rect 11072 27878 11100 28966
rect 11152 28416 11204 28422
rect 11152 28358 11204 28364
rect 11060 27872 11112 27878
rect 11060 27814 11112 27820
rect 10692 27600 10744 27606
rect 10692 27542 10744 27548
rect 11072 27402 11100 27814
rect 10876 27396 10928 27402
rect 10876 27338 10928 27344
rect 11060 27396 11112 27402
rect 11060 27338 11112 27344
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 10244 26314 10272 26930
rect 10324 26852 10376 26858
rect 10324 26794 10376 26800
rect 10232 26308 10284 26314
rect 10232 26250 10284 26256
rect 10244 25770 10272 26250
rect 10232 25764 10284 25770
rect 10232 25706 10284 25712
rect 10232 24200 10284 24206
rect 10232 24142 10284 24148
rect 10244 23866 10272 24142
rect 10232 23860 10284 23866
rect 10232 23802 10284 23808
rect 10336 23118 10364 26794
rect 10888 26790 10916 27338
rect 11072 26926 11100 27338
rect 11164 27334 11192 28358
rect 11244 27464 11296 27470
rect 11244 27406 11296 27412
rect 11152 27328 11204 27334
rect 11152 27270 11204 27276
rect 11164 27130 11192 27270
rect 11152 27124 11204 27130
rect 11152 27066 11204 27072
rect 11256 27062 11284 27406
rect 11244 27056 11296 27062
rect 11244 26998 11296 27004
rect 11060 26920 11112 26926
rect 11060 26862 11112 26868
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10888 26450 10916 26726
rect 11256 26450 11284 26998
rect 10876 26444 10928 26450
rect 10876 26386 10928 26392
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 10508 26376 10560 26382
rect 10508 26318 10560 26324
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 10428 25945 10456 26182
rect 10520 26042 10548 26318
rect 10508 26036 10560 26042
rect 10508 25978 10560 25984
rect 10414 25936 10470 25945
rect 10414 25871 10416 25880
rect 10468 25871 10470 25880
rect 10416 25842 10468 25848
rect 10416 25220 10468 25226
rect 10416 25162 10468 25168
rect 10428 24138 10456 25162
rect 10416 24132 10468 24138
rect 10416 24074 10468 24080
rect 10520 23866 10548 25978
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 10876 25152 10928 25158
rect 10876 25094 10928 25100
rect 10888 24954 10916 25094
rect 10876 24948 10928 24954
rect 10876 24890 10928 24896
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 10508 23860 10560 23866
rect 10508 23802 10560 23808
rect 10324 23112 10376 23118
rect 10324 23054 10376 23060
rect 10336 22778 10364 23054
rect 10416 22976 10468 22982
rect 10416 22918 10468 22924
rect 10428 22778 10456 22918
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10416 22772 10468 22778
rect 10416 22714 10468 22720
rect 10152 22066 10272 22094
rect 9784 21894 9812 22066
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9588 21412 9640 21418
rect 9588 21354 9640 21360
rect 9496 21072 9548 21078
rect 9496 21014 9548 21020
rect 9496 20936 9548 20942
rect 9416 20896 9496 20924
rect 9496 20878 9548 20884
rect 9508 19836 9536 20878
rect 9600 19990 9628 21354
rect 9692 21146 9720 21490
rect 9784 21418 9812 21830
rect 9772 21412 9824 21418
rect 9772 21354 9824 21360
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9784 20602 9812 21354
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9588 19984 9640 19990
rect 9588 19926 9640 19932
rect 9876 19922 9904 21966
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9968 20058 9996 20198
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9864 19916 9916 19922
rect 9784 19876 9864 19904
rect 9508 19808 9628 19836
rect 9404 19440 9456 19446
rect 9404 19382 9456 19388
rect 9416 18748 9444 19382
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9508 18970 9536 19314
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9600 18850 9628 19808
rect 9784 18970 9812 19876
rect 9864 19858 9916 19864
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9876 19378 9904 19722
rect 10060 19514 10088 21558
rect 10152 20942 10180 21830
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9600 18822 9812 18850
rect 9496 18760 9548 18766
rect 9416 18720 9496 18748
rect 9496 18702 9548 18708
rect 9324 18652 9444 18680
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8588 16658 8616 17002
rect 9048 16998 9076 17614
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9324 17270 9352 17478
rect 9312 17264 9364 17270
rect 9312 17206 9364 17212
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 9048 16250 9076 16934
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8404 12974 8524 13002
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11558 6776 12038
rect 7024 11898 7052 12106
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7484 11762 7512 12378
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 11082 6776 11494
rect 7852 11218 7880 12650
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7944 11694 7972 12038
rect 8034 11996 8342 12005
rect 8034 11994 8040 11996
rect 8096 11994 8120 11996
rect 8176 11994 8200 11996
rect 8256 11994 8280 11996
rect 8336 11994 8342 11996
rect 8096 11942 8098 11994
rect 8278 11942 8280 11994
rect 8034 11940 8040 11942
rect 8096 11940 8120 11942
rect 8176 11940 8200 11942
rect 8256 11940 8280 11942
rect 8336 11940 8342 11942
rect 8034 11931 8342 11940
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6564 8566 6592 8774
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 6458 5948 6734
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5184 5914 5212 6258
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 5920 5710 5948 6394
rect 6196 6390 6224 6598
rect 6564 6458 6592 7346
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6748 6390 6776 11018
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10130 7696 10950
rect 7852 10742 7880 11154
rect 7944 11150 7972 11630
rect 8404 11150 8432 12854
rect 8496 12850 8524 12974
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8496 11830 8524 12786
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7944 10674 7972 11086
rect 8034 10908 8342 10917
rect 8034 10906 8040 10908
rect 8096 10906 8120 10908
rect 8176 10906 8200 10908
rect 8256 10906 8280 10908
rect 8336 10906 8342 10908
rect 8096 10854 8098 10906
rect 8278 10854 8280 10906
rect 8034 10852 8040 10854
rect 8096 10852 8120 10854
rect 8176 10852 8200 10854
rect 8256 10852 8280 10854
rect 8336 10852 8342 10854
rect 8034 10843 8342 10852
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7288 9648 7340 9654
rect 7286 9616 7288 9625
rect 7340 9616 7342 9625
rect 7012 9580 7064 9586
rect 7944 9586 7972 9862
rect 8034 9820 8342 9829
rect 8034 9818 8040 9820
rect 8096 9818 8120 9820
rect 8176 9818 8200 9820
rect 8256 9818 8280 9820
rect 8336 9818 8342 9820
rect 8096 9766 8098 9818
rect 8278 9766 8280 9818
rect 8034 9764 8040 9766
rect 8096 9764 8120 9766
rect 8176 9764 8200 9766
rect 8256 9764 8280 9766
rect 8336 9764 8342 9766
rect 8034 9755 8342 9764
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 7286 9551 7342 9560
rect 7932 9580 7984 9586
rect 7012 9522 7064 9528
rect 7932 9522 7984 9528
rect 7024 9178 7052 9522
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7576 8974 7604 9318
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7564 8968 7616 8974
rect 7944 8945 7972 9386
rect 8312 9178 8340 9590
rect 8404 9586 8432 9998
rect 8588 9654 8616 13330
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8680 12782 8708 13194
rect 9048 12850 9076 13874
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8680 11880 8708 12718
rect 8864 12714 8892 12786
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8760 11892 8812 11898
rect 8680 11852 8760 11880
rect 8760 11834 8812 11840
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8680 10674 8708 11086
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 7564 8910 7616 8916
rect 7930 8936 7986 8945
rect 7208 8634 7236 8910
rect 7930 8871 7986 8880
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7944 8566 7972 8871
rect 8312 8838 8340 8978
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8034 8732 8342 8741
rect 8034 8730 8040 8732
rect 8096 8730 8120 8732
rect 8176 8730 8200 8732
rect 8256 8730 8280 8732
rect 8336 8730 8342 8732
rect 8096 8678 8098 8730
rect 8278 8678 8280 8730
rect 8034 8676 8040 8678
rect 8096 8676 8120 8678
rect 8176 8676 8200 8678
rect 8256 8676 8280 8678
rect 8336 8676 8342 8678
rect 8034 8667 8342 8676
rect 7932 8560 7984 8566
rect 7932 8502 7984 8508
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7944 7546 7972 7754
rect 8034 7644 8342 7653
rect 8034 7642 8040 7644
rect 8096 7642 8120 7644
rect 8176 7642 8200 7644
rect 8256 7642 8280 7644
rect 8336 7642 8342 7644
rect 8096 7590 8098 7642
rect 8278 7590 8280 7642
rect 8034 7588 8040 7590
rect 8096 7588 8120 7590
rect 8176 7588 8200 7590
rect 8256 7588 8280 7590
rect 8336 7588 8342 7590
rect 8034 7579 8342 7588
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7208 6798 7236 7278
rect 8404 6866 8432 9522
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 6184 6384 6236 6390
rect 6184 6326 6236 6332
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6196 6118 6224 6326
rect 7024 6322 7052 6734
rect 7208 6322 7236 6734
rect 8496 6730 8524 8774
rect 8588 8430 8616 9046
rect 8772 8634 8800 9114
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8034 6556 8342 6565
rect 8034 6554 8040 6556
rect 8096 6554 8120 6556
rect 8176 6554 8200 6556
rect 8256 6554 8280 6556
rect 8336 6554 8342 6556
rect 8096 6502 8098 6554
rect 8278 6502 8280 6554
rect 8034 6500 8040 6502
rect 8096 6500 8120 6502
rect 8176 6500 8200 6502
rect 8256 6500 8280 6502
rect 8336 6500 8342 6502
rect 8034 6491 8342 6500
rect 8496 6322 8524 6666
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5914 6224 6054
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 4492 4924 4800 4933
rect 4492 4922 4498 4924
rect 4554 4922 4578 4924
rect 4634 4922 4658 4924
rect 4714 4922 4738 4924
rect 4794 4922 4800 4924
rect 4554 4870 4556 4922
rect 4736 4870 4738 4922
rect 4492 4868 4498 4870
rect 4554 4868 4578 4870
rect 4634 4868 4658 4870
rect 4714 4868 4738 4870
rect 4794 4868 4800 4870
rect 4492 4859 4800 4868
rect 6472 4826 6500 5646
rect 6656 5370 6684 5646
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4826 6776 4966
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 4492 3836 4800 3845
rect 4492 3834 4498 3836
rect 4554 3834 4578 3836
rect 4634 3834 4658 3836
rect 4714 3834 4738 3836
rect 4794 3834 4800 3836
rect 4554 3782 4556 3834
rect 4736 3782 4738 3834
rect 4492 3780 4498 3782
rect 4554 3780 4578 3782
rect 4634 3780 4658 3782
rect 4714 3780 4738 3782
rect 4794 3780 4800 3782
rect 4492 3771 4800 3780
rect 4172 2746 4292 2774
rect 4264 2446 4292 2746
rect 4492 2748 4800 2757
rect 4492 2746 4498 2748
rect 4554 2746 4578 2748
rect 4634 2746 4658 2748
rect 4714 2746 4738 2748
rect 4794 2746 4800 2748
rect 4554 2694 4556 2746
rect 4736 2694 4738 2746
rect 4492 2692 4498 2694
rect 4554 2692 4578 2694
rect 4634 2692 4658 2694
rect 4714 2692 4738 2694
rect 4794 2692 4800 2694
rect 4492 2683 4800 2692
rect 6748 2650 6776 4762
rect 7116 4622 7144 5102
rect 7208 4690 7236 5170
rect 7852 5166 7880 5510
rect 7944 5370 7972 5646
rect 8034 5468 8342 5477
rect 8034 5466 8040 5468
rect 8096 5466 8120 5468
rect 8176 5466 8200 5468
rect 8256 5466 8280 5468
rect 8336 5466 8342 5468
rect 8096 5414 8098 5466
rect 8278 5414 8280 5466
rect 8034 5412 8040 5414
rect 8096 5412 8120 5414
rect 8176 5412 8200 5414
rect 8256 5412 8280 5414
rect 8336 5412 8342 5414
rect 8034 5403 8342 5412
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 8496 5030 8524 6258
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 8034 4380 8342 4389
rect 8034 4378 8040 4380
rect 8096 4378 8120 4380
rect 8176 4378 8200 4380
rect 8256 4378 8280 4380
rect 8336 4378 8342 4380
rect 8096 4326 8098 4378
rect 8278 4326 8280 4378
rect 8034 4324 8040 4326
rect 8096 4324 8120 4326
rect 8176 4324 8200 4326
rect 8256 4324 8280 4326
rect 8336 4324 8342 4326
rect 8034 4315 8342 4324
rect 8034 3292 8342 3301
rect 8034 3290 8040 3292
rect 8096 3290 8120 3292
rect 8176 3290 8200 3292
rect 8256 3290 8280 3292
rect 8336 3290 8342 3292
rect 8096 3238 8098 3290
rect 8278 3238 8280 3290
rect 8034 3236 8040 3238
rect 8096 3236 8120 3238
rect 8176 3236 8200 3238
rect 8256 3236 8280 3238
rect 8336 3236 8342 3238
rect 8034 3227 8342 3236
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 8588 2446 8616 8366
rect 8772 7410 8800 8570
rect 8864 7546 8892 11018
rect 9048 10674 9076 11154
rect 9140 11150 9168 14962
rect 9324 14822 9352 15302
rect 9416 14929 9444 18652
rect 9508 18426 9536 18702
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9692 17610 9720 18362
rect 9588 17604 9640 17610
rect 9588 17546 9640 17552
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9508 16794 9536 17138
rect 9600 16998 9628 17546
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9692 15706 9720 17546
rect 9784 17542 9812 18822
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9968 17678 9996 18022
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9876 16794 9904 17206
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9876 16250 9904 16458
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9692 15162 9720 15642
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9402 14920 9458 14929
rect 9402 14855 9458 14864
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14346 9352 14758
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9324 13870 9352 14282
rect 9508 13938 9536 14554
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9600 14278 9628 14418
rect 9692 14414 9720 14962
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9600 13802 9628 14214
rect 9692 14074 9720 14350
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9784 13954 9812 15030
rect 9692 13926 9812 13954
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9600 13258 9628 13738
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9692 12102 9720 13926
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9784 12238 9812 13806
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9784 11898 9812 12174
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9876 11286 9904 16186
rect 9968 13870 9996 17614
rect 10060 17270 10088 19450
rect 10244 19242 10272 22066
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10428 18426 10456 22714
rect 10520 21690 10548 23802
rect 10704 23118 10732 24006
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10796 23050 10824 23462
rect 10888 23202 10916 24890
rect 10980 23322 11008 25910
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 10888 23174 11008 23202
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10520 20942 10548 21626
rect 10612 21146 10640 21898
rect 10600 21140 10652 21146
rect 10600 21082 10652 21088
rect 10796 21078 10824 22986
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10520 20466 10548 20878
rect 10888 20874 10916 21286
rect 10876 20868 10928 20874
rect 10876 20810 10928 20816
rect 10600 20800 10652 20806
rect 10600 20742 10652 20748
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10612 19854 10640 20742
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10796 19786 10824 20198
rect 10784 19780 10836 19786
rect 10784 19722 10836 19728
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 10048 17264 10100 17270
rect 10048 17206 10100 17212
rect 10060 16794 10088 17206
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10612 16726 10640 17750
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 16998 10732 17478
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10600 16720 10652 16726
rect 10600 16662 10652 16668
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10060 16250 10088 16390
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10152 14414 10180 14758
rect 10244 14618 10272 14894
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10152 13870 10180 13942
rect 10428 13870 10456 16186
rect 10704 15502 10732 16934
rect 10796 15978 10824 19722
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10888 18086 10916 19654
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10692 15496 10744 15502
rect 10888 15473 10916 17614
rect 10980 16250 11008 23174
rect 11348 19334 11376 29446
rect 12912 29238 12940 29582
rect 13004 29306 13032 29650
rect 12992 29300 13044 29306
rect 12992 29242 13044 29248
rect 12900 29232 12952 29238
rect 12900 29174 12952 29180
rect 12624 29028 12676 29034
rect 12624 28970 12676 28976
rect 11576 28860 11884 28869
rect 11576 28858 11582 28860
rect 11638 28858 11662 28860
rect 11718 28858 11742 28860
rect 11798 28858 11822 28860
rect 11878 28858 11884 28860
rect 11638 28806 11640 28858
rect 11820 28806 11822 28858
rect 11576 28804 11582 28806
rect 11638 28804 11662 28806
rect 11718 28804 11742 28806
rect 11798 28804 11822 28806
rect 11878 28804 11884 28806
rect 11576 28795 11884 28804
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 11796 28552 11848 28558
rect 11796 28494 11848 28500
rect 11808 28082 11836 28494
rect 12164 28416 12216 28422
rect 12164 28358 12216 28364
rect 12176 28150 12204 28358
rect 12164 28144 12216 28150
rect 12164 28086 12216 28092
rect 11796 28076 11848 28082
rect 11796 28018 11848 28024
rect 11576 27772 11884 27781
rect 11576 27770 11582 27772
rect 11638 27770 11662 27772
rect 11718 27770 11742 27772
rect 11798 27770 11822 27772
rect 11878 27770 11884 27772
rect 11638 27718 11640 27770
rect 11820 27718 11822 27770
rect 11576 27716 11582 27718
rect 11638 27716 11662 27718
rect 11718 27716 11742 27718
rect 11798 27716 11822 27718
rect 11878 27716 11884 27718
rect 11576 27707 11884 27716
rect 12072 27396 12124 27402
rect 12072 27338 12124 27344
rect 11980 27056 12032 27062
rect 12084 27044 12112 27338
rect 12452 27062 12480 28562
rect 12532 28416 12584 28422
rect 12532 28358 12584 28364
rect 12032 27016 12112 27044
rect 11980 26998 12032 27004
rect 11980 26920 12032 26926
rect 11980 26862 12032 26868
rect 11576 26684 11884 26693
rect 11576 26682 11582 26684
rect 11638 26682 11662 26684
rect 11718 26682 11742 26684
rect 11798 26682 11822 26684
rect 11878 26682 11884 26684
rect 11638 26630 11640 26682
rect 11820 26630 11822 26682
rect 11576 26628 11582 26630
rect 11638 26628 11662 26630
rect 11718 26628 11742 26630
rect 11798 26628 11822 26630
rect 11878 26628 11884 26630
rect 11576 26619 11884 26628
rect 11992 26586 12020 26862
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11532 26042 11560 26318
rect 11520 26036 11572 26042
rect 11520 25978 11572 25984
rect 12084 25974 12112 27016
rect 12440 27056 12492 27062
rect 12440 26998 12492 27004
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12360 26586 12388 26930
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12360 26450 12388 26522
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12268 26246 12296 26318
rect 12256 26240 12308 26246
rect 12256 26182 12308 26188
rect 12072 25968 12124 25974
rect 11978 25936 12034 25945
rect 12072 25910 12124 25916
rect 11978 25871 12034 25880
rect 11576 25596 11884 25605
rect 11576 25594 11582 25596
rect 11638 25594 11662 25596
rect 11718 25594 11742 25596
rect 11798 25594 11822 25596
rect 11878 25594 11884 25596
rect 11638 25542 11640 25594
rect 11820 25542 11822 25594
rect 11576 25540 11582 25542
rect 11638 25540 11662 25542
rect 11718 25540 11742 25542
rect 11798 25540 11822 25542
rect 11878 25540 11884 25542
rect 11576 25531 11884 25540
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 11440 24410 11468 24686
rect 11576 24508 11884 24517
rect 11576 24506 11582 24508
rect 11638 24506 11662 24508
rect 11718 24506 11742 24508
rect 11798 24506 11822 24508
rect 11878 24506 11884 24508
rect 11638 24454 11640 24506
rect 11820 24454 11822 24506
rect 11576 24452 11582 24454
rect 11638 24452 11662 24454
rect 11718 24452 11742 24454
rect 11798 24452 11822 24454
rect 11878 24452 11884 24454
rect 11576 24443 11884 24452
rect 11428 24404 11480 24410
rect 11428 24346 11480 24352
rect 11576 23420 11884 23429
rect 11576 23418 11582 23420
rect 11638 23418 11662 23420
rect 11718 23418 11742 23420
rect 11798 23418 11822 23420
rect 11878 23418 11884 23420
rect 11638 23366 11640 23418
rect 11820 23366 11822 23418
rect 11576 23364 11582 23366
rect 11638 23364 11662 23366
rect 11718 23364 11742 23366
rect 11798 23364 11822 23366
rect 11878 23364 11884 23366
rect 11576 23355 11884 23364
rect 11992 22710 12020 25871
rect 12164 25832 12216 25838
rect 12164 25774 12216 25780
rect 12176 25294 12204 25774
rect 12268 25702 12296 26182
rect 12544 25906 12572 28358
rect 12636 27470 12664 28970
rect 12912 28558 12940 29174
rect 12992 29096 13044 29102
rect 12992 29038 13044 29044
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 13004 28422 13032 29038
rect 13372 28558 13400 29718
rect 13636 28960 13688 28966
rect 13688 28908 13860 28914
rect 13636 28902 13860 28908
rect 13648 28886 13860 28902
rect 13832 28626 13860 28886
rect 13820 28620 13872 28626
rect 13820 28562 13872 28568
rect 13360 28552 13412 28558
rect 13360 28494 13412 28500
rect 12992 28416 13044 28422
rect 12992 28358 13044 28364
rect 12900 28076 12952 28082
rect 12900 28018 12952 28024
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 12912 27674 12940 28018
rect 12900 27668 12952 27674
rect 12900 27610 12952 27616
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 13004 27130 13032 28018
rect 12992 27124 13044 27130
rect 12992 27066 13044 27072
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12728 26518 12756 26930
rect 12808 26784 12860 26790
rect 12808 26726 12860 26732
rect 12716 26512 12768 26518
rect 12716 26454 12768 26460
rect 12728 26314 12756 26454
rect 12820 26382 12848 26726
rect 12808 26376 12860 26382
rect 12808 26318 12860 26324
rect 12716 26308 12768 26314
rect 12716 26250 12768 26256
rect 12624 25968 12676 25974
rect 12624 25910 12676 25916
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 12164 25288 12216 25294
rect 12164 25230 12216 25236
rect 12268 25226 12296 25638
rect 12256 25220 12308 25226
rect 12256 25162 12308 25168
rect 12532 25152 12584 25158
rect 12636 25140 12664 25910
rect 12584 25112 12664 25140
rect 12820 25684 12848 26318
rect 13372 26042 13400 28494
rect 13728 28076 13780 28082
rect 13728 28018 13780 28024
rect 13740 27538 13768 28018
rect 13820 27872 13872 27878
rect 13820 27814 13872 27820
rect 13728 27532 13780 27538
rect 13728 27474 13780 27480
rect 13360 26036 13412 26042
rect 13360 25978 13412 25984
rect 12900 25696 12952 25702
rect 12820 25656 12900 25684
rect 12532 25094 12584 25100
rect 12544 24410 12572 25094
rect 12820 24818 12848 25656
rect 12900 25638 12952 25644
rect 13544 25288 13596 25294
rect 13544 25230 13596 25236
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12544 24138 12572 24346
rect 12716 24268 12768 24274
rect 12716 24210 12768 24216
rect 12532 24132 12584 24138
rect 12532 24074 12584 24080
rect 12728 23662 12756 24210
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 11980 22704 12032 22710
rect 11980 22646 12032 22652
rect 11576 22332 11884 22341
rect 11576 22330 11582 22332
rect 11638 22330 11662 22332
rect 11718 22330 11742 22332
rect 11798 22330 11822 22332
rect 11878 22330 11884 22332
rect 11638 22278 11640 22330
rect 11820 22278 11822 22330
rect 11576 22276 11582 22278
rect 11638 22276 11662 22278
rect 11718 22276 11742 22278
rect 11798 22276 11822 22278
rect 11878 22276 11884 22278
rect 11576 22267 11884 22276
rect 11992 22234 12020 22646
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 11576 21244 11884 21253
rect 11576 21242 11582 21244
rect 11638 21242 11662 21244
rect 11718 21242 11742 21244
rect 11798 21242 11822 21244
rect 11878 21242 11884 21244
rect 11638 21190 11640 21242
rect 11820 21190 11822 21242
rect 11576 21188 11582 21190
rect 11638 21188 11662 21190
rect 11718 21188 11742 21190
rect 11798 21188 11822 21190
rect 11878 21188 11884 21190
rect 11576 21179 11884 21188
rect 12452 21146 12480 21490
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11992 20602 12020 20878
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11576 20156 11884 20165
rect 11576 20154 11582 20156
rect 11638 20154 11662 20156
rect 11718 20154 11742 20156
rect 11798 20154 11822 20156
rect 11878 20154 11884 20156
rect 11638 20102 11640 20154
rect 11820 20102 11822 20154
rect 11576 20100 11582 20102
rect 11638 20100 11662 20102
rect 11718 20100 11742 20102
rect 11798 20100 11822 20102
rect 11878 20100 11884 20102
rect 11576 20091 11884 20100
rect 11518 19816 11574 19825
rect 11518 19751 11520 19760
rect 11572 19751 11574 19760
rect 11520 19722 11572 19728
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 11256 19306 11376 19334
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 17746 11100 18022
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10692 15438 10744 15444
rect 10874 15464 10930 15473
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10428 13530 10456 13806
rect 10520 13530 10548 14350
rect 10612 14074 10640 14962
rect 10704 14890 10732 15438
rect 10874 15399 10930 15408
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10336 12986 10364 13262
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 12374 9996 12582
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9968 12220 9996 12310
rect 10048 12232 10100 12238
rect 9968 12192 10048 12220
rect 10048 12174 10100 12180
rect 10060 11762 10088 12174
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10152 11558 10180 12106
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 8090 8984 8434
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 9048 6322 9076 8910
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7546 9168 7822
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9232 7410 9260 9590
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9232 7002 9260 7346
rect 9416 7342 9444 10474
rect 9508 10266 9536 10610
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9692 9178 9720 9590
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9600 8838 9628 8910
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9784 8566 9812 11018
rect 10336 10062 10364 11834
rect 10428 11830 10456 13466
rect 10612 12850 10640 13670
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10704 12238 10732 14826
rect 10888 14618 10916 14962
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10980 14482 11008 14758
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10704 11150 10732 12174
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10796 11082 10824 12174
rect 10888 11914 10916 14214
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10980 12238 11008 13466
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10888 11886 11192 11914
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10888 10810 10916 11698
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10520 9722 10548 9998
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10796 9178 10824 9998
rect 10980 9586 11008 11494
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10980 9382 11008 9522
rect 11072 9518 11100 11766
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9784 7546 9812 8502
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9784 7342 9812 7482
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9232 6798 9260 6938
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9232 6458 9260 6734
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9324 6322 9352 7210
rect 9416 6934 9444 7278
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9404 6928 9456 6934
rect 9404 6870 9456 6876
rect 9416 6662 9444 6870
rect 9600 6780 9628 6938
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9680 6792 9732 6798
rect 9600 6752 9680 6780
rect 9680 6734 9732 6740
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9048 5914 9076 6258
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9048 5710 9076 5850
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9324 4690 9352 6258
rect 9784 4690 9812 6870
rect 9876 6730 9904 7890
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10152 7206 10180 7686
rect 10336 7410 10364 7686
rect 10704 7478 10732 8230
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10152 6746 10180 7142
rect 10612 6934 10640 7346
rect 10704 7206 10732 7414
rect 10888 7392 10916 7822
rect 10980 7410 11008 9318
rect 11072 9178 11100 9454
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11072 8634 11100 9114
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11072 7546 11100 8570
rect 11164 7818 11192 11886
rect 11256 9625 11284 19306
rect 11576 19068 11884 19077
rect 11576 19066 11582 19068
rect 11638 19066 11662 19068
rect 11718 19066 11742 19068
rect 11798 19066 11822 19068
rect 11878 19066 11884 19068
rect 11638 19014 11640 19066
rect 11820 19014 11822 19066
rect 11576 19012 11582 19014
rect 11638 19012 11662 19014
rect 11718 19012 11742 19014
rect 11798 19012 11822 19014
rect 11878 19012 11884 19014
rect 11576 19003 11884 19012
rect 11980 18352 12032 18358
rect 11980 18294 12032 18300
rect 11576 17980 11884 17989
rect 11576 17978 11582 17980
rect 11638 17978 11662 17980
rect 11718 17978 11742 17980
rect 11798 17978 11822 17980
rect 11878 17978 11884 17980
rect 11638 17926 11640 17978
rect 11820 17926 11822 17978
rect 11576 17924 11582 17926
rect 11638 17924 11662 17926
rect 11718 17924 11742 17926
rect 11798 17924 11822 17926
rect 11878 17924 11884 17926
rect 11576 17915 11884 17924
rect 11992 17882 12020 18294
rect 12084 18290 12112 19450
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11900 17202 11928 17818
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11900 17082 11928 17138
rect 11900 17054 12020 17082
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11440 16590 11468 16934
rect 11576 16892 11884 16901
rect 11576 16890 11582 16892
rect 11638 16890 11662 16892
rect 11718 16890 11742 16892
rect 11798 16890 11822 16892
rect 11878 16890 11884 16892
rect 11638 16838 11640 16890
rect 11820 16838 11822 16890
rect 11576 16836 11582 16838
rect 11638 16836 11662 16838
rect 11718 16836 11742 16838
rect 11798 16836 11822 16838
rect 11878 16836 11884 16838
rect 11576 16827 11884 16836
rect 11428 16584 11480 16590
rect 11888 16584 11940 16590
rect 11428 16526 11480 16532
rect 11886 16552 11888 16561
rect 11940 16552 11942 16561
rect 11886 16487 11942 16496
rect 11992 16114 12020 17054
rect 12176 16590 12204 17478
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11576 15804 11884 15813
rect 11576 15802 11582 15804
rect 11638 15802 11662 15804
rect 11718 15802 11742 15804
rect 11798 15802 11822 15804
rect 11878 15802 11884 15804
rect 11638 15750 11640 15802
rect 11820 15750 11822 15802
rect 11576 15748 11582 15750
rect 11638 15748 11662 15750
rect 11718 15748 11742 15750
rect 11798 15748 11822 15750
rect 11878 15748 11884 15750
rect 11576 15739 11884 15748
rect 11992 15162 12020 15846
rect 12176 15366 12204 16526
rect 12544 16250 12572 23054
rect 13004 22778 13032 24142
rect 13176 23248 13228 23254
rect 13176 23190 13228 23196
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 12900 21684 12952 21690
rect 12900 21626 12952 21632
rect 12912 21554 12940 21626
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 12716 21480 12768 21486
rect 12768 21428 12848 21434
rect 12716 21422 12848 21428
rect 12728 21406 12848 21422
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12636 20602 12664 20878
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 12820 20466 12848 21406
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 12820 19802 12848 20402
rect 12912 20058 12940 21490
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12820 19786 12940 19802
rect 12820 19780 12952 19786
rect 12820 19774 12900 19780
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12636 16794 12664 18158
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12636 16114 12664 16526
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 14414 11376 14758
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11334 12336 11390 12345
rect 11334 12271 11390 12280
rect 11348 12238 11376 12271
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11348 11558 11376 12174
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11348 11218 11376 11494
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11242 9616 11298 9625
rect 11242 9551 11298 9560
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 10796 7364 10916 7392
rect 10968 7404 11020 7410
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10796 6798 10824 7364
rect 10968 7346 11020 7352
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 10060 6718 10180 6746
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10060 5370 10088 6718
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 6186 10180 6598
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9784 4146 9812 4626
rect 10060 4554 10088 5306
rect 10520 4826 10548 6734
rect 10796 6254 10824 6734
rect 10888 6322 10916 7210
rect 10980 6390 11008 7346
rect 11348 7206 11376 7482
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11256 6798 11284 7142
rect 11440 7002 11468 14962
rect 12176 14958 12204 15302
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 11576 14716 11884 14725
rect 11576 14714 11582 14716
rect 11638 14714 11662 14716
rect 11718 14714 11742 14716
rect 11798 14714 11822 14716
rect 11878 14714 11884 14716
rect 11638 14662 11640 14714
rect 11820 14662 11822 14714
rect 11576 14660 11582 14662
rect 11638 14660 11662 14662
rect 11718 14660 11742 14662
rect 11798 14660 11822 14662
rect 11878 14660 11884 14662
rect 11576 14651 11884 14660
rect 11610 14512 11666 14521
rect 11610 14447 11666 14456
rect 11624 14414 11652 14447
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11532 13802 11560 14010
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11624 13734 11652 14214
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11576 13628 11884 13637
rect 11576 13626 11582 13628
rect 11638 13626 11662 13628
rect 11718 13626 11742 13628
rect 11798 13626 11822 13628
rect 11878 13626 11884 13628
rect 11638 13574 11640 13626
rect 11820 13574 11822 13626
rect 11576 13572 11582 13574
rect 11638 13572 11662 13574
rect 11718 13572 11742 13574
rect 11798 13572 11822 13574
rect 11878 13572 11884 13574
rect 11576 13563 11884 13572
rect 11992 12918 12020 14282
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 13870 12664 14214
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12728 13326 12756 19654
rect 12820 17678 12848 19774
rect 12900 19722 12952 19728
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12820 16590 12848 17614
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12912 17338 12940 17478
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 13004 17202 13032 22714
rect 13188 22098 13216 23190
rect 13280 23186 13308 24754
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13188 21486 13216 22034
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 13280 20466 13308 23122
rect 13372 21894 13400 24686
rect 13556 23730 13584 25230
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13452 23588 13504 23594
rect 13452 23530 13504 23536
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13372 21554 13400 21830
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13280 18358 13308 20402
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 13372 19718 13400 20198
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13268 18352 13320 18358
rect 13188 18312 13268 18340
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13188 16658 13216 18312
rect 13268 18294 13320 18300
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 13188 16182 13216 16594
rect 13280 16590 13308 17614
rect 13372 16697 13400 19654
rect 13358 16688 13414 16697
rect 13358 16623 13414 16632
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13176 16176 13228 16182
rect 13176 16118 13228 16124
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12820 13870 12848 15914
rect 12912 15094 12940 15982
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 13004 15026 13032 15846
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 13188 13462 13216 16118
rect 13280 16114 13308 16526
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13464 15162 13492 23530
rect 13556 23118 13584 23666
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13556 22710 13584 23054
rect 13544 22704 13596 22710
rect 13544 22646 13596 22652
rect 13556 21486 13584 22646
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13556 21146 13584 21422
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13556 19922 13584 19994
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13556 17814 13584 19858
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 13556 16658 13584 17750
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13556 16114 13584 16594
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13452 15156 13504 15162
rect 13372 15116 13452 15144
rect 12808 13456 12860 13462
rect 12808 13398 12860 13404
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11576 12540 11884 12549
rect 11576 12538 11582 12540
rect 11638 12538 11662 12540
rect 11718 12538 11742 12540
rect 11798 12538 11822 12540
rect 11878 12538 11884 12540
rect 11638 12486 11640 12538
rect 11820 12486 11822 12538
rect 11576 12484 11582 12486
rect 11638 12484 11662 12486
rect 11718 12484 11742 12486
rect 11798 12484 11822 12486
rect 11878 12484 11884 12486
rect 11576 12475 11884 12484
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11716 12238 11744 12378
rect 11520 12232 11572 12238
rect 11704 12232 11756 12238
rect 11572 12192 11652 12220
rect 11520 12174 11572 12180
rect 11520 12096 11572 12102
rect 11624 12084 11652 12192
rect 11704 12174 11756 12180
rect 11992 12084 12020 12854
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12084 12442 12112 12786
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12636 12238 12664 13126
rect 12820 12782 12848 13398
rect 13372 13326 13400 15116
rect 13452 15098 13504 15104
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13556 14618 13584 14962
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 11624 12056 12020 12084
rect 11520 12038 11572 12044
rect 11532 11898 11560 12038
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11576 11452 11884 11461
rect 11576 11450 11582 11452
rect 11638 11450 11662 11452
rect 11718 11450 11742 11452
rect 11798 11450 11822 11452
rect 11878 11450 11884 11452
rect 11638 11398 11640 11450
rect 11820 11398 11822 11450
rect 11576 11396 11582 11398
rect 11638 11396 11662 11398
rect 11718 11396 11742 11398
rect 11798 11396 11822 11398
rect 11878 11396 11884 11398
rect 11576 11387 11884 11396
rect 11992 10538 12020 12056
rect 12820 11762 12848 12718
rect 13372 12238 13400 13262
rect 13464 12850 13492 13262
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13004 11762 13032 12174
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11576 10364 11884 10373
rect 11576 10362 11582 10364
rect 11638 10362 11662 10364
rect 11718 10362 11742 10364
rect 11798 10362 11822 10364
rect 11878 10362 11884 10364
rect 11638 10310 11640 10362
rect 11820 10310 11822 10362
rect 11576 10308 11582 10310
rect 11638 10308 11662 10310
rect 11718 10308 11742 10310
rect 11798 10308 11822 10310
rect 11878 10308 11884 10310
rect 11576 10299 11884 10308
rect 12728 10266 12756 10950
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12268 9518 12296 9930
rect 12360 9722 12388 9998
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 11576 9276 11884 9285
rect 11576 9274 11582 9276
rect 11638 9274 11662 9276
rect 11718 9274 11742 9276
rect 11798 9274 11822 9276
rect 11878 9274 11884 9276
rect 11638 9222 11640 9274
rect 11820 9222 11822 9274
rect 11576 9220 11582 9222
rect 11638 9220 11662 9222
rect 11718 9220 11742 9222
rect 11798 9220 11822 9222
rect 11878 9220 11884 9222
rect 11576 9211 11884 9220
rect 12268 8566 12296 9454
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 11576 8188 11884 8197
rect 11576 8186 11582 8188
rect 11638 8186 11662 8188
rect 11718 8186 11742 8188
rect 11798 8186 11822 8188
rect 11878 8186 11884 8188
rect 11638 8134 11640 8186
rect 11820 8134 11822 8186
rect 11576 8132 11582 8134
rect 11638 8132 11662 8134
rect 11718 8132 11742 8134
rect 11798 8132 11822 8134
rect 11878 8132 11884 8134
rect 11576 8123 11884 8132
rect 12452 8090 12480 9998
rect 12820 9586 12848 11494
rect 12898 11248 12954 11257
rect 13188 11234 13216 11698
rect 13188 11206 13400 11234
rect 13556 11218 13584 12582
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 12898 11183 12900 11192
rect 12952 11183 12954 11192
rect 12900 11154 12952 11160
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12912 10674 12940 11018
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12912 10470 12940 10610
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12532 9512 12584 9518
rect 12584 9472 12664 9500
rect 12532 9454 12584 9460
rect 12636 9382 12664 9472
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12544 7546 12572 9318
rect 12912 8838 12940 10406
rect 13004 10062 13032 10950
rect 13188 10266 13216 11086
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 13096 9518 13124 9930
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12636 7274 12664 8774
rect 13096 8430 13124 9454
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 13096 8090 13124 8366
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13004 7478 13032 7686
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 11576 7100 11884 7109
rect 11576 7098 11582 7100
rect 11638 7098 11662 7100
rect 11718 7098 11742 7100
rect 11798 7098 11822 7100
rect 11878 7098 11884 7100
rect 11638 7046 11640 7098
rect 11820 7046 11822 7098
rect 11576 7044 11582 7046
rect 11638 7044 11662 7046
rect 11718 7044 11742 7046
rect 11798 7044 11822 7046
rect 11878 7044 11884 7046
rect 11576 7035 11884 7044
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11348 6458 11376 6734
rect 12360 6662 12388 7142
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6458 12388 6598
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 12452 6322 12480 6734
rect 12728 6458 12756 7346
rect 12912 7002 12940 7346
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10612 5914 10640 6190
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10520 4622 10548 4762
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10612 4554 10640 5850
rect 10888 5370 10916 6258
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 10060 4010 10088 4490
rect 10612 4282 10640 4490
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10060 3194 10088 3946
rect 10612 3466 10640 4218
rect 10980 4146 11008 6190
rect 12728 6186 12756 6394
rect 13188 6322 13216 7278
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13280 6458 13308 6734
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10980 4026 11008 4082
rect 10888 3998 11008 4026
rect 11440 4010 11468 6054
rect 11576 6012 11884 6021
rect 11576 6010 11582 6012
rect 11638 6010 11662 6012
rect 11718 6010 11742 6012
rect 11798 6010 11822 6012
rect 11878 6010 11884 6012
rect 11638 5958 11640 6010
rect 11820 5958 11822 6010
rect 11576 5956 11582 5958
rect 11638 5956 11662 5958
rect 11718 5956 11742 5958
rect 11798 5956 11822 5958
rect 11878 5956 11884 5958
rect 11576 5947 11884 5956
rect 13188 5642 13216 6258
rect 13280 5710 13308 6258
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 11576 4924 11884 4933
rect 11576 4922 11582 4924
rect 11638 4922 11662 4924
rect 11718 4922 11742 4924
rect 11798 4922 11822 4924
rect 11878 4922 11884 4924
rect 11638 4870 11640 4922
rect 11820 4870 11822 4922
rect 11576 4868 11582 4870
rect 11638 4868 11662 4870
rect 11718 4868 11742 4870
rect 11798 4868 11822 4870
rect 11878 4868 11884 4870
rect 11576 4859 11884 4868
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11428 4004 11480 4010
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10612 3194 10640 3402
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10888 3058 10916 3998
rect 11428 3946 11480 3952
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10980 3602 11008 3878
rect 11440 3602 11468 3946
rect 11576 3836 11884 3845
rect 11576 3834 11582 3836
rect 11638 3834 11662 3836
rect 11718 3834 11742 3836
rect 11798 3834 11822 3836
rect 11878 3834 11884 3836
rect 11638 3782 11640 3834
rect 11820 3782 11822 3834
rect 11576 3780 11582 3782
rect 11638 3780 11662 3782
rect 11718 3780 11742 3782
rect 11798 3780 11822 3782
rect 11878 3780 11884 3782
rect 11576 3771 11884 3780
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11992 3534 12020 4082
rect 12636 3534 12664 4626
rect 13372 3618 13400 11206
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13648 10674 13676 12038
rect 13740 11762 13768 27474
rect 13832 27470 13860 27814
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 13924 26246 13952 30126
rect 17960 30116 18012 30122
rect 17960 30058 18012 30064
rect 16028 30048 16080 30054
rect 16028 29990 16080 29996
rect 15660 29776 15712 29782
rect 15660 29718 15712 29724
rect 15118 29404 15426 29413
rect 15118 29402 15124 29404
rect 15180 29402 15204 29404
rect 15260 29402 15284 29404
rect 15340 29402 15364 29404
rect 15420 29402 15426 29404
rect 15180 29350 15182 29402
rect 15362 29350 15364 29402
rect 15118 29348 15124 29350
rect 15180 29348 15204 29350
rect 15260 29348 15284 29350
rect 15340 29348 15364 29350
rect 15420 29348 15426 29350
rect 15118 29339 15426 29348
rect 15672 29102 15700 29718
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 15476 28960 15528 28966
rect 15476 28902 15528 28908
rect 14830 28656 14886 28665
rect 14830 28591 14832 28600
rect 14884 28591 14886 28600
rect 14832 28562 14884 28568
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 14568 27674 14596 28494
rect 15118 28316 15426 28325
rect 15118 28314 15124 28316
rect 15180 28314 15204 28316
rect 15260 28314 15284 28316
rect 15340 28314 15364 28316
rect 15420 28314 15426 28316
rect 15180 28262 15182 28314
rect 15362 28262 15364 28314
rect 15118 28260 15124 28262
rect 15180 28260 15204 28262
rect 15260 28260 15284 28262
rect 15340 28260 15364 28262
rect 15420 28260 15426 28262
rect 15118 28251 15426 28260
rect 15488 28218 15516 28902
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 15856 28218 15884 28494
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 15844 28212 15896 28218
rect 15844 28154 15896 28160
rect 14832 28144 14884 28150
rect 14832 28086 14884 28092
rect 14556 27668 14608 27674
rect 14556 27610 14608 27616
rect 14648 27668 14700 27674
rect 14648 27610 14700 27616
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14096 26784 14148 26790
rect 14096 26726 14148 26732
rect 14108 26314 14136 26726
rect 14384 26586 14412 26998
rect 14372 26580 14424 26586
rect 14372 26522 14424 26528
rect 14096 26308 14148 26314
rect 14096 26250 14148 26256
rect 14280 26308 14332 26314
rect 14280 26250 14332 26256
rect 13912 26240 13964 26246
rect 13912 26182 13964 26188
rect 13924 26042 13952 26182
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13924 25158 13952 25978
rect 14004 25968 14056 25974
rect 14004 25910 14056 25916
rect 13912 25152 13964 25158
rect 13912 25094 13964 25100
rect 13924 24818 13952 25094
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 14016 24750 14044 25910
rect 14108 25906 14136 26250
rect 14292 26042 14320 26250
rect 14280 26036 14332 26042
rect 14280 25978 14332 25984
rect 14384 25906 14412 26522
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 14372 25900 14424 25906
rect 14372 25842 14424 25848
rect 14464 25900 14516 25906
rect 14464 25842 14516 25848
rect 14108 25498 14136 25842
rect 14096 25492 14148 25498
rect 14096 25434 14148 25440
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 14016 24206 14044 24686
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 13912 24132 13964 24138
rect 13912 24074 13964 24080
rect 13924 21690 13952 24074
rect 14476 23866 14504 25842
rect 14660 23866 14688 27610
rect 14844 26858 14872 28086
rect 14924 28076 14976 28082
rect 14924 28018 14976 28024
rect 14832 26852 14884 26858
rect 14832 26794 14884 26800
rect 14832 25832 14884 25838
rect 14832 25774 14884 25780
rect 14844 24954 14872 25774
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14740 24676 14792 24682
rect 14740 24618 14792 24624
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14648 23860 14700 23866
rect 14648 23802 14700 23808
rect 14372 23724 14424 23730
rect 14372 23666 14424 23672
rect 14188 23588 14240 23594
rect 14188 23530 14240 23536
rect 14200 23322 14228 23530
rect 14384 23322 14412 23666
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14096 23044 14148 23050
rect 14096 22986 14148 22992
rect 14108 21690 14136 22986
rect 14200 22030 14228 23258
rect 14384 23118 14412 23258
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14752 22094 14780 24618
rect 14832 23520 14884 23526
rect 14832 23462 14884 23468
rect 14844 22778 14872 23462
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14936 22098 14964 28018
rect 15660 27600 15712 27606
rect 15660 27542 15712 27548
rect 15118 27228 15426 27237
rect 15118 27226 15124 27228
rect 15180 27226 15204 27228
rect 15260 27226 15284 27228
rect 15340 27226 15364 27228
rect 15420 27226 15426 27228
rect 15180 27174 15182 27226
rect 15362 27174 15364 27226
rect 15118 27172 15124 27174
rect 15180 27172 15204 27174
rect 15260 27172 15284 27174
rect 15340 27172 15364 27174
rect 15420 27172 15426 27174
rect 15118 27163 15426 27172
rect 15672 27130 15700 27542
rect 15844 27328 15896 27334
rect 15844 27270 15896 27276
rect 15856 27130 15884 27270
rect 15660 27124 15712 27130
rect 15660 27066 15712 27072
rect 15844 27124 15896 27130
rect 15844 27066 15896 27072
rect 15200 26988 15252 26994
rect 15200 26930 15252 26936
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 15568 26988 15620 26994
rect 15568 26930 15620 26936
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 15028 26042 15056 26862
rect 15212 26586 15240 26930
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15200 26580 15252 26586
rect 15200 26522 15252 26528
rect 15304 26382 15332 26726
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15396 26228 15424 26930
rect 15580 26450 15608 26930
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 15396 26200 15516 26228
rect 15118 26140 15426 26149
rect 15118 26138 15124 26140
rect 15180 26138 15204 26140
rect 15260 26138 15284 26140
rect 15340 26138 15364 26140
rect 15420 26138 15426 26140
rect 15180 26086 15182 26138
rect 15362 26086 15364 26138
rect 15118 26084 15124 26086
rect 15180 26084 15204 26086
rect 15260 26084 15284 26086
rect 15340 26084 15364 26086
rect 15420 26084 15426 26086
rect 15118 26075 15426 26084
rect 15016 26036 15068 26042
rect 15016 25978 15068 25984
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15304 25140 15332 25842
rect 15384 25764 15436 25770
rect 15488 25752 15516 26200
rect 15580 25906 15608 26386
rect 15672 26382 15700 27066
rect 15856 26382 15884 27066
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15844 26376 15896 26382
rect 15844 26318 15896 26324
rect 15660 26240 15712 26246
rect 15660 26182 15712 26188
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15436 25724 15516 25752
rect 15384 25706 15436 25712
rect 15580 25498 15608 25842
rect 15568 25492 15620 25498
rect 15568 25434 15620 25440
rect 15672 25294 15700 26182
rect 15856 25945 15884 26318
rect 15842 25936 15898 25945
rect 15842 25871 15898 25880
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15304 25112 15516 25140
rect 15118 25052 15426 25061
rect 15118 25050 15124 25052
rect 15180 25050 15204 25052
rect 15260 25050 15284 25052
rect 15340 25050 15364 25052
rect 15420 25050 15426 25052
rect 15180 24998 15182 25050
rect 15362 24998 15364 25050
rect 15118 24996 15124 24998
rect 15180 24996 15204 24998
rect 15260 24996 15284 24998
rect 15340 24996 15364 24998
rect 15420 24996 15426 24998
rect 15118 24987 15426 24996
rect 15488 24886 15516 25112
rect 15476 24880 15528 24886
rect 15476 24822 15528 24828
rect 15016 24064 15068 24070
rect 15016 24006 15068 24012
rect 15028 23202 15056 24006
rect 15118 23964 15426 23973
rect 15118 23962 15124 23964
rect 15180 23962 15204 23964
rect 15260 23962 15284 23964
rect 15340 23962 15364 23964
rect 15420 23962 15426 23964
rect 15180 23910 15182 23962
rect 15362 23910 15364 23962
rect 15118 23908 15124 23910
rect 15180 23908 15204 23910
rect 15260 23908 15284 23910
rect 15340 23908 15364 23910
rect 15420 23908 15426 23910
rect 15118 23899 15426 23908
rect 15488 23202 15516 24822
rect 15844 23792 15896 23798
rect 15844 23734 15896 23740
rect 15752 23588 15804 23594
rect 15752 23530 15804 23536
rect 15028 23186 15148 23202
rect 15028 23180 15160 23186
rect 15028 23174 15108 23180
rect 15108 23122 15160 23128
rect 15396 23174 15516 23202
rect 15396 23118 15424 23174
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15028 22642 15056 23054
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15118 22876 15426 22885
rect 15118 22874 15124 22876
rect 15180 22874 15204 22876
rect 15260 22874 15284 22876
rect 15340 22874 15364 22876
rect 15420 22874 15426 22876
rect 15180 22822 15182 22874
rect 15362 22822 15364 22874
rect 15118 22820 15124 22822
rect 15180 22820 15204 22822
rect 15260 22820 15284 22822
rect 15340 22820 15364 22822
rect 15420 22820 15426 22822
rect 15118 22811 15426 22820
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 14752 22066 14872 22094
rect 14188 22024 14240 22030
rect 14188 21966 14240 21972
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14476 21706 14504 21966
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14384 21690 14504 21706
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 14372 21684 14504 21690
rect 14424 21678 14504 21684
rect 14372 21626 14424 21632
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13832 19378 13860 19654
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13924 19258 13952 19858
rect 14016 19417 14044 21490
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14108 20534 14136 20878
rect 14188 20868 14240 20874
rect 14188 20810 14240 20816
rect 14096 20528 14148 20534
rect 14096 20470 14148 20476
rect 14200 20466 14228 20810
rect 14292 20806 14320 21626
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14384 21350 14412 21490
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14384 20874 14412 21286
rect 14568 20874 14596 21898
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14372 20868 14424 20874
rect 14556 20868 14608 20874
rect 14372 20810 14424 20816
rect 14476 20828 14556 20856
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14292 20602 14320 20742
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14002 19408 14058 19417
rect 14002 19343 14058 19352
rect 13832 19230 13952 19258
rect 13832 17882 13860 19230
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13832 17066 13860 17818
rect 13924 17354 13952 19110
rect 14016 18086 14044 19343
rect 14200 18698 14228 20402
rect 14476 19922 14504 20828
rect 14556 20810 14608 20816
rect 14556 20256 14608 20262
rect 14556 20198 14608 20204
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14568 19854 14596 20198
rect 14660 19990 14688 20878
rect 14648 19984 14700 19990
rect 14648 19926 14700 19932
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14660 19378 14688 19926
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 14108 17678 14136 18566
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14292 17678 14320 18022
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 13924 17326 14044 17354
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13924 16794 13952 17138
rect 14016 16810 14044 17326
rect 14108 16998 14136 17478
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 13912 16788 13964 16794
rect 14016 16782 14136 16810
rect 13912 16730 13964 16736
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 12238 13860 16390
rect 13924 16114 13952 16730
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13740 11558 13768 11698
rect 13924 11626 13952 15302
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14016 14006 14044 14962
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 14108 12434 14136 16782
rect 14292 14414 14320 16934
rect 14384 14498 14412 18158
rect 14464 17604 14516 17610
rect 14464 17546 14516 17552
rect 14476 15910 14504 17546
rect 14660 17338 14688 18226
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14556 16448 14608 16454
rect 14752 16436 14780 21966
rect 14608 16408 14780 16436
rect 14556 16390 14608 16396
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14660 15570 14688 15846
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14660 15026 14688 15506
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14384 14470 14596 14498
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14292 13938 14320 14350
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14384 12986 14412 13466
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14476 12442 14504 12922
rect 14016 12406 14136 12434
rect 14464 12436 14516 12442
rect 13912 11620 13964 11626
rect 13912 11562 13964 11568
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13464 9042 13492 10610
rect 13740 10554 13768 11494
rect 13648 10526 13768 10554
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 9994 13584 10406
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13648 8906 13676 10526
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10198 13768 10406
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13740 8906 13768 9590
rect 13832 9042 13860 10066
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13924 9518 13952 9862
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13648 8430 13676 8842
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13832 6730 13860 8978
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13924 7818 13952 8434
rect 13912 7812 13964 7818
rect 13912 7754 13964 7760
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13832 5846 13860 6666
rect 13924 6118 13952 6938
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13832 5370 13860 5646
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13556 3738 13584 4014
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13648 3618 13676 3674
rect 13372 3590 13676 3618
rect 13372 3534 13400 3590
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11532 3194 11560 3402
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 12544 3058 12572 3334
rect 12636 3194 12664 3470
rect 13924 3194 13952 3470
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 11576 2748 11884 2757
rect 11576 2746 11582 2748
rect 11638 2746 11662 2748
rect 11718 2746 11742 2748
rect 11798 2746 11822 2748
rect 11878 2746 11884 2748
rect 11638 2694 11640 2746
rect 11820 2694 11822 2746
rect 11576 2692 11582 2694
rect 11638 2692 11662 2694
rect 11718 2692 11742 2694
rect 11798 2692 11822 2694
rect 11878 2692 11884 2694
rect 11576 2683 11884 2692
rect 14016 2650 14044 12406
rect 14464 12378 14516 12384
rect 14568 12170 14596 14470
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14660 12986 14688 14282
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14752 12986 14780 13670
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14752 12850 14780 12922
rect 14740 12844 14792 12850
rect 14660 12804 14740 12832
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14568 11898 14596 12106
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14660 11150 14688 12804
rect 14740 12786 14792 12792
rect 14844 12434 14872 22066
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 15118 21788 15426 21797
rect 15118 21786 15124 21788
rect 15180 21786 15204 21788
rect 15260 21786 15284 21788
rect 15340 21786 15364 21788
rect 15420 21786 15426 21788
rect 15180 21734 15182 21786
rect 15362 21734 15364 21786
rect 15118 21732 15124 21734
rect 15180 21732 15204 21734
rect 15260 21732 15284 21734
rect 15340 21732 15364 21734
rect 15420 21732 15426 21734
rect 15118 21723 15426 21732
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 14936 16250 14964 21490
rect 15396 20856 15424 21558
rect 15396 20828 15516 20856
rect 15118 20700 15426 20709
rect 15118 20698 15124 20700
rect 15180 20698 15204 20700
rect 15260 20698 15284 20700
rect 15340 20698 15364 20700
rect 15420 20698 15426 20700
rect 15180 20646 15182 20698
rect 15362 20646 15364 20698
rect 15118 20644 15124 20646
rect 15180 20644 15204 20646
rect 15260 20644 15284 20646
rect 15340 20644 15364 20646
rect 15420 20644 15426 20646
rect 15118 20635 15426 20644
rect 15118 19612 15426 19621
rect 15118 19610 15124 19612
rect 15180 19610 15204 19612
rect 15260 19610 15284 19612
rect 15340 19610 15364 19612
rect 15420 19610 15426 19612
rect 15180 19558 15182 19610
rect 15362 19558 15364 19610
rect 15118 19556 15124 19558
rect 15180 19556 15204 19558
rect 15260 19556 15284 19558
rect 15340 19556 15364 19558
rect 15420 19556 15426 19558
rect 15118 19547 15426 19556
rect 15488 18970 15516 20828
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 15028 18290 15056 18634
rect 15118 18524 15426 18533
rect 15118 18522 15124 18524
rect 15180 18522 15204 18524
rect 15260 18522 15284 18524
rect 15340 18522 15364 18524
rect 15420 18522 15426 18524
rect 15180 18470 15182 18522
rect 15362 18470 15364 18522
rect 15118 18468 15124 18470
rect 15180 18468 15204 18470
rect 15260 18468 15284 18470
rect 15340 18468 15364 18470
rect 15420 18468 15426 18470
rect 15118 18459 15426 18468
rect 15488 18358 15516 18906
rect 15580 18834 15608 19654
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15672 18714 15700 22918
rect 15764 22710 15792 23530
rect 15856 23322 15884 23734
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15752 22704 15804 22710
rect 15752 22646 15804 22652
rect 16040 19174 16068 29990
rect 17972 29646 18000 30058
rect 18660 29948 18968 29957
rect 18660 29946 18666 29948
rect 18722 29946 18746 29948
rect 18802 29946 18826 29948
rect 18882 29946 18906 29948
rect 18962 29946 18968 29948
rect 18722 29894 18724 29946
rect 18904 29894 18906 29946
rect 18660 29892 18666 29894
rect 18722 29892 18746 29894
rect 18802 29892 18826 29894
rect 18882 29892 18906 29894
rect 18962 29892 18968 29894
rect 18660 29883 18968 29892
rect 19996 29850 20024 30194
rect 22652 30116 22704 30122
rect 22652 30058 22704 30064
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 22008 30048 22060 30054
rect 22008 29990 22060 29996
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 18236 29708 18288 29714
rect 18236 29650 18288 29656
rect 16856 29640 16908 29646
rect 16856 29582 16908 29588
rect 17868 29640 17920 29646
rect 17868 29582 17920 29588
rect 17960 29640 18012 29646
rect 17960 29582 18012 29588
rect 16868 29306 16896 29582
rect 17224 29504 17276 29510
rect 17224 29446 17276 29452
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 16580 29232 16632 29238
rect 16580 29174 16632 29180
rect 16212 28688 16264 28694
rect 16212 28630 16264 28636
rect 16224 28529 16252 28630
rect 16304 28552 16356 28558
rect 16210 28520 16266 28529
rect 16304 28494 16356 28500
rect 16210 28455 16212 28464
rect 16264 28455 16266 28464
rect 16212 28426 16264 28432
rect 16224 28395 16252 28426
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 16132 25498 16160 27406
rect 16212 27328 16264 27334
rect 16212 27270 16264 27276
rect 16224 26246 16252 27270
rect 16316 26586 16344 28494
rect 16592 27062 16620 29174
rect 16868 29170 16896 29242
rect 17236 29170 17264 29446
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16948 29164 17000 29170
rect 16948 29106 17000 29112
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 16960 28490 16988 29106
rect 17880 29102 17908 29582
rect 17972 29170 18000 29582
rect 17960 29164 18012 29170
rect 17960 29106 18012 29112
rect 17868 29096 17920 29102
rect 17868 29038 17920 29044
rect 18248 28626 18276 29650
rect 19156 29232 19208 29238
rect 19156 29174 19208 29180
rect 18660 28860 18968 28869
rect 18660 28858 18666 28860
rect 18722 28858 18746 28860
rect 18802 28858 18826 28860
rect 18882 28858 18906 28860
rect 18962 28858 18968 28860
rect 18722 28806 18724 28858
rect 18904 28806 18906 28858
rect 18660 28804 18666 28806
rect 18722 28804 18746 28806
rect 18802 28804 18826 28806
rect 18882 28804 18906 28806
rect 18962 28804 18968 28806
rect 18660 28795 18968 28804
rect 19168 28626 19196 29174
rect 19616 29164 19668 29170
rect 19616 29106 19668 29112
rect 19248 29028 19300 29034
rect 19248 28970 19300 28976
rect 19260 28694 19288 28970
rect 19628 28762 19656 29106
rect 19984 29028 20036 29034
rect 19984 28970 20036 28976
rect 19800 28960 19852 28966
rect 19800 28902 19852 28908
rect 19616 28756 19668 28762
rect 19616 28698 19668 28704
rect 19248 28688 19300 28694
rect 19248 28630 19300 28636
rect 18236 28620 18288 28626
rect 18236 28562 18288 28568
rect 19156 28620 19208 28626
rect 19156 28562 19208 28568
rect 16948 28484 17000 28490
rect 16948 28426 17000 28432
rect 16672 28008 16724 28014
rect 16670 27976 16672 27985
rect 16724 27976 16726 27985
rect 16670 27911 16726 27920
rect 16580 27056 16632 27062
rect 16580 26998 16632 27004
rect 16672 27056 16724 27062
rect 16672 26998 16724 27004
rect 16304 26580 16356 26586
rect 16304 26522 16356 26528
rect 16592 26314 16620 26998
rect 16684 26382 16712 26998
rect 17132 26784 17184 26790
rect 17132 26726 17184 26732
rect 18144 26784 18196 26790
rect 18144 26726 18196 26732
rect 17144 26382 17172 26726
rect 17408 26512 17460 26518
rect 17408 26454 17460 26460
rect 16672 26376 16724 26382
rect 16948 26376 17000 26382
rect 16672 26318 16724 26324
rect 16946 26344 16948 26353
rect 17132 26376 17184 26382
rect 17000 26344 17002 26353
rect 16580 26308 16632 26314
rect 16580 26250 16632 26256
rect 16212 26240 16264 26246
rect 16212 26182 16264 26188
rect 16120 25492 16172 25498
rect 16120 25434 16172 25440
rect 16684 25362 16712 26318
rect 17132 26318 17184 26324
rect 16946 26279 17002 26288
rect 16764 25968 16816 25974
rect 16764 25910 16816 25916
rect 16776 25770 16804 25910
rect 17224 25832 17276 25838
rect 17224 25774 17276 25780
rect 16764 25764 16816 25770
rect 16764 25706 16816 25712
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16396 25152 16448 25158
rect 16396 25094 16448 25100
rect 16302 23216 16358 23225
rect 16302 23151 16358 23160
rect 16316 23118 16344 23151
rect 16304 23112 16356 23118
rect 16304 23054 16356 23060
rect 16408 22574 16436 25094
rect 17236 24614 17264 25774
rect 17420 25498 17448 26454
rect 18050 26344 18106 26353
rect 18156 26314 18184 26726
rect 18050 26279 18106 26288
rect 18144 26308 18196 26314
rect 18064 25838 18092 26279
rect 18144 26250 18196 26256
rect 18052 25832 18104 25838
rect 18248 25786 18276 28562
rect 19156 28416 19208 28422
rect 19156 28358 19208 28364
rect 19168 28082 19196 28358
rect 19812 28218 19840 28902
rect 19996 28422 20024 28970
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19800 28212 19852 28218
rect 19800 28154 19852 28160
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 19616 28008 19668 28014
rect 19616 27950 19668 27956
rect 18512 27872 18564 27878
rect 18512 27814 18564 27820
rect 18420 26784 18472 26790
rect 18420 26726 18472 26732
rect 18328 26512 18380 26518
rect 18328 26454 18380 26460
rect 18340 26382 18368 26454
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18328 25968 18380 25974
rect 18328 25910 18380 25916
rect 18052 25774 18104 25780
rect 18156 25758 18276 25786
rect 17408 25492 17460 25498
rect 17408 25434 17460 25440
rect 17684 25220 17736 25226
rect 17684 25162 17736 25168
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17236 23730 17264 24006
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 17040 23588 17092 23594
rect 17040 23530 17092 23536
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16488 23112 16540 23118
rect 16488 23054 16540 23060
rect 16396 22568 16448 22574
rect 16396 22510 16448 22516
rect 16500 21418 16528 23054
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 16684 22778 16712 22986
rect 16672 22772 16724 22778
rect 16672 22714 16724 22720
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16488 21412 16540 21418
rect 16488 21354 16540 21360
rect 16592 21146 16620 21422
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16408 20602 16436 20878
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16132 19514 16160 19790
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 16592 19174 16620 20538
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16684 19378 16712 19654
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16776 19258 16804 23462
rect 17052 23322 17080 23530
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17040 23316 17092 23322
rect 17040 23258 17092 23264
rect 16948 23180 17000 23186
rect 16948 23122 17000 23128
rect 16960 22642 16988 23122
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16948 22636 17000 22642
rect 16948 22578 17000 22584
rect 16868 21962 16896 22578
rect 16856 21956 16908 21962
rect 16856 21898 16908 21904
rect 16868 20942 16896 21898
rect 17512 21894 17540 23462
rect 17500 21888 17552 21894
rect 17498 21856 17500 21865
rect 17552 21856 17554 21865
rect 17498 21791 17554 21800
rect 16948 21684 17000 21690
rect 16948 21626 17000 21632
rect 16960 21078 16988 21626
rect 17040 21548 17092 21554
rect 17040 21490 17092 21496
rect 16948 21072 17000 21078
rect 16948 21014 17000 21020
rect 16856 20936 16908 20942
rect 16856 20878 16908 20884
rect 16868 19378 16896 20878
rect 17052 19514 17080 21490
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17144 21146 17172 21422
rect 17328 21146 17356 21422
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 17328 20602 17356 21082
rect 17420 20942 17448 21286
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17696 20602 17724 25162
rect 18156 22778 18184 25758
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18248 25498 18276 25638
rect 18236 25492 18288 25498
rect 18236 25434 18288 25440
rect 18248 25158 18276 25434
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 18144 22772 18196 22778
rect 18144 22714 18196 22720
rect 17868 22500 17920 22506
rect 17868 22442 17920 22448
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17316 20596 17368 20602
rect 17316 20538 17368 20544
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17696 19990 17724 20538
rect 17788 20262 17816 21422
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17684 19984 17736 19990
rect 17684 19926 17736 19932
rect 17316 19780 17368 19786
rect 17316 19722 17368 19728
rect 17328 19514 17356 19722
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16684 19230 16804 19258
rect 16868 19258 16896 19314
rect 16868 19230 16988 19258
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16316 18902 16344 19110
rect 16304 18896 16356 18902
rect 16304 18838 16356 18844
rect 15580 18686 15700 18714
rect 15580 18630 15608 18686
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15580 18426 15608 18566
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15476 18352 15528 18358
rect 15476 18294 15528 18300
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 15856 17542 15884 18566
rect 16316 17610 16344 18838
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16592 17746 16620 18158
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15118 17436 15426 17445
rect 15118 17434 15124 17436
rect 15180 17434 15204 17436
rect 15260 17434 15284 17436
rect 15340 17434 15364 17436
rect 15420 17434 15426 17436
rect 15180 17382 15182 17434
rect 15362 17382 15364 17434
rect 15118 17380 15124 17382
rect 15180 17380 15204 17382
rect 15260 17380 15284 17382
rect 15340 17380 15364 17382
rect 15420 17380 15426 17382
rect 15118 17371 15426 17380
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15212 16454 15240 17274
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15118 16348 15426 16357
rect 15118 16346 15124 16348
rect 15180 16346 15204 16348
rect 15260 16346 15284 16348
rect 15340 16346 15364 16348
rect 15420 16346 15426 16348
rect 15180 16294 15182 16346
rect 15362 16294 15364 16346
rect 15118 16292 15124 16294
rect 15180 16292 15204 16294
rect 15260 16292 15284 16294
rect 15340 16292 15364 16294
rect 15420 16292 15426 16294
rect 15118 16283 15426 16292
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 15028 15366 15056 16118
rect 15488 15502 15516 17070
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15580 15638 15608 17002
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16224 15978 16252 16186
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 15118 15260 15426 15269
rect 15118 15258 15124 15260
rect 15180 15258 15204 15260
rect 15260 15258 15284 15260
rect 15340 15258 15364 15260
rect 15420 15258 15426 15260
rect 15180 15206 15182 15258
rect 15362 15206 15364 15258
rect 15118 15204 15124 15206
rect 15180 15204 15204 15206
rect 15260 15204 15284 15206
rect 15340 15204 15364 15206
rect 15420 15204 15426 15206
rect 15118 15195 15426 15204
rect 15488 14346 15516 15438
rect 16316 14822 16344 17546
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16408 15706 16436 16390
rect 16500 15706 16528 16458
rect 16592 16250 16620 17478
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16394 15464 16450 15473
rect 16394 15399 16450 15408
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15118 14172 15426 14181
rect 15118 14170 15124 14172
rect 15180 14170 15204 14172
rect 15260 14170 15284 14172
rect 15340 14170 15364 14172
rect 15420 14170 15426 14172
rect 15180 14118 15182 14170
rect 15362 14118 15364 14170
rect 15118 14116 15124 14118
rect 15180 14116 15204 14118
rect 15260 14116 15284 14118
rect 15340 14116 15364 14118
rect 15420 14116 15426 14118
rect 15118 14107 15426 14116
rect 15580 14074 15608 14350
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15396 13954 15424 14010
rect 15672 13954 15700 14758
rect 15396 13926 15700 13954
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15856 13190 15884 13874
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15118 13084 15426 13093
rect 15118 13082 15124 13084
rect 15180 13082 15204 13084
rect 15260 13082 15284 13084
rect 15340 13082 15364 13084
rect 15420 13082 15426 13084
rect 15180 13030 15182 13082
rect 15362 13030 15364 13082
rect 15118 13028 15124 13030
rect 15180 13028 15204 13030
rect 15260 13028 15284 13030
rect 15340 13028 15364 13030
rect 15420 13028 15426 13030
rect 15118 13019 15426 13028
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 14844 12406 14964 12434
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14200 10810 14228 11086
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14384 10577 14412 11086
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14554 10704 14610 10713
rect 14554 10639 14556 10648
rect 14608 10639 14610 10648
rect 14556 10610 14608 10616
rect 14370 10568 14426 10577
rect 14370 10503 14426 10512
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14108 9110 14136 9522
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14108 8498 14136 9046
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14108 8022 14136 8434
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14200 7478 14228 9318
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14476 8974 14504 9046
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14108 6458 14136 7142
rect 14292 6866 14320 7686
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 14384 7002 14412 7414
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14200 6322 14228 6734
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14200 5914 14228 6258
rect 14292 6254 14320 6802
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14292 4622 14320 6190
rect 14476 5914 14504 7958
rect 14568 6458 14596 9454
rect 14660 9450 14688 10950
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14752 8498 14780 12038
rect 14936 9586 14964 12406
rect 15028 11218 15056 12650
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15120 12374 15148 12582
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15396 12306 15424 12718
rect 15856 12442 15884 13126
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 16040 12238 16068 12582
rect 16408 12374 16436 15399
rect 16500 12850 16528 15642
rect 16684 15502 16712 19230
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16776 18834 16804 19110
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16776 18086 16804 18770
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 16868 18290 16896 18566
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16960 18222 16988 19230
rect 17052 18766 17080 19450
rect 17696 19334 17724 19926
rect 17788 19922 17816 20198
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17604 19306 17724 19334
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17130 17776 17186 17785
rect 17130 17711 17132 17720
rect 17184 17711 17186 17720
rect 17132 17682 17184 17688
rect 17144 17338 17172 17682
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 17224 17060 17276 17066
rect 17224 17002 17276 17008
rect 17236 16726 17264 17002
rect 17224 16720 17276 16726
rect 17224 16662 17276 16668
rect 17328 16454 17356 18022
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 17236 15366 17264 16118
rect 17328 16046 17356 16390
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 16776 15162 16804 15302
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17052 12986 17080 14350
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16500 12238 16528 12378
rect 15568 12232 15620 12238
rect 15382 12200 15438 12209
rect 15568 12174 15620 12180
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 15382 12135 15384 12144
rect 15436 12135 15438 12144
rect 15384 12106 15436 12112
rect 15118 11996 15426 12005
rect 15118 11994 15124 11996
rect 15180 11994 15204 11996
rect 15260 11994 15284 11996
rect 15340 11994 15364 11996
rect 15420 11994 15426 11996
rect 15180 11942 15182 11994
rect 15362 11942 15364 11994
rect 15118 11940 15124 11942
rect 15180 11940 15204 11942
rect 15260 11940 15284 11942
rect 15340 11940 15364 11942
rect 15420 11940 15426 11942
rect 15118 11931 15426 11940
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15118 10908 15426 10917
rect 15118 10906 15124 10908
rect 15180 10906 15204 10908
rect 15260 10906 15284 10908
rect 15340 10906 15364 10908
rect 15420 10906 15426 10908
rect 15180 10854 15182 10906
rect 15362 10854 15364 10906
rect 15118 10852 15124 10854
rect 15180 10852 15204 10854
rect 15260 10852 15284 10854
rect 15340 10852 15364 10854
rect 15420 10852 15426 10854
rect 15118 10843 15426 10852
rect 15118 9820 15426 9829
rect 15118 9818 15124 9820
rect 15180 9818 15204 9820
rect 15260 9818 15284 9820
rect 15340 9818 15364 9820
rect 15420 9818 15426 9820
rect 15180 9766 15182 9818
rect 15362 9766 15364 9818
rect 15118 9764 15124 9766
rect 15180 9764 15204 9766
rect 15260 9764 15284 9766
rect 15340 9764 15364 9766
rect 15420 9764 15426 9766
rect 15118 9755 15426 9764
rect 15290 9616 15346 9625
rect 14924 9580 14976 9586
rect 15290 9551 15292 9560
rect 14924 9522 14976 9528
rect 15344 9551 15346 9560
rect 15292 9522 15344 9528
rect 14936 9466 14964 9522
rect 14936 9438 15148 9466
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14844 8634 14872 8978
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14660 7546 14688 8434
rect 14844 8022 14872 8570
rect 14936 8566 14964 9318
rect 15120 9042 15148 9438
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15118 8732 15426 8741
rect 15118 8730 15124 8732
rect 15180 8730 15204 8732
rect 15260 8730 15284 8732
rect 15340 8730 15364 8732
rect 15420 8730 15426 8732
rect 15180 8678 15182 8730
rect 15362 8678 15364 8730
rect 15118 8676 15124 8678
rect 15180 8676 15204 8678
rect 15260 8676 15284 8678
rect 15340 8676 15364 8678
rect 15420 8676 15426 8678
rect 15118 8667 15426 8676
rect 15488 8634 15516 8774
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 14832 8016 14884 8022
rect 14832 7958 14884 7964
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14752 6662 14780 7414
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14384 4826 14412 5306
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14292 4146 14320 4558
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14108 3126 14136 3878
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14108 2854 14136 3062
rect 14384 3058 14412 4422
rect 14476 4078 14504 4694
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14568 4146 14596 4558
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14476 3194 14504 3470
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14936 3058 14964 4150
rect 15028 4010 15056 8230
rect 15488 7886 15516 8434
rect 15580 8362 15608 12174
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15672 8090 15700 8434
rect 15764 8090 15792 9998
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15660 7880 15712 7886
rect 15764 7868 15792 8026
rect 15712 7840 15792 7868
rect 15936 7880 15988 7886
rect 15660 7822 15712 7828
rect 15936 7822 15988 7828
rect 15118 7644 15426 7653
rect 15118 7642 15124 7644
rect 15180 7642 15204 7644
rect 15260 7642 15284 7644
rect 15340 7642 15364 7644
rect 15420 7642 15426 7644
rect 15180 7590 15182 7642
rect 15362 7590 15364 7642
rect 15118 7588 15124 7590
rect 15180 7588 15204 7590
rect 15260 7588 15284 7590
rect 15340 7588 15364 7590
rect 15420 7588 15426 7590
rect 15118 7579 15426 7588
rect 15118 6556 15426 6565
rect 15118 6554 15124 6556
rect 15180 6554 15204 6556
rect 15260 6554 15284 6556
rect 15340 6554 15364 6556
rect 15420 6554 15426 6556
rect 15180 6502 15182 6554
rect 15362 6502 15364 6554
rect 15118 6500 15124 6502
rect 15180 6500 15204 6502
rect 15260 6500 15284 6502
rect 15340 6500 15364 6502
rect 15420 6500 15426 6502
rect 15118 6491 15426 6500
rect 15488 6390 15516 7822
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15764 7206 15792 7686
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15856 6934 15884 7754
rect 15948 7274 15976 7822
rect 16040 7750 16068 8910
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15672 6322 15700 6734
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15856 6254 15884 6870
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6390 16068 6734
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 15844 6248 15896 6254
rect 16592 6225 16620 11018
rect 16684 8566 16712 12038
rect 17052 11762 17080 12922
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17236 11354 17264 15302
rect 17328 14958 17356 15982
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17420 15026 17448 15438
rect 17604 15094 17632 19306
rect 17788 18834 17816 19858
rect 17880 18970 17908 22442
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17972 21622 18000 21830
rect 18248 21706 18276 25094
rect 18340 24274 18368 25910
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18340 23866 18368 24210
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 18340 22030 18368 22714
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 18156 21678 18276 21706
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 18064 19417 18092 20198
rect 18156 19922 18184 21678
rect 18340 21146 18368 21966
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18156 19446 18184 19654
rect 18144 19440 18196 19446
rect 18050 19408 18106 19417
rect 18144 19382 18196 19388
rect 18050 19343 18106 19352
rect 18064 19310 18092 19343
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 18064 18834 18092 19246
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 17788 18426 17816 18770
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17788 17882 17816 18362
rect 18064 17882 18092 18770
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18156 16726 18184 18294
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18156 16130 18184 16662
rect 18248 16590 18276 18566
rect 18340 18426 18368 18566
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18432 17864 18460 26726
rect 18524 19938 18552 27814
rect 18660 27772 18968 27781
rect 18660 27770 18666 27772
rect 18722 27770 18746 27772
rect 18802 27770 18826 27772
rect 18882 27770 18906 27772
rect 18962 27770 18968 27772
rect 18722 27718 18724 27770
rect 18904 27718 18906 27770
rect 18660 27716 18666 27718
rect 18722 27716 18746 27718
rect 18802 27716 18826 27718
rect 18882 27716 18906 27718
rect 18962 27716 18968 27718
rect 18660 27707 18968 27716
rect 19628 27674 19656 27950
rect 19892 27872 19944 27878
rect 19892 27814 19944 27820
rect 19616 27668 19668 27674
rect 19616 27610 19668 27616
rect 19708 27600 19760 27606
rect 19708 27542 19760 27548
rect 19248 27532 19300 27538
rect 19248 27474 19300 27480
rect 19260 26994 19288 27474
rect 19616 27328 19668 27334
rect 19616 27270 19668 27276
rect 19628 27130 19656 27270
rect 19616 27124 19668 27130
rect 19616 27066 19668 27072
rect 19432 27056 19484 27062
rect 19432 26998 19484 27004
rect 19248 26988 19300 26994
rect 19168 26948 19248 26976
rect 19064 26784 19116 26790
rect 19064 26726 19116 26732
rect 18660 26684 18968 26693
rect 18660 26682 18666 26684
rect 18722 26682 18746 26684
rect 18802 26682 18826 26684
rect 18882 26682 18906 26684
rect 18962 26682 18968 26684
rect 18722 26630 18724 26682
rect 18904 26630 18906 26682
rect 18660 26628 18666 26630
rect 18722 26628 18746 26630
rect 18802 26628 18826 26630
rect 18882 26628 18906 26630
rect 18962 26628 18968 26630
rect 18660 26619 18968 26628
rect 18972 26512 19024 26518
rect 18972 26454 19024 26460
rect 18984 26314 19012 26454
rect 19076 26382 19104 26726
rect 19064 26376 19116 26382
rect 19064 26318 19116 26324
rect 18880 26308 18932 26314
rect 18880 26250 18932 26256
rect 18972 26308 19024 26314
rect 18972 26250 19024 26256
rect 18892 25974 18920 26250
rect 18880 25968 18932 25974
rect 18880 25910 18932 25916
rect 18660 25596 18968 25605
rect 18660 25594 18666 25596
rect 18722 25594 18746 25596
rect 18802 25594 18826 25596
rect 18882 25594 18906 25596
rect 18962 25594 18968 25596
rect 18722 25542 18724 25594
rect 18904 25542 18906 25594
rect 18660 25540 18666 25542
rect 18722 25540 18746 25542
rect 18802 25540 18826 25542
rect 18882 25540 18906 25542
rect 18962 25540 18968 25542
rect 18660 25531 18968 25540
rect 19076 24614 19104 26318
rect 19168 25906 19196 26948
rect 19248 26930 19300 26936
rect 19444 26518 19472 26998
rect 19720 26994 19748 27542
rect 19904 27470 19932 27814
rect 19800 27464 19852 27470
rect 19800 27406 19852 27412
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 19708 26988 19760 26994
rect 19708 26930 19760 26936
rect 19616 26852 19668 26858
rect 19616 26794 19668 26800
rect 19432 26512 19484 26518
rect 19432 26454 19484 26460
rect 19628 26382 19656 26794
rect 19812 26586 19840 27406
rect 19904 27033 19932 27406
rect 19890 27024 19946 27033
rect 19890 26959 19946 26968
rect 19800 26580 19852 26586
rect 19800 26522 19852 26528
rect 19904 26450 19932 26959
rect 19892 26444 19944 26450
rect 19892 26386 19944 26392
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19800 26376 19852 26382
rect 19800 26318 19852 26324
rect 19708 26308 19760 26314
rect 19708 26250 19760 26256
rect 19248 26240 19300 26246
rect 19248 26182 19300 26188
rect 19260 26042 19288 26182
rect 19248 26036 19300 26042
rect 19248 25978 19300 25984
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19260 25498 19288 25978
rect 19720 25906 19748 26250
rect 19708 25900 19760 25906
rect 19708 25842 19760 25848
rect 19248 25492 19300 25498
rect 19248 25434 19300 25440
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 18660 24508 18968 24517
rect 18660 24506 18666 24508
rect 18722 24506 18746 24508
rect 18802 24506 18826 24508
rect 18882 24506 18906 24508
rect 18962 24506 18968 24508
rect 18722 24454 18724 24506
rect 18904 24454 18906 24506
rect 18660 24452 18666 24454
rect 18722 24452 18746 24454
rect 18802 24452 18826 24454
rect 18882 24452 18906 24454
rect 18962 24452 18968 24454
rect 18660 24443 18968 24452
rect 19076 24206 19104 24550
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 18660 23420 18968 23429
rect 18660 23418 18666 23420
rect 18722 23418 18746 23420
rect 18802 23418 18826 23420
rect 18882 23418 18906 23420
rect 18962 23418 18968 23420
rect 18722 23366 18724 23418
rect 18904 23366 18906 23418
rect 18660 23364 18666 23366
rect 18722 23364 18746 23366
rect 18802 23364 18826 23366
rect 18882 23364 18906 23366
rect 18962 23364 18968 23366
rect 18660 23355 18968 23364
rect 19168 23322 19196 23802
rect 19156 23316 19208 23322
rect 19156 23258 19208 23264
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18984 22930 19012 23054
rect 19260 22964 19288 24346
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19352 23254 19380 23462
rect 19340 23248 19392 23254
rect 19340 23190 19392 23196
rect 19444 23118 19472 23666
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19168 22936 19288 22964
rect 19340 22976 19392 22982
rect 18984 22902 19104 22930
rect 18660 22332 18968 22341
rect 18660 22330 18666 22332
rect 18722 22330 18746 22332
rect 18802 22330 18826 22332
rect 18882 22330 18906 22332
rect 18962 22330 18968 22332
rect 18722 22278 18724 22330
rect 18904 22278 18906 22330
rect 18660 22276 18666 22278
rect 18722 22276 18746 22278
rect 18802 22276 18826 22278
rect 18882 22276 18906 22278
rect 18962 22276 18968 22278
rect 18660 22267 18968 22276
rect 19076 22234 19104 22902
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18984 21865 19012 21966
rect 19168 21962 19196 22936
rect 19340 22918 19392 22924
rect 19352 22778 19380 22918
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19260 22098 19288 22578
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19156 21956 19208 21962
rect 19156 21898 19208 21904
rect 18970 21856 19026 21865
rect 18970 21791 19026 21800
rect 18984 21706 19012 21791
rect 18984 21678 19104 21706
rect 18696 21616 18748 21622
rect 18696 21558 18748 21564
rect 18708 21418 18736 21558
rect 18696 21412 18748 21418
rect 18696 21354 18748 21360
rect 18660 21244 18968 21253
rect 18660 21242 18666 21244
rect 18722 21242 18746 21244
rect 18802 21242 18826 21244
rect 18882 21242 18906 21244
rect 18962 21242 18968 21244
rect 18722 21190 18724 21242
rect 18904 21190 18906 21242
rect 18660 21188 18666 21190
rect 18722 21188 18746 21190
rect 18802 21188 18826 21190
rect 18882 21188 18906 21190
rect 18962 21188 18968 21190
rect 18660 21179 18968 21188
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 20466 18736 20742
rect 19076 20466 19104 21678
rect 19260 20806 19288 22034
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19352 21146 19380 21354
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 19260 20262 19288 20742
rect 19248 20256 19300 20262
rect 19248 20198 19300 20204
rect 18660 20156 18968 20165
rect 18660 20154 18666 20156
rect 18722 20154 18746 20156
rect 18802 20154 18826 20156
rect 18882 20154 18906 20156
rect 18962 20154 18968 20156
rect 18722 20102 18724 20154
rect 18904 20102 18906 20154
rect 18660 20100 18666 20102
rect 18722 20100 18746 20102
rect 18802 20100 18826 20102
rect 18882 20100 18906 20102
rect 18962 20100 18968 20102
rect 18660 20091 18968 20100
rect 18524 19910 18644 19938
rect 18616 19854 18644 19910
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18660 19068 18968 19077
rect 18660 19066 18666 19068
rect 18722 19066 18746 19068
rect 18802 19066 18826 19068
rect 18882 19066 18906 19068
rect 18962 19066 18968 19068
rect 18722 19014 18724 19066
rect 18904 19014 18906 19066
rect 18660 19012 18666 19014
rect 18722 19012 18746 19014
rect 18802 19012 18826 19014
rect 18882 19012 18906 19014
rect 18962 19012 18968 19014
rect 18660 19003 18968 19012
rect 18660 17980 18968 17989
rect 18660 17978 18666 17980
rect 18722 17978 18746 17980
rect 18802 17978 18826 17980
rect 18882 17978 18906 17980
rect 18962 17978 18968 17980
rect 18722 17926 18724 17978
rect 18904 17926 18906 17978
rect 18660 17924 18666 17926
rect 18722 17924 18746 17926
rect 18802 17924 18826 17926
rect 18882 17924 18906 17926
rect 18962 17924 18968 17926
rect 18660 17915 18968 17924
rect 18696 17876 18748 17882
rect 18340 17836 18696 17864
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18248 16250 18276 16526
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18064 16102 18184 16130
rect 18064 15638 18092 16102
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17328 13258 17356 14282
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17328 11762 17356 13194
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17144 10742 17172 11086
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17328 10266 17356 11086
rect 17420 10810 17448 14962
rect 17604 11626 17632 15030
rect 17972 15026 18000 15370
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 18050 14920 18106 14929
rect 18050 14855 18052 14864
rect 18104 14855 18106 14864
rect 18052 14826 18104 14832
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17592 11620 17644 11626
rect 17592 11562 17644 11568
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16776 9926 16804 9998
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16776 8294 16804 9862
rect 17420 9722 17448 10610
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17604 9654 17632 11562
rect 17788 11354 17816 12038
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 17052 9382 17080 9522
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16960 7410 16988 8230
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16672 7336 16724 7342
rect 16670 7304 16672 7313
rect 16724 7304 16726 7313
rect 16670 7239 16726 7248
rect 17052 7206 17080 9318
rect 17604 8974 17632 9590
rect 17788 9042 17816 9862
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17236 8498 17264 8570
rect 17604 8498 17632 8774
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16776 6458 16804 6734
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 17052 6322 17080 7142
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 15844 6190 15896 6196
rect 16578 6216 16634 6225
rect 15856 5914 15884 6190
rect 16578 6151 16634 6160
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15120 5778 15148 5850
rect 16868 5778 16896 6258
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17052 5710 17080 6258
rect 17144 5914 17172 7278
rect 17236 7002 17264 7346
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15118 5468 15426 5477
rect 15118 5466 15124 5468
rect 15180 5466 15204 5468
rect 15260 5466 15284 5468
rect 15340 5466 15364 5468
rect 15420 5466 15426 5468
rect 15180 5414 15182 5466
rect 15362 5414 15364 5466
rect 15118 5412 15124 5414
rect 15180 5412 15204 5414
rect 15260 5412 15284 5414
rect 15340 5412 15364 5414
rect 15420 5412 15426 5414
rect 15118 5403 15426 5412
rect 15488 4826 15516 5578
rect 17052 5574 17080 5646
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 17052 5370 17080 5510
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15212 4622 15240 4762
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15118 4380 15426 4389
rect 15118 4378 15124 4380
rect 15180 4378 15204 4380
rect 15260 4378 15284 4380
rect 15340 4378 15364 4380
rect 15420 4378 15426 4380
rect 15180 4326 15182 4378
rect 15362 4326 15364 4378
rect 15118 4324 15124 4326
rect 15180 4324 15204 4326
rect 15260 4324 15284 4326
rect 15340 4324 15364 4326
rect 15420 4324 15426 4326
rect 15118 4315 15426 4324
rect 15948 4282 15976 5102
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15200 4208 15252 4214
rect 15200 4150 15252 4156
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 15212 3738 15240 4150
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15304 3398 15332 3878
rect 15856 3670 15884 3878
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 16592 3602 16620 3674
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16396 3528 16448 3534
rect 16394 3496 16396 3505
rect 16448 3496 16450 3505
rect 16394 3431 16450 3440
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15568 3392 15620 3398
rect 16776 3346 16804 4150
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17236 3602 17264 3878
rect 17328 3670 17356 8298
rect 17880 7546 17908 12106
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17788 6934 17816 7346
rect 17776 6928 17828 6934
rect 17776 6870 17828 6876
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17512 6662 17540 6802
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17512 5642 17540 6598
rect 17788 6186 17816 6870
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17972 5846 18000 6666
rect 18064 6644 18092 14826
rect 18156 13326 18184 15982
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18248 15162 18276 15370
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18248 10810 18276 15098
rect 18340 12918 18368 17836
rect 18696 17818 18748 17824
rect 19260 17814 19288 19858
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19248 17808 19300 17814
rect 18510 17776 18566 17785
rect 19248 17750 19300 17756
rect 18510 17711 18566 17720
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18432 16114 18460 17070
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18432 14618 18460 14962
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18524 13172 18552 17711
rect 18660 16892 18968 16901
rect 18660 16890 18666 16892
rect 18722 16890 18746 16892
rect 18802 16890 18826 16892
rect 18882 16890 18906 16892
rect 18962 16890 18968 16892
rect 18722 16838 18724 16890
rect 18904 16838 18906 16890
rect 18660 16836 18666 16838
rect 18722 16836 18746 16838
rect 18802 16836 18826 16838
rect 18882 16836 18906 16838
rect 18962 16836 18968 16838
rect 18660 16827 18968 16836
rect 19260 16810 19288 17750
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19352 17202 19380 17614
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19076 16782 19288 16810
rect 19352 16794 19380 17138
rect 19340 16788 19392 16794
rect 18604 16516 18656 16522
rect 18604 16458 18656 16464
rect 18616 16114 18644 16458
rect 19076 16114 19104 16782
rect 19340 16730 19392 16736
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18660 15804 18968 15813
rect 18660 15802 18666 15804
rect 18722 15802 18746 15804
rect 18802 15802 18826 15804
rect 18882 15802 18906 15804
rect 18962 15802 18968 15804
rect 18722 15750 18724 15802
rect 18904 15750 18906 15802
rect 18660 15748 18666 15750
rect 18722 15748 18746 15750
rect 18802 15748 18826 15750
rect 18882 15748 18906 15750
rect 18962 15748 18968 15750
rect 18660 15739 18968 15748
rect 19076 15366 19104 16050
rect 19168 16046 19196 16662
rect 19444 16572 19472 18566
rect 19536 17218 19564 25230
rect 19616 23860 19668 23866
rect 19616 23802 19668 23808
rect 19628 23118 19656 23802
rect 19597 23112 19656 23118
rect 19649 23072 19656 23112
rect 19597 23054 19649 23060
rect 19720 22982 19748 25842
rect 19812 25770 19840 26318
rect 19904 25838 19932 26386
rect 19892 25832 19944 25838
rect 19892 25774 19944 25780
rect 19800 25764 19852 25770
rect 19800 25706 19852 25712
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19812 24614 19840 25230
rect 19800 24608 19852 24614
rect 19800 24550 19852 24556
rect 19812 24206 19840 24550
rect 19800 24200 19852 24206
rect 19800 24142 19852 24148
rect 19812 23662 19840 24142
rect 19996 24070 20024 28358
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19800 23656 19852 23662
rect 19800 23598 19852 23604
rect 19708 22976 19760 22982
rect 19708 22918 19760 22924
rect 19616 22500 19668 22506
rect 19616 22442 19668 22448
rect 19628 22030 19656 22442
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19708 21956 19760 21962
rect 19708 21898 19760 21904
rect 19720 21690 19748 21898
rect 19708 21684 19760 21690
rect 19708 21626 19760 21632
rect 19536 17190 19748 17218
rect 19616 16584 19668 16590
rect 19444 16544 19616 16572
rect 19616 16526 19668 16532
rect 19248 16516 19300 16522
rect 19248 16458 19300 16464
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 18660 14716 18968 14725
rect 18660 14714 18666 14716
rect 18722 14714 18746 14716
rect 18802 14714 18826 14716
rect 18882 14714 18906 14716
rect 18962 14714 18968 14716
rect 18722 14662 18724 14714
rect 18904 14662 18906 14714
rect 18660 14660 18666 14662
rect 18722 14660 18746 14662
rect 18802 14660 18826 14662
rect 18882 14660 18906 14662
rect 18962 14660 18968 14662
rect 18660 14651 18968 14660
rect 18660 13628 18968 13637
rect 18660 13626 18666 13628
rect 18722 13626 18746 13628
rect 18802 13626 18826 13628
rect 18882 13626 18906 13628
rect 18962 13626 18968 13628
rect 18722 13574 18724 13626
rect 18904 13574 18906 13626
rect 18660 13572 18666 13574
rect 18722 13572 18746 13574
rect 18802 13572 18826 13574
rect 18882 13572 18906 13574
rect 18962 13572 18968 13574
rect 18660 13563 18968 13572
rect 18432 13144 18552 13172
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18340 12714 18368 12854
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18432 12345 18460 13144
rect 19076 12986 19104 15302
rect 19260 14618 19288 16458
rect 19628 15978 19656 16526
rect 19616 15972 19668 15978
rect 19616 15914 19668 15920
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19352 13462 19380 13806
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19352 12866 19380 13398
rect 19260 12850 19380 12866
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 19248 12844 19380 12850
rect 19300 12838 19380 12844
rect 19248 12786 19300 12792
rect 18524 12646 18552 12786
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18524 12442 18552 12582
rect 18660 12540 18968 12549
rect 18660 12538 18666 12540
rect 18722 12538 18746 12540
rect 18802 12538 18826 12540
rect 18882 12538 18906 12540
rect 18962 12538 18968 12540
rect 18722 12486 18724 12538
rect 18904 12486 18906 12538
rect 18660 12484 18666 12486
rect 18722 12484 18746 12486
rect 18802 12484 18826 12486
rect 18882 12484 18906 12486
rect 18962 12484 18968 12486
rect 18660 12475 18968 12484
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18418 12336 18474 12345
rect 18418 12271 18474 12280
rect 18432 11898 18460 12271
rect 18524 12102 18552 12378
rect 19352 12238 19380 12838
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19536 12238 19564 12378
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18524 11830 18552 12038
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18432 11234 18460 11698
rect 18524 11354 18552 11766
rect 19260 11762 19288 12038
rect 19352 11898 19380 12038
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 18660 11452 18968 11461
rect 18660 11450 18666 11452
rect 18722 11450 18746 11452
rect 18802 11450 18826 11452
rect 18882 11450 18906 11452
rect 18962 11450 18968 11452
rect 18722 11398 18724 11450
rect 18904 11398 18906 11450
rect 18660 11396 18666 11398
rect 18722 11396 18746 11398
rect 18802 11396 18826 11398
rect 18882 11396 18906 11398
rect 18962 11396 18968 11398
rect 18660 11387 18968 11396
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 19168 11286 19196 11630
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19156 11280 19208 11286
rect 18432 11218 18552 11234
rect 19156 11222 19208 11228
rect 18432 11212 18564 11218
rect 18432 11206 18512 11212
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18326 10704 18382 10713
rect 18326 10639 18382 10648
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 6798 18276 7686
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18064 6616 18276 6644
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17788 4758 17816 5510
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17788 4214 17816 4694
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 17788 4078 17816 4150
rect 17972 4146 18000 5782
rect 18064 5370 18092 6326
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 18064 4214 18092 5306
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17316 3664 17368 3670
rect 17316 3606 17368 3612
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17880 3534 17908 3878
rect 17684 3528 17736 3534
rect 17682 3496 17684 3505
rect 17868 3528 17920 3534
rect 17736 3496 17738 3505
rect 17868 3470 17920 3476
rect 17972 3466 18000 3878
rect 17682 3431 17738 3440
rect 17960 3460 18012 3466
rect 15568 3334 15620 3340
rect 15118 3292 15426 3301
rect 15118 3290 15124 3292
rect 15180 3290 15204 3292
rect 15260 3290 15284 3292
rect 15340 3290 15364 3292
rect 15420 3290 15426 3292
rect 15180 3238 15182 3290
rect 15362 3238 15364 3290
rect 15118 3236 15124 3238
rect 15180 3236 15204 3238
rect 15260 3236 15284 3238
rect 15340 3236 15364 3238
rect 15420 3236 15426 3238
rect 15118 3227 15426 3236
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 15580 2922 15608 3334
rect 16592 3318 16804 3346
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 14936 2446 14964 2586
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 16592 2378 16620 3318
rect 17696 3194 17724 3431
rect 17960 3402 18012 3408
rect 18064 3398 18092 4150
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16776 2378 16804 2790
rect 18064 2774 18092 3334
rect 18156 3058 18184 3606
rect 18248 3058 18276 6616
rect 18340 6322 18368 10639
rect 18432 6458 18460 11206
rect 18512 11154 18564 11160
rect 19168 11150 19196 11222
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19260 10742 19288 11562
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 18660 10364 18968 10373
rect 18660 10362 18666 10364
rect 18722 10362 18746 10364
rect 18802 10362 18826 10364
rect 18882 10362 18906 10364
rect 18962 10362 18968 10364
rect 18722 10310 18724 10362
rect 18904 10310 18906 10362
rect 18660 10308 18666 10310
rect 18722 10308 18746 10310
rect 18802 10308 18826 10310
rect 18882 10308 18906 10310
rect 18962 10308 18968 10310
rect 18660 10299 18968 10308
rect 19352 10062 19380 10950
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19340 10056 19392 10062
rect 19338 10024 19340 10033
rect 19392 10024 19394 10033
rect 19338 9959 19394 9968
rect 19444 9926 19472 10610
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 18708 9654 18736 9862
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18660 9276 18968 9285
rect 18660 9274 18666 9276
rect 18722 9274 18746 9276
rect 18802 9274 18826 9276
rect 18882 9274 18906 9276
rect 18962 9274 18968 9276
rect 18722 9222 18724 9274
rect 18904 9222 18906 9274
rect 18660 9220 18666 9222
rect 18722 9220 18746 9222
rect 18802 9220 18826 9222
rect 18882 9220 18906 9222
rect 18962 9220 18968 9222
rect 18660 9211 18968 9220
rect 18660 8188 18968 8197
rect 18660 8186 18666 8188
rect 18722 8186 18746 8188
rect 18802 8186 18826 8188
rect 18882 8186 18906 8188
rect 18962 8186 18968 8188
rect 18722 8134 18724 8186
rect 18904 8134 18906 8186
rect 18660 8132 18666 8134
rect 18722 8132 18746 8134
rect 18802 8132 18826 8134
rect 18882 8132 18906 8134
rect 18962 8132 18968 8134
rect 18660 8123 18968 8132
rect 19444 7886 19472 9862
rect 19628 9654 19656 15642
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19432 7880 19484 7886
rect 19484 7840 19564 7868
rect 19432 7822 19484 7828
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19444 7410 19472 7686
rect 19536 7546 19564 7840
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19628 7410 19656 8026
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 18616 7290 18644 7346
rect 18524 7262 18644 7290
rect 18524 7002 18552 7262
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 18660 7100 18968 7109
rect 18660 7098 18666 7100
rect 18722 7098 18746 7100
rect 18802 7098 18826 7100
rect 18882 7098 18906 7100
rect 18962 7098 18968 7100
rect 18722 7046 18724 7098
rect 18904 7046 18906 7098
rect 18660 7044 18666 7046
rect 18722 7044 18746 7046
rect 18802 7044 18826 7046
rect 18882 7044 18906 7046
rect 18962 7044 18968 7046
rect 18660 7035 18968 7044
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18340 5370 18368 6258
rect 18524 5778 18552 6802
rect 19352 6798 19380 7142
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 18616 6458 18644 6734
rect 19260 6458 19288 6734
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19064 6248 19116 6254
rect 19116 6196 19196 6202
rect 19064 6190 19196 6196
rect 19076 6174 19196 6190
rect 18660 6012 18968 6021
rect 18660 6010 18666 6012
rect 18722 6010 18746 6012
rect 18802 6010 18826 6012
rect 18882 6010 18906 6012
rect 18962 6010 18968 6012
rect 18722 5958 18724 6010
rect 18904 5958 18906 6010
rect 18660 5956 18666 5958
rect 18722 5956 18746 5958
rect 18802 5956 18826 5958
rect 18882 5956 18906 5958
rect 18962 5956 18968 5958
rect 18660 5947 18968 5956
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 19168 5030 19196 6174
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19260 5030 19288 6054
rect 19352 5778 19380 6326
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19444 5710 19472 7346
rect 19522 6896 19578 6905
rect 19522 6831 19524 6840
rect 19576 6831 19578 6840
rect 19524 6802 19576 6808
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19524 6724 19576 6730
rect 19524 6666 19576 6672
rect 19536 5914 19564 6666
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19628 5778 19656 6734
rect 19616 5772 19668 5778
rect 19616 5714 19668 5720
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 18660 4924 18968 4933
rect 18660 4922 18666 4924
rect 18722 4922 18746 4924
rect 18802 4922 18826 4924
rect 18882 4922 18906 4924
rect 18962 4922 18968 4924
rect 18722 4870 18724 4922
rect 18904 4870 18906 4922
rect 18660 4868 18666 4870
rect 18722 4868 18746 4870
rect 18802 4868 18826 4870
rect 18882 4868 18906 4870
rect 18962 4868 18968 4870
rect 18660 4859 18968 4868
rect 19168 4690 19196 4966
rect 19260 4826 19288 4966
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 18660 3836 18968 3845
rect 18660 3834 18666 3836
rect 18722 3834 18746 3836
rect 18802 3834 18826 3836
rect 18882 3834 18906 3836
rect 18962 3834 18968 3836
rect 18722 3782 18724 3834
rect 18904 3782 18906 3834
rect 18660 3780 18666 3782
rect 18722 3780 18746 3782
rect 18802 3780 18826 3782
rect 18882 3780 18906 3782
rect 18962 3780 18968 3782
rect 18660 3771 18968 3780
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 18984 3126 19012 3470
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18064 2746 18276 2774
rect 18248 2514 18276 2746
rect 18660 2748 18968 2757
rect 18660 2746 18666 2748
rect 18722 2746 18746 2748
rect 18802 2746 18826 2748
rect 18882 2746 18906 2748
rect 18962 2746 18968 2748
rect 18722 2694 18724 2746
rect 18904 2694 18906 2746
rect 18660 2692 18666 2694
rect 18722 2692 18746 2694
rect 18802 2692 18826 2694
rect 18882 2692 18906 2694
rect 18962 2692 18968 2694
rect 18660 2683 18968 2692
rect 19168 2514 19196 4626
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19352 4010 19380 4490
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 19260 2446 19288 2790
rect 19720 2774 19748 17190
rect 19628 2746 19748 2774
rect 19628 2650 19656 2746
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 19812 2514 19840 23598
rect 19892 23520 19944 23526
rect 19892 23462 19944 23468
rect 19904 23322 19932 23462
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 19996 23118 20024 24006
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19892 22432 19944 22438
rect 19892 22374 19944 22380
rect 19904 22098 19932 22374
rect 19892 22092 19944 22098
rect 19892 22034 19944 22040
rect 19904 21418 19932 22034
rect 19892 21412 19944 21418
rect 19892 21354 19944 21360
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19904 20262 19932 20402
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 19904 18698 19932 20198
rect 19996 19378 20024 23054
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19892 18692 19944 18698
rect 19892 18634 19944 18640
rect 19904 18086 19932 18634
rect 19996 18358 20024 19314
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19904 15706 19932 18022
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19904 13938 19932 14418
rect 20088 14278 20116 29990
rect 20168 29640 20220 29646
rect 20168 29582 20220 29588
rect 20180 28082 20208 29582
rect 22020 29170 22048 29990
rect 22100 29844 22152 29850
rect 22100 29786 22152 29792
rect 21456 29164 21508 29170
rect 21456 29106 21508 29112
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 21468 28994 21496 29106
rect 21376 28966 21496 28994
rect 21272 28960 21324 28966
rect 21272 28902 21324 28908
rect 21284 28626 21312 28902
rect 21272 28620 21324 28626
rect 21272 28562 21324 28568
rect 21272 28416 21324 28422
rect 21272 28358 21324 28364
rect 20720 28212 20772 28218
rect 20720 28154 20772 28160
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 20168 27872 20220 27878
rect 20168 27814 20220 27820
rect 20180 27334 20208 27814
rect 20444 27464 20496 27470
rect 20444 27406 20496 27412
rect 20168 27328 20220 27334
rect 20168 27270 20220 27276
rect 20456 27130 20484 27406
rect 20444 27124 20496 27130
rect 20444 27066 20496 27072
rect 20352 27056 20404 27062
rect 20166 27024 20222 27033
rect 20352 26998 20404 27004
rect 20166 26959 20168 26968
rect 20220 26959 20222 26968
rect 20260 26988 20312 26994
rect 20168 26930 20220 26936
rect 20260 26930 20312 26936
rect 20272 26042 20300 26930
rect 20364 26518 20392 26998
rect 20352 26512 20404 26518
rect 20352 26454 20404 26460
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20260 26036 20312 26042
rect 20260 25978 20312 25984
rect 20456 25974 20484 26318
rect 20444 25968 20496 25974
rect 20444 25910 20496 25916
rect 20732 23594 20760 28154
rect 21284 28082 21312 28358
rect 21376 28150 21404 28966
rect 21824 28620 21876 28626
rect 21824 28562 21876 28568
rect 21364 28144 21416 28150
rect 21364 28086 21416 28092
rect 21548 28144 21600 28150
rect 21548 28086 21600 28092
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 20996 27328 21048 27334
rect 20996 27270 21048 27276
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20824 26042 20852 26318
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 20916 25906 20944 26862
rect 21008 26586 21036 27270
rect 21284 27062 21312 28018
rect 21272 27056 21324 27062
rect 21272 26998 21324 27004
rect 21272 26920 21324 26926
rect 21376 26908 21404 28086
rect 21560 27606 21588 28086
rect 21732 27940 21784 27946
rect 21732 27882 21784 27888
rect 21744 27606 21772 27882
rect 21548 27600 21600 27606
rect 21548 27542 21600 27548
rect 21732 27600 21784 27606
rect 21732 27542 21784 27548
rect 21324 26880 21404 26908
rect 21272 26862 21324 26868
rect 20996 26580 21048 26586
rect 20996 26522 21048 26528
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 20916 25498 20944 25842
rect 20904 25492 20956 25498
rect 20824 25452 20904 25480
rect 20824 23866 20852 25452
rect 20904 25434 20956 25440
rect 21284 25226 21312 26862
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21560 26518 21588 26726
rect 21548 26512 21600 26518
rect 21548 26454 21600 26460
rect 21364 26240 21416 26246
rect 21364 26182 21416 26188
rect 21376 25974 21404 26182
rect 21364 25968 21416 25974
rect 21364 25910 21416 25916
rect 21376 25498 21404 25910
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 20996 25220 21048 25226
rect 20996 25162 21048 25168
rect 21272 25220 21324 25226
rect 21272 25162 21324 25168
rect 20904 24132 20956 24138
rect 20904 24074 20956 24080
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 20720 23588 20772 23594
rect 20720 23530 20772 23536
rect 20824 23322 20852 23802
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20824 22778 20852 23258
rect 20916 23118 20944 24074
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20916 21554 20944 21830
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20824 21010 20852 21490
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20824 20482 20852 20946
rect 20916 20534 20944 21286
rect 20732 20454 20852 20482
rect 20904 20528 20956 20534
rect 20904 20470 20956 20476
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20640 19854 20668 20198
rect 20732 19922 20760 20454
rect 20812 20392 20864 20398
rect 21008 20380 21036 25162
rect 21836 24818 21864 28562
rect 22112 28558 22140 29786
rect 22664 29646 22692 30058
rect 24400 30048 24452 30054
rect 24400 29990 24452 29996
rect 22836 29708 22888 29714
rect 22836 29650 22888 29656
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22202 29404 22510 29413
rect 22202 29402 22208 29404
rect 22264 29402 22288 29404
rect 22344 29402 22368 29404
rect 22424 29402 22448 29404
rect 22504 29402 22510 29404
rect 22264 29350 22266 29402
rect 22446 29350 22448 29402
rect 22202 29348 22208 29350
rect 22264 29348 22288 29350
rect 22344 29348 22368 29350
rect 22424 29348 22448 29350
rect 22504 29348 22510 29350
rect 22202 29339 22510 29348
rect 22664 29170 22692 29582
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 22560 28416 22612 28422
rect 22560 28358 22612 28364
rect 22202 28316 22510 28325
rect 22202 28314 22208 28316
rect 22264 28314 22288 28316
rect 22344 28314 22368 28316
rect 22424 28314 22448 28316
rect 22504 28314 22510 28316
rect 22264 28262 22266 28314
rect 22446 28262 22448 28314
rect 22202 28260 22208 28262
rect 22264 28260 22288 28262
rect 22344 28260 22368 28262
rect 22424 28260 22448 28262
rect 22504 28260 22510 28262
rect 22202 28251 22510 28260
rect 22572 28082 22600 28358
rect 22664 28150 22692 29106
rect 22848 28966 22876 29650
rect 22836 28960 22888 28966
rect 22836 28902 22888 28908
rect 23020 28960 23072 28966
rect 23020 28902 23072 28908
rect 23756 28960 23808 28966
rect 23756 28902 23808 28908
rect 22652 28144 22704 28150
rect 22652 28086 22704 28092
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 22112 26234 22140 28018
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22652 27396 22704 27402
rect 22652 27338 22704 27344
rect 22202 27228 22510 27237
rect 22202 27226 22208 27228
rect 22264 27226 22288 27228
rect 22344 27226 22368 27228
rect 22424 27226 22448 27228
rect 22504 27226 22510 27228
rect 22264 27174 22266 27226
rect 22446 27174 22448 27226
rect 22202 27172 22208 27174
rect 22264 27172 22288 27174
rect 22344 27172 22368 27174
rect 22424 27172 22448 27174
rect 22504 27172 22510 27174
rect 22202 27163 22510 27172
rect 22192 26852 22244 26858
rect 22192 26794 22244 26800
rect 22204 26450 22232 26794
rect 22376 26784 22428 26790
rect 22376 26726 22428 26732
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22388 26586 22416 26726
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 22192 26444 22244 26450
rect 22192 26386 22244 26392
rect 22572 26353 22600 26726
rect 22664 26489 22692 27338
rect 22756 26994 22784 27814
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22650 26480 22706 26489
rect 22650 26415 22706 26424
rect 22558 26344 22614 26353
rect 22558 26279 22614 26288
rect 22020 26206 22140 26234
rect 22020 25362 22048 26206
rect 22202 26140 22510 26149
rect 22202 26138 22208 26140
rect 22264 26138 22288 26140
rect 22344 26138 22368 26140
rect 22424 26138 22448 26140
rect 22504 26138 22510 26140
rect 22264 26086 22266 26138
rect 22446 26086 22448 26138
rect 22202 26084 22208 26086
rect 22264 26084 22288 26086
rect 22344 26084 22368 26086
rect 22424 26084 22448 26086
rect 22504 26084 22510 26086
rect 22202 26075 22510 26084
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21836 24206 21864 24754
rect 22020 24274 22048 25298
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22202 25052 22510 25061
rect 22202 25050 22208 25052
rect 22264 25050 22288 25052
rect 22344 25050 22368 25052
rect 22424 25050 22448 25052
rect 22504 25050 22510 25052
rect 22264 24998 22266 25050
rect 22446 24998 22448 25050
rect 22202 24996 22208 24998
rect 22264 24996 22288 24998
rect 22344 24996 22368 24998
rect 22424 24996 22448 24998
rect 22504 24996 22510 24998
rect 22202 24987 22510 24996
rect 22572 24954 22600 25230
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22008 24268 22060 24274
rect 22008 24210 22060 24216
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21836 23866 21864 24142
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 21732 23792 21784 23798
rect 21732 23734 21784 23740
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 21088 23180 21140 23186
rect 21088 23122 21140 23128
rect 21100 22982 21128 23122
rect 21192 23118 21220 23462
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21088 22976 21140 22982
rect 21086 22944 21088 22953
rect 21140 22944 21142 22953
rect 21086 22879 21142 22888
rect 21088 22704 21140 22710
rect 21088 22646 21140 22652
rect 21100 22022 21128 22646
rect 21192 22137 21220 23054
rect 21272 23044 21324 23050
rect 21272 22986 21324 22992
rect 21178 22128 21234 22137
rect 21178 22063 21234 22072
rect 21180 22024 21232 22030
rect 21100 21994 21180 22022
rect 21100 21010 21128 21994
rect 21180 21966 21232 21972
rect 21178 21856 21234 21865
rect 21178 21791 21234 21800
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 20864 20352 21036 20380
rect 20812 20334 20864 20340
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20536 19780 20588 19786
rect 20536 19722 20588 19728
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20364 19514 20392 19654
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20456 19122 20484 19382
rect 20548 19310 20576 19722
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20456 19094 20576 19122
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 18290 20392 18566
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20364 16114 20392 16730
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20258 16008 20314 16017
rect 20258 15943 20314 15952
rect 20272 15706 20300 15943
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20272 15026 20300 15642
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 20088 12646 20116 14214
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20272 13462 20300 13806
rect 20260 13456 20312 13462
rect 20260 13398 20312 13404
rect 20272 13002 20300 13398
rect 20180 12986 20300 13002
rect 20180 12980 20312 12986
rect 20180 12974 20260 12980
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19904 11354 19932 11630
rect 20088 11558 20116 12378
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20088 11354 20116 11494
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20088 11150 20116 11290
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19904 9674 19932 11018
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19996 10266 20024 10542
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19904 9646 20024 9674
rect 19996 7954 20024 9646
rect 20076 8560 20128 8566
rect 20074 8528 20076 8537
rect 20128 8528 20130 8537
rect 20074 8463 20130 8472
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19996 7750 20024 7890
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19996 6905 20024 7686
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 19982 6896 20038 6905
rect 19982 6831 20038 6840
rect 19892 6452 19944 6458
rect 19892 6394 19944 6400
rect 19904 6186 19932 6394
rect 19996 6254 20024 6831
rect 20088 6322 20116 7482
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19892 6180 19944 6186
rect 19892 6122 19944 6128
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20088 3738 20116 4558
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20180 2774 20208 12974
rect 20260 12922 20312 12928
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20272 12442 20300 12582
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20364 10538 20392 16050
rect 20548 15978 20576 19094
rect 20640 18850 20668 19790
rect 20732 18970 20760 19858
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20640 18834 20760 18850
rect 20640 18828 20772 18834
rect 20640 18822 20720 18828
rect 20720 18770 20772 18776
rect 20732 18057 20760 18770
rect 20824 18766 20852 20334
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20824 18358 20852 18702
rect 21008 18630 21036 19790
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20916 18290 20944 18566
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20718 18048 20774 18057
rect 20718 17983 20774 17992
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20732 16726 20760 17138
rect 20720 16720 20772 16726
rect 20626 16688 20682 16697
rect 20720 16662 20772 16668
rect 20626 16623 20682 16632
rect 20640 16590 20668 16623
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20548 13954 20576 15914
rect 20824 15314 20852 18158
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20732 15286 20852 15314
rect 20628 14884 20680 14890
rect 20628 14826 20680 14832
rect 20640 14657 20668 14826
rect 20626 14648 20682 14657
rect 20626 14583 20682 14592
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20640 14074 20668 14418
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20444 13932 20496 13938
rect 20548 13926 20668 13954
rect 20444 13874 20496 13880
rect 20456 13734 20484 13874
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20456 13394 20484 13670
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20352 10532 20404 10538
rect 20352 10474 20404 10480
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20272 4826 20300 8434
rect 20456 8378 20484 11698
rect 20548 8498 20576 13126
rect 20640 10810 20668 13926
rect 20732 11898 20760 15286
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20824 14346 20852 15030
rect 20916 14414 20944 16594
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20824 14074 20852 14282
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20824 12986 20852 13806
rect 20902 13016 20958 13025
rect 20812 12980 20864 12986
rect 20902 12951 20958 12960
rect 20812 12922 20864 12928
rect 20916 12918 20944 12951
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 20812 12164 20864 12170
rect 20812 12106 20864 12112
rect 20824 11898 20852 12106
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20824 11762 20852 11834
rect 20916 11762 20944 12650
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20732 10266 20760 10542
rect 20824 10470 20852 10746
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20640 9382 20668 9998
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20732 9722 20760 9930
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20824 9586 20852 10406
rect 20916 9994 20944 10406
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20916 9586 20944 9930
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20640 9110 20668 9318
rect 20628 9104 20680 9110
rect 20628 9046 20680 9052
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20456 8350 20668 8378
rect 20352 7812 20404 7818
rect 20352 7754 20404 7760
rect 20364 7410 20392 7754
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20456 6798 20484 7414
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20456 6322 20484 6734
rect 20548 6458 20576 6734
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20548 6186 20576 6394
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20548 4690 20576 5714
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 20640 4622 20668 8350
rect 20824 7392 20852 9522
rect 20916 9382 20944 9522
rect 21008 9489 21036 18566
rect 21100 18086 21128 18838
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 21192 17134 21220 21791
rect 21284 17338 21312 22986
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 21364 22092 21416 22098
rect 21351 22040 21364 22080
rect 21351 22034 21416 22040
rect 21351 21978 21379 22034
rect 21351 21950 21404 21978
rect 21376 21690 21404 21950
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21376 20874 21404 21286
rect 21560 21026 21588 22578
rect 21640 22092 21692 22098
rect 21640 22034 21692 22040
rect 21652 21486 21680 22034
rect 21744 21554 21772 23734
rect 21836 23118 21864 23802
rect 22020 23798 22048 24210
rect 22100 24064 22152 24070
rect 22100 24006 22152 24012
rect 22112 23798 22140 24006
rect 22202 23964 22510 23973
rect 22202 23962 22208 23964
rect 22264 23962 22288 23964
rect 22344 23962 22368 23964
rect 22424 23962 22448 23964
rect 22504 23962 22510 23964
rect 22264 23910 22266 23962
rect 22446 23910 22448 23962
rect 22202 23908 22208 23910
rect 22264 23908 22288 23910
rect 22344 23908 22368 23910
rect 22424 23908 22448 23910
rect 22504 23908 22510 23910
rect 22202 23899 22510 23908
rect 22008 23792 22060 23798
rect 22008 23734 22060 23740
rect 22100 23792 22152 23798
rect 22100 23734 22152 23740
rect 22560 23792 22612 23798
rect 22560 23734 22612 23740
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 21836 22642 21864 23054
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21916 22500 21968 22506
rect 21916 22442 21968 22448
rect 21824 22160 21876 22166
rect 21824 22102 21876 22108
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21560 20998 21680 21026
rect 21652 20942 21680 20998
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21364 20868 21416 20874
rect 21364 20810 21416 20816
rect 21376 19174 21404 20810
rect 21652 20466 21680 20878
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21376 18698 21404 19110
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21468 18290 21496 18702
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21284 15162 21312 17274
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21376 16114 21404 16526
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21376 15502 21404 16050
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 21100 14346 21128 14894
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21100 12850 21128 14010
rect 21192 13326 21220 14214
rect 21284 13938 21312 15098
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21272 13796 21324 13802
rect 21272 13738 21324 13744
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21284 11218 21312 13738
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21376 12714 21404 13262
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21284 10674 21312 11154
rect 21468 10674 21496 18226
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21560 10810 21588 17546
rect 21652 16998 21680 20266
rect 21836 19854 21864 22102
rect 21928 22094 21956 22442
rect 22020 22234 22048 22918
rect 22202 22876 22510 22885
rect 22202 22874 22208 22876
rect 22264 22874 22288 22876
rect 22344 22874 22368 22876
rect 22424 22874 22448 22876
rect 22504 22874 22510 22876
rect 22264 22822 22266 22874
rect 22446 22822 22448 22874
rect 22202 22820 22208 22822
rect 22264 22820 22288 22822
rect 22344 22820 22368 22822
rect 22424 22820 22448 22822
rect 22504 22820 22510 22822
rect 22202 22811 22510 22820
rect 22572 22642 22600 23734
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 22008 22094 22060 22098
rect 21928 22092 22060 22094
rect 21928 22066 22008 22092
rect 22008 22034 22060 22040
rect 22202 21788 22510 21797
rect 22202 21786 22208 21788
rect 22264 21786 22288 21788
rect 22344 21786 22368 21788
rect 22424 21786 22448 21788
rect 22504 21786 22510 21788
rect 22264 21734 22266 21786
rect 22446 21734 22448 21786
rect 22202 21732 22208 21734
rect 22264 21732 22288 21734
rect 22344 21732 22368 21734
rect 22424 21732 22448 21734
rect 22504 21732 22510 21734
rect 22202 21723 22510 21732
rect 22560 21412 22612 21418
rect 22560 21354 22612 21360
rect 22202 20700 22510 20709
rect 22202 20698 22208 20700
rect 22264 20698 22288 20700
rect 22344 20698 22368 20700
rect 22424 20698 22448 20700
rect 22504 20698 22510 20700
rect 22264 20646 22266 20698
rect 22446 20646 22448 20698
rect 22202 20644 22208 20646
rect 22264 20644 22288 20646
rect 22344 20644 22368 20646
rect 22424 20644 22448 20646
rect 22504 20644 22510 20646
rect 22202 20635 22510 20644
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 22202 19612 22510 19621
rect 22202 19610 22208 19612
rect 22264 19610 22288 19612
rect 22344 19610 22368 19612
rect 22424 19610 22448 19612
rect 22504 19610 22510 19612
rect 22264 19558 22266 19610
rect 22446 19558 22448 19610
rect 22202 19556 22208 19558
rect 22264 19556 22288 19558
rect 22344 19556 22368 19558
rect 22424 19556 22448 19558
rect 22504 19556 22510 19558
rect 22202 19547 22510 19556
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21744 17678 21772 18906
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21744 17202 21772 17478
rect 21732 17196 21784 17202
rect 21732 17138 21784 17144
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21652 15026 21680 16934
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21638 14648 21694 14657
rect 21638 14583 21694 14592
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21652 10169 21680 14583
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21744 14346 21772 14418
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 21836 13802 21864 18566
rect 22202 18524 22510 18533
rect 22202 18522 22208 18524
rect 22264 18522 22288 18524
rect 22344 18522 22368 18524
rect 22424 18522 22448 18524
rect 22504 18522 22510 18524
rect 22264 18470 22266 18522
rect 22446 18470 22448 18522
rect 22202 18468 22208 18470
rect 22264 18468 22288 18470
rect 22344 18468 22368 18470
rect 22424 18468 22448 18470
rect 22504 18468 22510 18470
rect 22202 18459 22510 18468
rect 22202 17436 22510 17445
rect 22202 17434 22208 17436
rect 22264 17434 22288 17436
rect 22344 17434 22368 17436
rect 22424 17434 22448 17436
rect 22504 17434 22510 17436
rect 22264 17382 22266 17434
rect 22446 17382 22448 17434
rect 22202 17380 22208 17382
rect 22264 17380 22288 17382
rect 22344 17380 22368 17382
rect 22424 17380 22448 17382
rect 22504 17380 22510 17382
rect 22202 17371 22510 17380
rect 22008 17332 22060 17338
rect 22008 17274 22060 17280
rect 22020 17202 22048 17274
rect 22572 17202 22600 21354
rect 22664 17218 22692 26415
rect 22744 25764 22796 25770
rect 22744 25706 22796 25712
rect 22756 24206 22784 25706
rect 22848 25362 22876 28902
rect 23032 28558 23060 28902
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 23204 28484 23256 28490
rect 23204 28426 23256 28432
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 23216 28218 23244 28426
rect 23204 28212 23256 28218
rect 23204 28154 23256 28160
rect 23112 28144 23164 28150
rect 23112 28086 23164 28092
rect 23124 26518 23152 28086
rect 23216 27470 23244 28154
rect 23676 28082 23704 28426
rect 23768 28422 23796 28902
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23664 28076 23716 28082
rect 23664 28018 23716 28024
rect 23492 27878 23520 28018
rect 23480 27872 23532 27878
rect 23480 27814 23532 27820
rect 23676 27470 23704 28018
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23296 26784 23348 26790
rect 23296 26726 23348 26732
rect 23112 26512 23164 26518
rect 23112 26454 23164 26460
rect 23124 25498 23152 26454
rect 23308 25770 23336 26726
rect 23676 26586 23704 27406
rect 23572 26580 23624 26586
rect 23572 26522 23624 26528
rect 23664 26580 23716 26586
rect 23664 26522 23716 26528
rect 23584 26042 23612 26522
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23296 25764 23348 25770
rect 23296 25706 23348 25712
rect 23308 25498 23336 25706
rect 23112 25492 23164 25498
rect 23112 25434 23164 25440
rect 23296 25492 23348 25498
rect 23296 25434 23348 25440
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 23388 25220 23440 25226
rect 23388 25162 23440 25168
rect 22928 25152 22980 25158
rect 22928 25094 22980 25100
rect 22940 24886 22968 25094
rect 22928 24880 22980 24886
rect 22980 24840 23060 24868
rect 22928 24822 22980 24828
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 22928 23724 22980 23730
rect 22928 23666 22980 23672
rect 22940 23526 22968 23666
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22744 23316 22796 23322
rect 22744 23258 22796 23264
rect 22756 22506 22784 23258
rect 22836 22636 22888 22642
rect 22940 22624 22968 23462
rect 22888 22596 22968 22624
rect 22836 22578 22888 22584
rect 22744 22500 22796 22506
rect 22744 22442 22796 22448
rect 22756 21962 22784 22442
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22744 20052 22796 20058
rect 22744 19994 22796 20000
rect 22756 19854 22784 19994
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22836 19712 22888 19718
rect 22836 19654 22888 19660
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 22560 17196 22612 17202
rect 22664 17190 22784 17218
rect 22560 17138 22612 17144
rect 22572 16522 22600 17138
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 22112 12374 22140 16390
rect 22202 16348 22510 16357
rect 22202 16346 22208 16348
rect 22264 16346 22288 16348
rect 22344 16346 22368 16348
rect 22424 16346 22448 16348
rect 22504 16346 22510 16348
rect 22264 16294 22266 16346
rect 22446 16294 22448 16346
rect 22202 16292 22208 16294
rect 22264 16292 22288 16294
rect 22344 16292 22368 16294
rect 22424 16292 22448 16294
rect 22504 16292 22510 16294
rect 22202 16283 22510 16292
rect 22202 15260 22510 15269
rect 22202 15258 22208 15260
rect 22264 15258 22288 15260
rect 22344 15258 22368 15260
rect 22424 15258 22448 15260
rect 22504 15258 22510 15260
rect 22264 15206 22266 15258
rect 22446 15206 22448 15258
rect 22202 15204 22208 15206
rect 22264 15204 22288 15206
rect 22344 15204 22368 15206
rect 22424 15204 22448 15206
rect 22504 15204 22510 15206
rect 22202 15195 22510 15204
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22202 14172 22510 14181
rect 22202 14170 22208 14172
rect 22264 14170 22288 14172
rect 22344 14170 22368 14172
rect 22424 14170 22448 14172
rect 22504 14170 22510 14172
rect 22264 14118 22266 14170
rect 22446 14118 22448 14170
rect 22202 14116 22208 14118
rect 22264 14116 22288 14118
rect 22344 14116 22368 14118
rect 22424 14116 22448 14118
rect 22504 14116 22510 14118
rect 22202 14107 22510 14116
rect 22572 13326 22600 14214
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22202 13084 22510 13093
rect 22202 13082 22208 13084
rect 22264 13082 22288 13084
rect 22344 13082 22368 13084
rect 22424 13082 22448 13084
rect 22504 13082 22510 13084
rect 22264 13030 22266 13082
rect 22446 13030 22448 13082
rect 22202 13028 22208 13030
rect 22264 13028 22288 13030
rect 22344 13028 22368 13030
rect 22424 13028 22448 13030
rect 22504 13028 22510 13030
rect 22202 13019 22510 13028
rect 22100 12368 22152 12374
rect 22100 12310 22152 12316
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21928 10266 21956 10610
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 21638 10160 21694 10169
rect 21638 10095 21694 10104
rect 21652 10062 21680 10095
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 20994 9480 21050 9489
rect 20994 9415 21050 9424
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 22112 8634 22140 12106
rect 22202 11996 22510 12005
rect 22202 11994 22208 11996
rect 22264 11994 22288 11996
rect 22344 11994 22368 11996
rect 22424 11994 22448 11996
rect 22504 11994 22510 11996
rect 22264 11942 22266 11994
rect 22446 11942 22448 11994
rect 22202 11940 22208 11942
rect 22264 11940 22288 11942
rect 22344 11940 22368 11942
rect 22424 11940 22448 11942
rect 22504 11940 22510 11942
rect 22202 11931 22510 11940
rect 22202 10908 22510 10917
rect 22202 10906 22208 10908
rect 22264 10906 22288 10908
rect 22344 10906 22368 10908
rect 22424 10906 22448 10908
rect 22504 10906 22510 10908
rect 22264 10854 22266 10906
rect 22446 10854 22448 10906
rect 22202 10852 22208 10854
rect 22264 10852 22288 10854
rect 22344 10852 22368 10854
rect 22424 10852 22448 10854
rect 22504 10852 22510 10854
rect 22202 10843 22510 10852
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22296 10266 22324 10610
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22296 10010 22324 10202
rect 22204 9994 22324 10010
rect 22192 9988 22324 9994
rect 22244 9982 22324 9988
rect 22192 9930 22244 9936
rect 22202 9820 22510 9829
rect 22202 9818 22208 9820
rect 22264 9818 22288 9820
rect 22344 9818 22368 9820
rect 22424 9818 22448 9820
rect 22504 9818 22510 9820
rect 22264 9766 22266 9818
rect 22446 9766 22448 9818
rect 22202 9764 22208 9766
rect 22264 9764 22288 9766
rect 22344 9764 22368 9766
rect 22424 9764 22448 9766
rect 22504 9764 22510 9766
rect 22202 9755 22510 9764
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22480 9586 22508 9658
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22202 8732 22510 8741
rect 22202 8730 22208 8732
rect 22264 8730 22288 8732
rect 22344 8730 22368 8732
rect 22424 8730 22448 8732
rect 22504 8730 22510 8732
rect 22264 8678 22266 8730
rect 22446 8678 22448 8730
rect 22202 8676 22208 8678
rect 22264 8676 22288 8678
rect 22344 8676 22368 8678
rect 22424 8676 22448 8678
rect 22504 8676 22510 8678
rect 22202 8667 22510 8676
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21008 8090 21036 8434
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21914 7848 21970 7857
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 20824 7364 20944 7392
rect 20812 7268 20864 7274
rect 20812 7210 20864 7216
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20732 6390 20760 6802
rect 20824 6662 20852 7210
rect 20916 6798 20944 7364
rect 21192 7206 21220 7686
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21192 7002 21220 7142
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 21284 6730 21312 7822
rect 21914 7783 21916 7792
rect 21968 7783 21970 7792
rect 21916 7754 21968 7760
rect 21928 7546 21956 7754
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 22112 7478 22140 8434
rect 22388 7834 22416 8570
rect 22572 8430 22600 10406
rect 22664 8566 22692 16934
rect 22756 15994 22784 17190
rect 22848 16130 22876 19654
rect 22940 17954 22968 22596
rect 23032 19922 23060 24840
rect 23400 24818 23428 25162
rect 23388 24812 23440 24818
rect 23308 24772 23388 24800
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23216 23866 23244 24142
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23112 22704 23164 22710
rect 23112 22646 23164 22652
rect 23124 21622 23152 22646
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 23112 21480 23164 21486
rect 23112 21422 23164 21428
rect 23124 20330 23152 21422
rect 23112 20324 23164 20330
rect 23112 20266 23164 20272
rect 23020 19916 23072 19922
rect 23020 19858 23072 19864
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 23124 19378 23152 19790
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 23124 18358 23152 19110
rect 23216 18766 23244 19314
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 23112 18352 23164 18358
rect 23112 18294 23164 18300
rect 22940 17926 23060 17954
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 22940 16726 22968 16934
rect 22928 16720 22980 16726
rect 22928 16662 22980 16668
rect 22940 16250 22968 16662
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 22848 16102 22968 16130
rect 23032 16114 23060 17926
rect 23216 17202 23244 18702
rect 23204 17196 23256 17202
rect 23124 17156 23204 17184
rect 22756 15966 22876 15994
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22756 13462 22784 14486
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22744 12912 22796 12918
rect 22744 12854 22796 12860
rect 22756 10674 22784 12854
rect 22848 12170 22876 15966
rect 22836 12164 22888 12170
rect 22836 12106 22888 12112
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22744 10668 22796 10674
rect 22744 10610 22796 10616
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22756 10130 22784 10406
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22744 9988 22796 9994
rect 22744 9930 22796 9936
rect 22756 9382 22784 9930
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22652 8560 22704 8566
rect 22652 8502 22704 8508
rect 22560 8424 22612 8430
rect 22848 8378 22876 11834
rect 22940 10010 22968 16102
rect 23020 16108 23072 16114
rect 23020 16050 23072 16056
rect 23032 15706 23060 16050
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23020 13728 23072 13734
rect 23020 13670 23072 13676
rect 23032 13326 23060 13670
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 23032 12986 23060 13126
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 23032 10742 23060 11698
rect 23020 10736 23072 10742
rect 23020 10678 23072 10684
rect 23124 10130 23152 17156
rect 23204 17138 23256 17144
rect 23204 13184 23256 13190
rect 23204 13126 23256 13132
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 22940 9982 23060 10010
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22940 9722 22968 9862
rect 22928 9716 22980 9722
rect 22928 9658 22980 9664
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 22560 8366 22612 8372
rect 22756 8350 22876 8378
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22480 8090 22508 8230
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22652 7880 22704 7886
rect 22388 7806 22600 7834
rect 22652 7822 22704 7828
rect 22202 7644 22510 7653
rect 22202 7642 22208 7644
rect 22264 7642 22288 7644
rect 22344 7642 22368 7644
rect 22424 7642 22448 7644
rect 22504 7642 22510 7644
rect 22264 7590 22266 7642
rect 22446 7590 22448 7642
rect 22202 7588 22208 7590
rect 22264 7588 22288 7590
rect 22344 7588 22368 7590
rect 22424 7588 22448 7590
rect 22504 7588 22510 7590
rect 22202 7579 22510 7588
rect 22100 7472 22152 7478
rect 22100 7414 22152 7420
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 21272 6724 21324 6730
rect 21272 6666 21324 6672
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20732 4282 20760 4422
rect 20720 4276 20772 4282
rect 20720 4218 20772 4224
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20548 3058 20576 3334
rect 20732 3058 20760 4218
rect 20824 4078 20852 6190
rect 21100 6118 21128 6598
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20824 3738 20852 4014
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20916 3534 20944 4082
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 21008 3534 21036 3946
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 19904 2746 20208 2774
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 1952 2372 2004 2378
rect 1952 2314 2004 2320
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 1490 2136 1546 2145
rect 1490 2071 1546 2080
rect 1964 800 1992 2314
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 3896 800 3924 2246
rect 5828 800 5856 2246
rect 8034 2204 8342 2213
rect 8034 2202 8040 2204
rect 8096 2202 8120 2204
rect 8176 2202 8200 2204
rect 8256 2202 8280 2204
rect 8336 2202 8342 2204
rect 8096 2150 8098 2202
rect 8278 2150 8280 2202
rect 8034 2148 8040 2150
rect 8096 2148 8120 2150
rect 8176 2148 8200 2150
rect 8256 2148 8280 2150
rect 8336 2148 8342 2150
rect 8034 2139 8342 2148
rect 8404 800 8432 2246
rect 10336 800 10364 2246
rect 12268 800 12296 2314
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14844 800 14872 2246
rect 15118 2204 15426 2213
rect 15118 2202 15124 2204
rect 15180 2202 15204 2204
rect 15260 2202 15284 2204
rect 15340 2202 15364 2204
rect 15420 2202 15426 2204
rect 15180 2150 15182 2202
rect 15362 2150 15364 2202
rect 15118 2148 15124 2150
rect 15180 2148 15204 2150
rect 15260 2148 15284 2150
rect 15340 2148 15364 2150
rect 15420 2148 15426 2150
rect 15118 2139 15426 2148
rect 16776 800 16804 2314
rect 18708 800 18736 2382
rect 19904 2378 19932 2746
rect 20916 2650 20944 3470
rect 20996 3120 21048 3126
rect 21100 3108 21128 6054
rect 21192 5642 21220 6054
rect 21284 5914 21312 6666
rect 21376 6254 21404 6666
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21180 5636 21232 5642
rect 21180 5578 21232 5584
rect 21836 5234 21864 7142
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 22020 6458 22048 6734
rect 22202 6556 22510 6565
rect 22202 6554 22208 6556
rect 22264 6554 22288 6556
rect 22344 6554 22368 6556
rect 22424 6554 22448 6556
rect 22504 6554 22510 6556
rect 22264 6502 22266 6554
rect 22446 6502 22448 6554
rect 22202 6500 22208 6502
rect 22264 6500 22288 6502
rect 22344 6500 22368 6502
rect 22424 6500 22448 6502
rect 22504 6500 22510 6502
rect 22202 6491 22510 6500
rect 22008 6452 22060 6458
rect 22008 6394 22060 6400
rect 21916 5840 21968 5846
rect 21916 5782 21968 5788
rect 21928 5234 21956 5782
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 22020 4758 22048 6394
rect 22468 6180 22520 6186
rect 22468 6122 22520 6128
rect 22480 5574 22508 6122
rect 22572 5914 22600 7806
rect 22664 7342 22692 7822
rect 22756 7750 22784 8350
rect 22836 8288 22888 8294
rect 22836 8230 22888 8236
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22848 7410 22876 8230
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 22744 6792 22796 6798
rect 22796 6752 22876 6780
rect 22744 6734 22796 6740
rect 22744 6656 22796 6662
rect 22744 6598 22796 6604
rect 22756 6322 22784 6598
rect 22848 6390 22876 6752
rect 22836 6384 22888 6390
rect 22836 6326 22888 6332
rect 22744 6316 22796 6322
rect 22744 6258 22796 6264
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 22202 5468 22510 5477
rect 22202 5466 22208 5468
rect 22264 5466 22288 5468
rect 22344 5466 22368 5468
rect 22424 5466 22448 5468
rect 22504 5466 22510 5468
rect 22264 5414 22266 5466
rect 22446 5414 22448 5466
rect 22202 5412 22208 5414
rect 22264 5412 22288 5414
rect 22344 5412 22368 5414
rect 22424 5412 22448 5414
rect 22504 5412 22510 5414
rect 22202 5403 22510 5412
rect 22572 5370 22600 5850
rect 22560 5364 22612 5370
rect 22560 5306 22612 5312
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 22008 4752 22060 4758
rect 22008 4694 22060 4700
rect 22204 4570 22232 5238
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22468 5092 22520 5098
rect 22468 5034 22520 5040
rect 22480 4622 22508 5034
rect 22112 4542 22232 4570
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 21468 3534 21496 4014
rect 21836 3602 21864 4082
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21928 3534 21956 4082
rect 22112 3738 22140 4542
rect 22202 4380 22510 4389
rect 22202 4378 22208 4380
rect 22264 4378 22288 4380
rect 22344 4378 22368 4380
rect 22424 4378 22448 4380
rect 22504 4378 22510 4380
rect 22264 4326 22266 4378
rect 22446 4326 22448 4378
rect 22202 4324 22208 4326
rect 22264 4324 22288 4326
rect 22344 4324 22368 4326
rect 22424 4324 22448 4326
rect 22504 4324 22510 4326
rect 22202 4315 22510 4324
rect 22572 4282 22600 5170
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 22756 4010 22784 6258
rect 22848 5778 22876 6326
rect 22940 6186 22968 9318
rect 23032 8634 23060 9982
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 23216 7342 23244 13126
rect 23308 11898 23336 24772
rect 23388 24754 23440 24760
rect 23584 24274 23612 25978
rect 23768 24410 23796 28358
rect 23940 27940 23992 27946
rect 23940 27882 23992 27888
rect 23952 27062 23980 27882
rect 24308 27872 24360 27878
rect 24308 27814 24360 27820
rect 24320 27470 24348 27814
rect 24308 27464 24360 27470
rect 24308 27406 24360 27412
rect 23940 27056 23992 27062
rect 23940 26998 23992 27004
rect 23756 24404 23808 24410
rect 23756 24346 23808 24352
rect 23572 24268 23624 24274
rect 23572 24210 23624 24216
rect 23952 23662 23980 26998
rect 24320 26926 24348 27406
rect 24308 26920 24360 26926
rect 24308 26862 24360 26868
rect 24320 26790 24348 26862
rect 24308 26784 24360 26790
rect 24308 26726 24360 26732
rect 24216 24608 24268 24614
rect 24216 24550 24268 24556
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 24228 23118 24256 24550
rect 24216 23112 24268 23118
rect 24216 23054 24268 23060
rect 24228 22710 24256 23054
rect 24216 22704 24268 22710
rect 24216 22646 24268 22652
rect 24032 22500 24084 22506
rect 24032 22442 24084 22448
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23400 20942 23428 22374
rect 24044 21690 24072 22442
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 24136 21554 24164 21830
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23492 20534 23520 20742
rect 23480 20528 23532 20534
rect 23480 20470 23532 20476
rect 23492 19446 23520 20470
rect 23480 19440 23532 19446
rect 23480 19382 23532 19388
rect 23492 18834 23520 19382
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23388 17876 23440 17882
rect 23388 17818 23440 17824
rect 23400 17338 23428 17818
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23400 16590 23428 17274
rect 23584 17134 23612 21286
rect 23676 20942 23704 21422
rect 24044 21418 24072 21490
rect 24032 21412 24084 21418
rect 24032 21354 24084 21360
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23848 20800 23900 20806
rect 23848 20742 23900 20748
rect 23860 20466 23888 20742
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 23584 16590 23612 17070
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23400 15706 23428 16526
rect 23676 16250 23704 18906
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 23768 17270 23796 18158
rect 23756 17264 23808 17270
rect 23756 17206 23808 17212
rect 23768 16658 23796 17206
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23676 16046 23704 16186
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 23308 10674 23336 11630
rect 23400 11286 23428 15506
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23584 14074 23612 14758
rect 23572 14068 23624 14074
rect 23572 14010 23624 14016
rect 23480 13252 23532 13258
rect 23480 13194 23532 13200
rect 23492 12918 23520 13194
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23584 12850 23612 14010
rect 23664 12912 23716 12918
rect 23664 12854 23716 12860
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23492 11898 23520 12718
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23676 11762 23704 12854
rect 23860 12434 23888 20402
rect 24228 17218 24256 22646
rect 24136 17190 24256 17218
rect 24030 16552 24086 16561
rect 24030 16487 24086 16496
rect 24044 16250 24072 16487
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23952 15366 23980 15506
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23952 14618 23980 15302
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 23952 14414 23980 14554
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23952 13462 23980 14350
rect 24044 14006 24072 16186
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 23940 13456 23992 13462
rect 23940 13398 23992 13404
rect 23768 12406 23888 12434
rect 23768 11830 23796 12406
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23768 11354 23796 11766
rect 24044 11762 24072 12038
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 24032 11756 24084 11762
rect 24032 11698 24084 11704
rect 23756 11348 23808 11354
rect 23756 11290 23808 11296
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23400 10810 23428 11222
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23860 10674 23888 11698
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23952 11257 23980 11494
rect 23938 11248 23994 11257
rect 23938 11183 23994 11192
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23296 10532 23348 10538
rect 23296 10474 23348 10480
rect 23308 9994 23336 10474
rect 23400 10266 23428 10610
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23662 10024 23718 10033
rect 23296 9988 23348 9994
rect 23662 9959 23718 9968
rect 23296 9930 23348 9936
rect 23308 9654 23336 9930
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 23308 9178 23336 9590
rect 23480 9512 23532 9518
rect 23478 9480 23480 9489
rect 23532 9480 23534 9489
rect 23478 9415 23534 9424
rect 23676 9382 23704 9959
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23296 9172 23348 9178
rect 23296 9114 23348 9120
rect 23676 8634 23704 9318
rect 23860 9042 23888 9522
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23860 8838 23888 8978
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23676 7954 23704 8570
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23584 7002 23612 7346
rect 23572 6996 23624 7002
rect 23572 6938 23624 6944
rect 23676 6730 23704 7890
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23664 6724 23716 6730
rect 23664 6666 23716 6672
rect 23676 6390 23704 6666
rect 23664 6384 23716 6390
rect 23664 6326 23716 6332
rect 22928 6180 22980 6186
rect 22928 6122 22980 6128
rect 22836 5772 22888 5778
rect 22836 5714 22888 5720
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 23032 4010 23060 5306
rect 23768 5234 23796 7686
rect 23860 6730 23888 7822
rect 23848 6724 23900 6730
rect 23848 6666 23900 6672
rect 23860 6458 23888 6666
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 22744 4004 22796 4010
rect 22744 3946 22796 3952
rect 23020 4004 23072 4010
rect 23020 3946 23072 3952
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 22756 3534 22784 3946
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 21468 3194 21496 3470
rect 22202 3292 22510 3301
rect 22202 3290 22208 3292
rect 22264 3290 22288 3292
rect 22344 3290 22368 3292
rect 22424 3290 22448 3292
rect 22504 3290 22510 3292
rect 22264 3238 22266 3290
rect 22446 3238 22448 3290
rect 22202 3236 22208 3238
rect 22264 3236 22288 3238
rect 22344 3236 22368 3238
rect 22424 3236 22448 3238
rect 22504 3236 22510 3238
rect 22202 3227 22510 3236
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21048 3080 21128 3108
rect 20996 3062 21048 3068
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 21008 2446 21036 3062
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21836 2446 21864 2926
rect 22940 2582 22968 3878
rect 23032 3466 23060 3946
rect 23124 3670 23152 4966
rect 23400 4826 23428 5170
rect 23478 5128 23534 5137
rect 23478 5063 23480 5072
rect 23532 5063 23534 5072
rect 23480 5034 23532 5040
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23216 4146 23244 4422
rect 23492 4185 23520 5034
rect 23664 4752 23716 4758
rect 23664 4694 23716 4700
rect 23478 4176 23534 4185
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23296 4140 23348 4146
rect 23478 4111 23534 4120
rect 23296 4082 23348 4088
rect 23308 3738 23336 4082
rect 23492 3942 23520 4111
rect 23676 4078 23704 4694
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23112 3664 23164 3670
rect 23112 3606 23164 3612
rect 23492 3602 23520 3878
rect 23676 3738 23704 4014
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 23860 3534 23888 4082
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 23032 3194 23060 3402
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 24136 2774 24164 17190
rect 24308 17060 24360 17066
rect 24308 17002 24360 17008
rect 24320 16114 24348 17002
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24320 15026 24348 16050
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24308 14884 24360 14890
rect 24308 14826 24360 14832
rect 24320 14618 24348 14826
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24308 14340 24360 14346
rect 24308 14282 24360 14288
rect 24320 14074 24348 14282
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24228 13530 24256 13670
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24320 13326 24348 14010
rect 24308 13320 24360 13326
rect 24308 13262 24360 13268
rect 24412 10713 24440 29990
rect 24504 29850 24532 30194
rect 26344 30054 26372 30194
rect 26436 30122 26464 31965
rect 27620 30252 27672 30258
rect 27620 30194 27672 30200
rect 28264 30252 28316 30258
rect 28264 30194 28316 30200
rect 26424 30116 26476 30122
rect 26424 30058 26476 30064
rect 26332 30048 26384 30054
rect 26332 29990 26384 29996
rect 25744 29948 26052 29957
rect 25744 29946 25750 29948
rect 25806 29946 25830 29948
rect 25886 29946 25910 29948
rect 25966 29946 25990 29948
rect 26046 29946 26052 29948
rect 25806 29894 25808 29946
rect 25988 29894 25990 29946
rect 25744 29892 25750 29894
rect 25806 29892 25830 29894
rect 25886 29892 25910 29894
rect 25966 29892 25990 29894
rect 26046 29892 26052 29894
rect 25744 29883 26052 29892
rect 24492 29844 24544 29850
rect 24492 29786 24544 29792
rect 25744 28860 26052 28869
rect 25744 28858 25750 28860
rect 25806 28858 25830 28860
rect 25886 28858 25910 28860
rect 25966 28858 25990 28860
rect 26046 28858 26052 28860
rect 25806 28806 25808 28858
rect 25988 28806 25990 28858
rect 25744 28804 25750 28806
rect 25806 28804 25830 28806
rect 25886 28804 25910 28806
rect 25966 28804 25990 28806
rect 26046 28804 26052 28806
rect 25744 28795 26052 28804
rect 26344 28665 26372 29990
rect 27632 29510 27660 30194
rect 27896 30048 27948 30054
rect 27894 30016 27896 30025
rect 27948 30016 27950 30025
rect 27894 29951 27950 29960
rect 27620 29504 27672 29510
rect 27620 29446 27672 29452
rect 27632 29345 27660 29446
rect 27618 29336 27674 29345
rect 27618 29271 27674 29280
rect 28276 29034 28304 30194
rect 28368 30122 28396 31965
rect 29286 30492 29594 30501
rect 29286 30490 29292 30492
rect 29348 30490 29372 30492
rect 29428 30490 29452 30492
rect 29508 30490 29532 30492
rect 29588 30490 29594 30492
rect 29348 30438 29350 30490
rect 29530 30438 29532 30490
rect 29286 30436 29292 30438
rect 29348 30436 29372 30438
rect 29428 30436 29452 30438
rect 29508 30436 29532 30438
rect 29588 30436 29594 30438
rect 29286 30427 29594 30436
rect 28356 30116 28408 30122
rect 28356 30058 28408 30064
rect 30300 29646 30328 31965
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 28816 29504 28868 29510
rect 28816 29446 28868 29452
rect 28264 29028 28316 29034
rect 28264 28970 28316 28976
rect 26330 28656 26386 28665
rect 26330 28591 26386 28600
rect 28276 28529 28304 28970
rect 28262 28520 28318 28529
rect 28262 28455 28318 28464
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24504 28014 24532 28358
rect 24676 28212 24728 28218
rect 24676 28154 24728 28160
rect 24584 28144 24636 28150
rect 24584 28086 24636 28092
rect 24492 28008 24544 28014
rect 24492 27950 24544 27956
rect 24596 27470 24624 28086
rect 24688 27538 24716 28154
rect 28632 28076 28684 28082
rect 28632 28018 28684 28024
rect 28644 27985 28672 28018
rect 25502 27976 25558 27985
rect 28630 27976 28686 27985
rect 25502 27911 25558 27920
rect 26148 27940 26200 27946
rect 25516 27674 25544 27911
rect 28630 27911 28686 27920
rect 26148 27882 26200 27888
rect 25744 27772 26052 27781
rect 25744 27770 25750 27772
rect 25806 27770 25830 27772
rect 25886 27770 25910 27772
rect 25966 27770 25990 27772
rect 26046 27770 26052 27772
rect 25806 27718 25808 27770
rect 25988 27718 25990 27770
rect 25744 27716 25750 27718
rect 25806 27716 25830 27718
rect 25886 27716 25910 27718
rect 25966 27716 25990 27718
rect 26046 27716 26052 27718
rect 25744 27707 26052 27716
rect 25504 27668 25556 27674
rect 25504 27610 25556 27616
rect 24676 27532 24728 27538
rect 24676 27474 24728 27480
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24596 26926 24624 27406
rect 24688 27130 24716 27474
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 25596 27464 25648 27470
rect 25596 27406 25648 27412
rect 25148 27130 25176 27406
rect 24676 27124 24728 27130
rect 24676 27066 24728 27072
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 25044 27056 25096 27062
rect 25044 26998 25096 27004
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24584 26920 24636 26926
rect 24584 26862 24636 26868
rect 24492 26376 24544 26382
rect 24596 26364 24624 26862
rect 24872 26450 24900 26930
rect 24860 26444 24912 26450
rect 24860 26386 24912 26392
rect 24544 26336 24624 26364
rect 24492 26318 24544 26324
rect 24596 25294 24624 26336
rect 24952 25968 25004 25974
rect 25056 25956 25084 26998
rect 25148 26790 25176 27066
rect 25136 26784 25188 26790
rect 25136 26726 25188 26732
rect 25004 25928 25084 25956
rect 24952 25910 25004 25916
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24596 24138 24624 25230
rect 24964 24818 24992 25910
rect 25044 25424 25096 25430
rect 25044 25366 25096 25372
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24964 24274 24992 24754
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24584 24132 24636 24138
rect 24584 24074 24636 24080
rect 24860 24132 24912 24138
rect 24860 24074 24912 24080
rect 24872 23662 24900 24074
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24780 22778 24808 23054
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24780 22545 24808 22714
rect 24766 22536 24822 22545
rect 24766 22471 24822 22480
rect 24768 21956 24820 21962
rect 24768 21898 24820 21904
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24596 21010 24624 21830
rect 24780 21554 24808 21898
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 24492 20868 24544 20874
rect 24492 20810 24544 20816
rect 24504 20466 24532 20810
rect 24492 20460 24544 20466
rect 24492 20402 24544 20408
rect 24596 19378 24624 20946
rect 24780 20806 24808 21490
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 25056 20602 25084 25366
rect 25148 25294 25176 26726
rect 25608 26246 25636 27406
rect 26160 26994 26188 27882
rect 26148 26988 26200 26994
rect 26148 26930 26200 26936
rect 25744 26684 26052 26693
rect 25744 26682 25750 26684
rect 25806 26682 25830 26684
rect 25886 26682 25910 26684
rect 25966 26682 25990 26684
rect 26046 26682 26052 26684
rect 25806 26630 25808 26682
rect 25988 26630 25990 26682
rect 25744 26628 25750 26630
rect 25806 26628 25830 26630
rect 25886 26628 25910 26630
rect 25966 26628 25990 26630
rect 26046 26628 26052 26630
rect 25744 26619 26052 26628
rect 26160 26450 26188 26930
rect 28632 26784 28684 26790
rect 28632 26726 28684 26732
rect 26148 26444 26200 26450
rect 26148 26386 26200 26392
rect 25964 26376 26016 26382
rect 25964 26318 26016 26324
rect 25596 26240 25648 26246
rect 25596 26182 25648 26188
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 25148 24138 25176 25230
rect 25608 25226 25636 26182
rect 25976 25974 26004 26318
rect 26160 26042 26188 26386
rect 28644 26314 28672 26726
rect 28356 26308 28408 26314
rect 28356 26250 28408 26256
rect 28632 26308 28684 26314
rect 28632 26250 28684 26256
rect 26148 26036 26200 26042
rect 26200 25996 26280 26024
rect 26148 25978 26200 25984
rect 25964 25968 26016 25974
rect 25964 25910 26016 25916
rect 26148 25696 26200 25702
rect 26148 25638 26200 25644
rect 25744 25596 26052 25605
rect 25744 25594 25750 25596
rect 25806 25594 25830 25596
rect 25886 25594 25910 25596
rect 25966 25594 25990 25596
rect 26046 25594 26052 25596
rect 25806 25542 25808 25594
rect 25988 25542 25990 25594
rect 25744 25540 25750 25542
rect 25806 25540 25830 25542
rect 25886 25540 25910 25542
rect 25966 25540 25990 25542
rect 26046 25540 26052 25542
rect 25744 25531 26052 25540
rect 26160 25362 26188 25638
rect 26148 25356 26200 25362
rect 26148 25298 26200 25304
rect 26252 25294 26280 25996
rect 26884 25968 26936 25974
rect 26884 25910 26936 25916
rect 26896 25498 26924 25910
rect 27712 25764 27764 25770
rect 27712 25706 27764 25712
rect 27620 25696 27672 25702
rect 27620 25638 27672 25644
rect 27632 25498 27660 25638
rect 26884 25492 26936 25498
rect 26884 25434 26936 25440
rect 27620 25492 27672 25498
rect 27620 25434 27672 25440
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 26240 25288 26292 25294
rect 26240 25230 26292 25236
rect 25596 25220 25648 25226
rect 25596 25162 25648 25168
rect 25700 24954 25728 25230
rect 25688 24948 25740 24954
rect 25688 24890 25740 24896
rect 25688 24812 25740 24818
rect 25516 24772 25688 24800
rect 25320 24744 25372 24750
rect 25240 24704 25320 24732
rect 25240 24274 25268 24704
rect 25320 24686 25372 24692
rect 25412 24336 25464 24342
rect 25412 24278 25464 24284
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25136 24132 25188 24138
rect 25136 24074 25188 24080
rect 25148 23526 25176 24074
rect 25240 23866 25268 24210
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25240 23186 25268 23802
rect 25332 23730 25360 24142
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25228 23180 25280 23186
rect 25148 23140 25228 23168
rect 25148 22642 25176 23140
rect 25228 23122 25280 23128
rect 25332 23118 25360 23666
rect 25320 23112 25372 23118
rect 25320 23054 25372 23060
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 25332 22574 25360 23054
rect 25320 22568 25372 22574
rect 25320 22510 25372 22516
rect 25044 20596 25096 20602
rect 25044 20538 25096 20544
rect 24768 20392 24820 20398
rect 24768 20334 24820 20340
rect 24780 19786 24808 20334
rect 24768 19780 24820 19786
rect 24768 19722 24820 19728
rect 24584 19372 24636 19378
rect 24636 19320 24716 19334
rect 24584 19314 24716 19320
rect 24596 19306 24716 19314
rect 24780 19310 24808 19722
rect 24688 18970 24716 19306
rect 24768 19304 24820 19310
rect 24768 19246 24820 19252
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24492 17536 24544 17542
rect 24492 17478 24544 17484
rect 24504 14006 24532 17478
rect 24596 15638 24624 17614
rect 24584 15632 24636 15638
rect 24584 15574 24636 15580
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24596 14414 24624 15302
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24492 14000 24544 14006
rect 24492 13942 24544 13948
rect 24688 13938 24716 18566
rect 24964 18358 24992 18566
rect 24952 18352 25004 18358
rect 24952 18294 25004 18300
rect 24964 17678 24992 18294
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24780 16182 24808 16390
rect 25056 16250 25084 20538
rect 25332 16590 25360 22510
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 24768 16176 24820 16182
rect 24768 16118 24820 16124
rect 24780 15162 24808 16118
rect 25056 15502 25084 16186
rect 25424 15994 25452 24278
rect 25516 23662 25544 24772
rect 25688 24754 25740 24760
rect 25596 24608 25648 24614
rect 25596 24550 25648 24556
rect 25608 24206 25636 24550
rect 25744 24508 26052 24517
rect 25744 24506 25750 24508
rect 25806 24506 25830 24508
rect 25886 24506 25910 24508
rect 25966 24506 25990 24508
rect 26046 24506 26052 24508
rect 25806 24454 25808 24506
rect 25988 24454 25990 24506
rect 25744 24452 25750 24454
rect 25806 24452 25830 24454
rect 25886 24452 25910 24454
rect 25966 24452 25990 24454
rect 26046 24452 26052 24454
rect 25744 24443 26052 24452
rect 26252 24274 26280 25230
rect 26976 24608 27028 24614
rect 26976 24550 27028 24556
rect 26240 24268 26292 24274
rect 26240 24210 26292 24216
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 26160 23730 26188 24142
rect 26148 23724 26200 23730
rect 26148 23666 26200 23672
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25744 23420 26052 23429
rect 25744 23418 25750 23420
rect 25806 23418 25830 23420
rect 25886 23418 25910 23420
rect 25966 23418 25990 23420
rect 26046 23418 26052 23420
rect 25806 23366 25808 23418
rect 25988 23366 25990 23418
rect 25744 23364 25750 23366
rect 25806 23364 25830 23366
rect 25886 23364 25910 23366
rect 25966 23364 25990 23366
rect 26046 23364 26052 23366
rect 25744 23355 26052 23364
rect 25964 22976 26016 22982
rect 26160 22964 26188 23666
rect 26884 23588 26936 23594
rect 26884 23530 26936 23536
rect 26238 23216 26294 23225
rect 26238 23151 26240 23160
rect 26292 23151 26294 23160
rect 26240 23122 26292 23128
rect 26016 22936 26188 22964
rect 25964 22918 26016 22924
rect 25976 22778 26004 22918
rect 25964 22772 26016 22778
rect 25964 22714 26016 22720
rect 25596 22432 25648 22438
rect 25596 22374 25648 22380
rect 25608 22030 25636 22374
rect 25744 22332 26052 22341
rect 25744 22330 25750 22332
rect 25806 22330 25830 22332
rect 25886 22330 25910 22332
rect 25966 22330 25990 22332
rect 26046 22330 26052 22332
rect 25806 22278 25808 22330
rect 25988 22278 25990 22330
rect 25744 22276 25750 22278
rect 25806 22276 25830 22278
rect 25886 22276 25910 22278
rect 25966 22276 25990 22278
rect 26046 22276 26052 22278
rect 25744 22267 26052 22276
rect 26792 22094 26844 22098
rect 26896 22094 26924 23530
rect 26988 23186 27016 24550
rect 27528 23520 27580 23526
rect 27528 23462 27580 23468
rect 26976 23180 27028 23186
rect 26976 23122 27028 23128
rect 26792 22092 26924 22094
rect 26844 22066 26924 22092
rect 26792 22034 26844 22040
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 26896 21486 26924 22066
rect 26988 21894 27016 23122
rect 26976 21888 27028 21894
rect 26976 21830 27028 21836
rect 27252 21888 27304 21894
rect 27252 21830 27304 21836
rect 26424 21480 26476 21486
rect 26424 21422 26476 21428
rect 26884 21480 26936 21486
rect 26884 21422 26936 21428
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 25744 21244 26052 21253
rect 25744 21242 25750 21244
rect 25806 21242 25830 21244
rect 25886 21242 25910 21244
rect 25966 21242 25990 21244
rect 26046 21242 26052 21244
rect 25806 21190 25808 21242
rect 25988 21190 25990 21242
rect 25744 21188 25750 21190
rect 25806 21188 25830 21190
rect 25886 21188 25910 21190
rect 25966 21188 25990 21190
rect 26046 21188 26052 21190
rect 25744 21179 26052 21188
rect 26252 21146 26280 21286
rect 26056 21140 26108 21146
rect 26056 21082 26108 21088
rect 26240 21140 26292 21146
rect 26240 21082 26292 21088
rect 26068 21026 26096 21082
rect 26068 20998 26372 21026
rect 26436 21010 26464 21422
rect 26516 21412 26568 21418
rect 26516 21354 26568 21360
rect 26148 20800 26200 20806
rect 26148 20742 26200 20748
rect 25596 20528 25648 20534
rect 25596 20470 25648 20476
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25516 19990 25544 20198
rect 25608 20058 25636 20470
rect 26160 20466 26188 20742
rect 26148 20460 26200 20466
rect 26148 20402 26200 20408
rect 25744 20156 26052 20165
rect 25744 20154 25750 20156
rect 25806 20154 25830 20156
rect 25886 20154 25910 20156
rect 25966 20154 25990 20156
rect 26046 20154 26052 20156
rect 25806 20102 25808 20154
rect 25988 20102 25990 20154
rect 25744 20100 25750 20102
rect 25806 20100 25830 20102
rect 25886 20100 25910 20102
rect 25966 20100 25990 20102
rect 26046 20100 26052 20102
rect 25744 20091 26052 20100
rect 25596 20052 25648 20058
rect 25596 19994 25648 20000
rect 25504 19984 25556 19990
rect 25504 19926 25556 19932
rect 25744 19068 26052 19077
rect 25744 19066 25750 19068
rect 25806 19066 25830 19068
rect 25886 19066 25910 19068
rect 25966 19066 25990 19068
rect 26046 19066 26052 19068
rect 25806 19014 25808 19066
rect 25988 19014 25990 19066
rect 25744 19012 25750 19014
rect 25806 19012 25830 19014
rect 25886 19012 25910 19014
rect 25966 19012 25990 19014
rect 26046 19012 26052 19014
rect 25744 19003 26052 19012
rect 26160 18766 26188 20402
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 26252 20058 26280 20334
rect 26240 20052 26292 20058
rect 26240 19994 26292 20000
rect 26252 18834 26280 19994
rect 26344 19310 26372 20998
rect 26424 21004 26476 21010
rect 26424 20946 26476 20952
rect 26528 20942 26556 21354
rect 26700 21004 26752 21010
rect 26700 20946 26752 20952
rect 26516 20936 26568 20942
rect 26516 20878 26568 20884
rect 26332 19304 26384 19310
rect 26332 19246 26384 19252
rect 26240 18828 26292 18834
rect 26240 18770 26292 18776
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 25744 17980 26052 17989
rect 25744 17978 25750 17980
rect 25806 17978 25830 17980
rect 25886 17978 25910 17980
rect 25966 17978 25990 17980
rect 26046 17978 26052 17980
rect 25806 17926 25808 17978
rect 25988 17926 25990 17978
rect 25744 17924 25750 17926
rect 25806 17924 25830 17926
rect 25886 17924 25910 17926
rect 25966 17924 25990 17926
rect 26046 17924 26052 17926
rect 25744 17915 26052 17924
rect 25744 16892 26052 16901
rect 25744 16890 25750 16892
rect 25806 16890 25830 16892
rect 25886 16890 25910 16892
rect 25966 16890 25990 16892
rect 26046 16890 26052 16892
rect 25806 16838 25808 16890
rect 25988 16838 25990 16890
rect 25744 16836 25750 16838
rect 25806 16836 25830 16838
rect 25886 16836 25910 16838
rect 25966 16836 25990 16838
rect 26046 16836 26052 16838
rect 25744 16827 26052 16836
rect 26252 16658 26280 18770
rect 26528 18358 26556 20878
rect 26516 18352 26568 18358
rect 26516 18294 26568 18300
rect 26712 18222 26740 20946
rect 26700 18216 26752 18222
rect 26700 18158 26752 18164
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26344 17134 26372 17478
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 25332 15966 25452 15994
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 24860 15360 24912 15366
rect 24860 15302 24912 15308
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24780 14074 24808 14418
rect 24872 14414 24900 15302
rect 25228 14884 25280 14890
rect 25228 14826 25280 14832
rect 25042 14512 25098 14521
rect 25042 14447 25044 14456
rect 25096 14447 25098 14456
rect 25044 14418 25096 14424
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24584 13796 24636 13802
rect 24584 13738 24636 13744
rect 24596 13190 24624 13738
rect 24768 13456 24820 13462
rect 24768 13398 24820 13404
rect 24584 13184 24636 13190
rect 24584 13126 24636 13132
rect 24596 12646 24624 13126
rect 24780 12986 24808 13398
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24596 11830 24624 12582
rect 24676 12164 24728 12170
rect 24676 12106 24728 12112
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24688 11762 24716 12106
rect 24780 11762 24808 12922
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 24780 11354 24808 11698
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24398 10704 24454 10713
rect 24872 10674 24900 12242
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24398 10639 24454 10648
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24214 10568 24270 10577
rect 24214 10503 24216 10512
rect 24268 10503 24270 10512
rect 24860 10532 24912 10538
rect 24216 10474 24268 10480
rect 24860 10474 24912 10480
rect 24872 9178 24900 10474
rect 24964 9654 24992 11698
rect 25148 10810 25176 12786
rect 25240 12238 25268 14826
rect 25332 14278 25360 15966
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 25424 15502 25452 15846
rect 25744 15804 26052 15813
rect 25744 15802 25750 15804
rect 25806 15802 25830 15804
rect 25886 15802 25910 15804
rect 25966 15802 25990 15804
rect 26046 15802 26052 15804
rect 25806 15750 25808 15802
rect 25988 15750 25990 15802
rect 25744 15748 25750 15750
rect 25806 15748 25830 15750
rect 25886 15748 25910 15750
rect 25966 15748 25990 15750
rect 26046 15748 26052 15750
rect 25744 15739 26052 15748
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25504 14952 25556 14958
rect 25504 14894 25556 14900
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 25516 13326 25544 14894
rect 25744 14716 26052 14725
rect 25744 14714 25750 14716
rect 25806 14714 25830 14716
rect 25886 14714 25910 14716
rect 25966 14714 25990 14716
rect 26046 14714 26052 14716
rect 25806 14662 25808 14714
rect 25988 14662 25990 14714
rect 25744 14660 25750 14662
rect 25806 14660 25830 14662
rect 25886 14660 25910 14662
rect 25966 14660 25990 14662
rect 26046 14660 26052 14662
rect 25744 14651 26052 14660
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 25596 14340 25648 14346
rect 25596 14282 25648 14288
rect 25608 13530 25636 14282
rect 25744 13628 26052 13637
rect 25744 13626 25750 13628
rect 25806 13626 25830 13628
rect 25886 13626 25910 13628
rect 25966 13626 25990 13628
rect 26046 13626 26052 13628
rect 25806 13574 25808 13626
rect 25988 13574 25990 13626
rect 25744 13572 25750 13574
rect 25806 13572 25830 13574
rect 25886 13572 25910 13574
rect 25966 13572 25990 13574
rect 26046 13572 26052 13574
rect 25744 13563 26052 13572
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25504 13320 25556 13326
rect 25504 13262 25556 13268
rect 25516 12306 25544 13262
rect 25744 12540 26052 12549
rect 25744 12538 25750 12540
rect 25806 12538 25830 12540
rect 25886 12538 25910 12540
rect 25966 12538 25990 12540
rect 26046 12538 26052 12540
rect 25806 12486 25808 12538
rect 25988 12486 25990 12538
rect 25744 12484 25750 12486
rect 25806 12484 25830 12486
rect 25886 12484 25910 12486
rect 25966 12484 25990 12486
rect 26046 12484 26052 12486
rect 25744 12475 26052 12484
rect 26160 12442 26188 14554
rect 26344 14346 26372 17070
rect 26424 16788 26476 16794
rect 26424 16730 26476 16736
rect 26436 16454 26464 16730
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26252 12850 26280 13262
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 26148 12436 26200 12442
rect 26148 12378 26200 12384
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 26160 12238 26188 12378
rect 25228 12232 25280 12238
rect 25228 12174 25280 12180
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26148 12096 26200 12102
rect 26148 12038 26200 12044
rect 25744 11452 26052 11461
rect 25744 11450 25750 11452
rect 25806 11450 25830 11452
rect 25886 11450 25910 11452
rect 25966 11450 25990 11452
rect 26046 11450 26052 11452
rect 25806 11398 25808 11450
rect 25988 11398 25990 11450
rect 25744 11396 25750 11398
rect 25806 11396 25830 11398
rect 25886 11396 25910 11398
rect 25966 11396 25990 11398
rect 26046 11396 26052 11398
rect 25744 11387 26052 11396
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 25148 10266 25176 10542
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 25332 10130 25360 10610
rect 25516 10169 25544 11086
rect 25688 10668 25740 10674
rect 25688 10610 25740 10616
rect 25596 10532 25648 10538
rect 25596 10474 25648 10480
rect 25502 10160 25558 10169
rect 25320 10124 25372 10130
rect 25608 10130 25636 10474
rect 25700 10470 25728 10610
rect 25688 10464 25740 10470
rect 25688 10406 25740 10412
rect 25744 10364 26052 10373
rect 25744 10362 25750 10364
rect 25806 10362 25830 10364
rect 25886 10362 25910 10364
rect 25966 10362 25990 10364
rect 26046 10362 26052 10364
rect 25806 10310 25808 10362
rect 25988 10310 25990 10362
rect 25744 10308 25750 10310
rect 25806 10308 25830 10310
rect 25886 10308 25910 10310
rect 25966 10308 25990 10310
rect 26046 10308 26052 10310
rect 25744 10299 26052 10308
rect 25502 10095 25558 10104
rect 25596 10124 25648 10130
rect 25320 10066 25372 10072
rect 25332 9874 25360 10066
rect 25516 10062 25544 10095
rect 25596 10066 25648 10072
rect 25504 10056 25556 10062
rect 25504 9998 25556 10004
rect 25240 9846 25360 9874
rect 25412 9920 25464 9926
rect 25412 9862 25464 9868
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 25136 9648 25188 9654
rect 25136 9590 25188 9596
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24216 8832 24268 8838
rect 24216 8774 24268 8780
rect 24228 6458 24256 8774
rect 25148 7546 25176 9590
rect 25240 9586 25268 9846
rect 25424 9586 25452 9862
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 25412 9580 25464 9586
rect 25412 9522 25464 9528
rect 25228 8900 25280 8906
rect 25228 8842 25280 8848
rect 25240 8634 25268 8842
rect 25412 8832 25464 8838
rect 25412 8774 25464 8780
rect 25424 8634 25452 8774
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25516 7410 25544 9998
rect 25608 9586 25636 10066
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25608 9042 25636 9522
rect 25744 9276 26052 9285
rect 25744 9274 25750 9276
rect 25806 9274 25830 9276
rect 25886 9274 25910 9276
rect 25966 9274 25990 9276
rect 26046 9274 26052 9276
rect 25806 9222 25808 9274
rect 25988 9222 25990 9274
rect 25744 9220 25750 9222
rect 25806 9220 25830 9222
rect 25886 9220 25910 9222
rect 25966 9220 25990 9222
rect 26046 9220 26052 9222
rect 25744 9211 26052 9220
rect 25596 9036 25648 9042
rect 25596 8978 25648 8984
rect 25608 8498 25636 8978
rect 25596 8492 25648 8498
rect 25596 8434 25648 8440
rect 25596 8356 25648 8362
rect 25596 8298 25648 8304
rect 25608 8090 25636 8298
rect 25744 8188 26052 8197
rect 25744 8186 25750 8188
rect 25806 8186 25830 8188
rect 25886 8186 25910 8188
rect 25966 8186 25990 8188
rect 26046 8186 26052 8188
rect 25806 8134 25808 8186
rect 25988 8134 25990 8186
rect 25744 8132 25750 8134
rect 25806 8132 25830 8134
rect 25886 8132 25910 8134
rect 25966 8132 25990 8134
rect 26046 8132 26052 8134
rect 25744 8123 26052 8132
rect 26160 8090 26188 12038
rect 26436 8974 26464 16390
rect 26516 13864 26568 13870
rect 26516 13806 26568 13812
rect 26528 13530 26556 13806
rect 26516 13524 26568 13530
rect 26516 13466 26568 13472
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26620 12986 26648 13262
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26712 12170 26740 18158
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 26804 16726 26832 16934
rect 26792 16720 26844 16726
rect 26792 16662 26844 16668
rect 26804 16522 26832 16662
rect 26792 16516 26844 16522
rect 26792 16458 26844 16464
rect 26896 16402 26924 21422
rect 26988 21078 27016 21830
rect 26976 21072 27028 21078
rect 26976 21014 27028 21020
rect 26976 20528 27028 20534
rect 26976 20470 27028 20476
rect 26988 17542 27016 20470
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 27080 18086 27108 18566
rect 27172 18290 27200 18566
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27068 18080 27120 18086
rect 27068 18022 27120 18028
rect 26976 17536 27028 17542
rect 26976 17478 27028 17484
rect 26804 16374 26924 16402
rect 26700 12164 26752 12170
rect 26700 12106 26752 12112
rect 26712 11694 26740 12106
rect 26700 11688 26752 11694
rect 26700 11630 26752 11636
rect 26516 9920 26568 9926
rect 26516 9862 26568 9868
rect 26528 9625 26556 9862
rect 26514 9616 26570 9625
rect 26514 9551 26570 9560
rect 26424 8968 26476 8974
rect 26424 8910 26476 8916
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 25976 7546 26004 7686
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 25504 7404 25556 7410
rect 25504 7346 25556 7352
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 25608 7002 25636 7142
rect 25744 7100 26052 7109
rect 25744 7098 25750 7100
rect 25806 7098 25830 7100
rect 25886 7098 25910 7100
rect 25966 7098 25990 7100
rect 26046 7098 26052 7100
rect 25806 7046 25808 7098
rect 25988 7046 25990 7098
rect 25744 7044 25750 7046
rect 25806 7044 25830 7046
rect 25886 7044 25910 7046
rect 25966 7044 25990 7046
rect 26046 7044 26052 7046
rect 25744 7035 26052 7044
rect 25596 6996 25648 7002
rect 25596 6938 25648 6944
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 25240 6186 25268 6598
rect 25228 6180 25280 6186
rect 25228 6122 25280 6128
rect 25744 6012 26052 6021
rect 25744 6010 25750 6012
rect 25806 6010 25830 6012
rect 25886 6010 25910 6012
rect 25966 6010 25990 6012
rect 26046 6010 26052 6012
rect 25806 5958 25808 6010
rect 25988 5958 25990 6010
rect 25744 5956 25750 5958
rect 25806 5956 25830 5958
rect 25886 5956 25910 5958
rect 25966 5956 25990 5958
rect 26046 5956 26052 5958
rect 25744 5947 26052 5956
rect 26804 5914 26832 16374
rect 27080 16250 27108 18022
rect 27264 17202 27292 21830
rect 27540 21486 27568 23462
rect 27724 23118 27752 25706
rect 28264 25152 28316 25158
rect 28264 25094 28316 25100
rect 27896 24404 27948 24410
rect 27896 24346 27948 24352
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27816 23186 27844 24006
rect 27804 23180 27856 23186
rect 27804 23122 27856 23128
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27620 21616 27672 21622
rect 27620 21558 27672 21564
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 27540 20806 27568 21422
rect 27632 21026 27660 21558
rect 27724 21146 27752 23054
rect 27712 21140 27764 21146
rect 27712 21082 27764 21088
rect 27632 21010 27752 21026
rect 27632 21004 27764 21010
rect 27632 20998 27712 21004
rect 27712 20946 27764 20952
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27528 20800 27580 20806
rect 27528 20742 27580 20748
rect 27632 20534 27660 20878
rect 27620 20528 27672 20534
rect 27620 20470 27672 20476
rect 27724 19394 27752 20946
rect 27816 20806 27844 23122
rect 27908 22438 27936 24346
rect 28276 23730 28304 25094
rect 28264 23724 28316 23730
rect 28264 23666 28316 23672
rect 28080 23180 28132 23186
rect 28080 23122 28132 23128
rect 28092 22642 28120 23122
rect 28276 22681 28304 23666
rect 28262 22672 28318 22681
rect 28080 22636 28132 22642
rect 28262 22607 28318 22616
rect 28080 22578 28132 22584
rect 27896 22432 27948 22438
rect 27896 22374 27948 22380
rect 27804 20800 27856 20806
rect 27804 20742 27856 20748
rect 27816 19990 27844 20742
rect 27804 19984 27856 19990
rect 27804 19926 27856 19932
rect 27816 19514 27844 19926
rect 27804 19508 27856 19514
rect 27804 19450 27856 19456
rect 27632 19366 27752 19394
rect 27436 19168 27488 19174
rect 27436 19110 27488 19116
rect 27252 17196 27304 17202
rect 27252 17138 27304 17144
rect 27448 16794 27476 19110
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 27540 17202 27568 18226
rect 27632 17218 27660 19366
rect 27712 19304 27764 19310
rect 27712 19246 27764 19252
rect 27724 18766 27752 19246
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 27724 18426 27752 18702
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 27816 17882 27844 19450
rect 27804 17876 27856 17882
rect 27804 17818 27856 17824
rect 27816 17678 27844 17818
rect 27908 17746 27936 22374
rect 28092 22098 28120 22578
rect 28080 22092 28132 22098
rect 28080 22034 28132 22040
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 28000 21690 28028 21830
rect 27988 21684 28040 21690
rect 27988 21626 28040 21632
rect 28092 21010 28120 22034
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28080 21004 28132 21010
rect 28080 20946 28132 20952
rect 27988 20256 28040 20262
rect 27988 20198 28040 20204
rect 28000 19854 28028 20198
rect 27988 19848 28040 19854
rect 27986 19816 27988 19825
rect 28040 19816 28042 19825
rect 27986 19751 28042 19760
rect 28000 18970 28028 19751
rect 28092 19310 28120 20946
rect 28184 20924 28212 21082
rect 28264 20936 28316 20942
rect 28184 20896 28264 20924
rect 28184 20262 28212 20896
rect 28264 20878 28316 20884
rect 28172 20256 28224 20262
rect 28172 20198 28224 20204
rect 28184 19718 28212 20198
rect 28172 19712 28224 19718
rect 28172 19654 28224 19660
rect 28184 19378 28212 19654
rect 28172 19372 28224 19378
rect 28172 19314 28224 19320
rect 28080 19304 28132 19310
rect 28080 19246 28132 19252
rect 27988 18964 28040 18970
rect 27988 18906 28040 18912
rect 28092 18902 28120 19246
rect 28172 19168 28224 19174
rect 28172 19110 28224 19116
rect 28080 18896 28132 18902
rect 28080 18838 28132 18844
rect 28184 18630 28212 19110
rect 28172 18624 28224 18630
rect 28172 18566 28224 18572
rect 27896 17740 27948 17746
rect 27896 17682 27948 17688
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27908 17338 27936 17682
rect 27896 17332 27948 17338
rect 27896 17274 27948 17280
rect 27528 17196 27580 17202
rect 27632 17190 27844 17218
rect 27528 17138 27580 17144
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27540 16674 27568 17138
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27448 16646 27568 16674
rect 27632 16658 27660 17070
rect 27620 16652 27672 16658
rect 27068 16244 27120 16250
rect 27068 16186 27120 16192
rect 27264 16046 27292 16594
rect 27448 16590 27476 16646
rect 27620 16594 27672 16600
rect 27436 16584 27488 16590
rect 27436 16526 27488 16532
rect 27344 16516 27396 16522
rect 27344 16458 27396 16464
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 27264 15502 27292 15982
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27356 15162 27384 16458
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27448 15042 27476 16526
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27356 15026 27476 15042
rect 27344 15020 27476 15026
rect 27396 15014 27476 15020
rect 27344 14962 27396 14968
rect 27356 14550 27384 14962
rect 27540 14958 27568 15302
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27344 14544 27396 14550
rect 27344 14486 27396 14492
rect 27448 14006 27476 14894
rect 27436 14000 27488 14006
rect 27436 13942 27488 13948
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 26884 12980 26936 12986
rect 26884 12922 26936 12928
rect 26896 10062 26924 12922
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27264 11898 27292 12786
rect 27252 11892 27304 11898
rect 27252 11834 27304 11840
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 27172 10674 27200 11154
rect 27356 11150 27384 13874
rect 27344 11144 27396 11150
rect 27344 11086 27396 11092
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 27172 7342 27200 10610
rect 27448 8634 27476 13942
rect 27540 12850 27568 14894
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27632 13802 27660 14214
rect 27620 13796 27672 13802
rect 27620 13738 27672 13744
rect 27724 12986 27752 16050
rect 27816 14618 27844 17190
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27908 14482 27936 17274
rect 28080 16652 28132 16658
rect 28080 16594 28132 16600
rect 28092 16046 28120 16594
rect 28080 16040 28132 16046
rect 28080 15982 28132 15988
rect 27896 14476 27948 14482
rect 27948 14436 28028 14464
rect 27896 14418 27948 14424
rect 27712 12980 27764 12986
rect 27712 12922 27764 12928
rect 27528 12844 27580 12850
rect 27528 12786 27580 12792
rect 27896 12844 27948 12850
rect 27896 12786 27948 12792
rect 27712 12776 27764 12782
rect 27712 12718 27764 12724
rect 27620 12096 27672 12102
rect 27620 12038 27672 12044
rect 27632 11354 27660 12038
rect 27724 11898 27752 12718
rect 27712 11892 27764 11898
rect 27712 11834 27764 11840
rect 27724 11778 27752 11834
rect 27724 11750 27844 11778
rect 27712 11688 27764 11694
rect 27712 11630 27764 11636
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27724 10810 27752 11630
rect 27816 11354 27844 11750
rect 27804 11348 27856 11354
rect 27804 11290 27856 11296
rect 27804 11076 27856 11082
rect 27804 11018 27856 11024
rect 27712 10804 27764 10810
rect 27712 10746 27764 10752
rect 27724 10062 27752 10746
rect 27816 10674 27844 11018
rect 27804 10668 27856 10674
rect 27804 10610 27856 10616
rect 27804 10464 27856 10470
rect 27804 10406 27856 10412
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27620 9988 27672 9994
rect 27620 9930 27672 9936
rect 27632 9738 27660 9930
rect 27540 9710 27660 9738
rect 27816 9722 27844 10406
rect 27804 9716 27856 9722
rect 27436 8628 27488 8634
rect 27436 8570 27488 8576
rect 27540 8430 27568 9710
rect 27804 9658 27856 9664
rect 27620 9444 27672 9450
rect 27620 9386 27672 9392
rect 27632 9178 27660 9386
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 27436 8424 27488 8430
rect 27436 8366 27488 8372
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27448 7886 27476 8366
rect 27540 8022 27568 8366
rect 27528 8016 27580 8022
rect 27528 7958 27580 7964
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 27448 7546 27476 7822
rect 27436 7540 27488 7546
rect 27436 7482 27488 7488
rect 27160 7336 27212 7342
rect 27160 7278 27212 7284
rect 27068 7200 27120 7206
rect 27068 7142 27120 7148
rect 27080 7002 27108 7142
rect 27068 6996 27120 7002
rect 27068 6938 27120 6944
rect 27632 6866 27660 9114
rect 27908 8945 27936 12786
rect 28000 12594 28028 14436
rect 28092 13870 28120 15982
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 28184 13818 28212 18566
rect 28368 17814 28396 26250
rect 28644 25945 28672 26250
rect 28630 25936 28686 25945
rect 28630 25871 28686 25880
rect 28540 25696 28592 25702
rect 28540 25638 28592 25644
rect 28448 25492 28500 25498
rect 28448 25434 28500 25440
rect 28460 23186 28488 25434
rect 28552 24614 28580 25638
rect 28540 24608 28592 24614
rect 28540 24550 28592 24556
rect 28552 24070 28580 24550
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28724 24064 28776 24070
rect 28724 24006 28776 24012
rect 28448 23180 28500 23186
rect 28448 23122 28500 23128
rect 28460 21962 28488 23122
rect 28552 23118 28580 24006
rect 28632 23520 28684 23526
rect 28632 23462 28684 23468
rect 28644 23225 28672 23462
rect 28630 23216 28686 23225
rect 28630 23151 28686 23160
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28460 20330 28488 21898
rect 28552 21690 28580 23054
rect 28540 21684 28592 21690
rect 28540 21626 28592 21632
rect 28736 21554 28764 24006
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 28736 21185 28764 21490
rect 28722 21176 28778 21185
rect 28722 21111 28778 21120
rect 28448 20324 28500 20330
rect 28448 20266 28500 20272
rect 28460 19174 28488 20266
rect 28448 19168 28500 19174
rect 28448 19110 28500 19116
rect 28722 19136 28778 19145
rect 28722 19071 28778 19080
rect 28736 18766 28764 19071
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 28736 17882 28764 18702
rect 28724 17876 28776 17882
rect 28724 17818 28776 17824
rect 28356 17808 28408 17814
rect 28356 17750 28408 17756
rect 28356 17536 28408 17542
rect 28356 17478 28408 17484
rect 28368 16114 28396 17478
rect 28724 16584 28776 16590
rect 28722 16552 28724 16561
rect 28776 16552 28778 16561
rect 28722 16487 28778 16496
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28264 16040 28316 16046
rect 28264 15982 28316 15988
rect 28276 14822 28304 15982
rect 28736 15706 28764 16487
rect 28724 15700 28776 15706
rect 28724 15642 28776 15648
rect 28264 14816 28316 14822
rect 28264 14758 28316 14764
rect 28276 13938 28304 14758
rect 28630 14376 28686 14385
rect 28630 14311 28686 14320
rect 28644 14074 28672 14311
rect 28632 14068 28684 14074
rect 28632 14010 28684 14016
rect 28446 13968 28502 13977
rect 28264 13932 28316 13938
rect 28446 13903 28448 13912
rect 28264 13874 28316 13880
rect 28500 13903 28502 13912
rect 28448 13874 28500 13880
rect 28092 12730 28120 13806
rect 28184 13790 28396 13818
rect 28172 13184 28224 13190
rect 28172 13126 28224 13132
rect 28184 12850 28212 13126
rect 28172 12844 28224 12850
rect 28172 12786 28224 12792
rect 28264 12776 28316 12782
rect 28092 12702 28212 12730
rect 28264 12718 28316 12724
rect 28000 12566 28120 12594
rect 27986 12472 28042 12481
rect 27986 12407 28042 12416
rect 27894 8936 27950 8945
rect 27894 8871 27950 8880
rect 27712 7812 27764 7818
rect 27712 7754 27764 7760
rect 27724 7546 27752 7754
rect 27712 7540 27764 7546
rect 27712 7482 27764 7488
rect 27896 7200 27948 7206
rect 27896 7142 27948 7148
rect 27908 7002 27936 7142
rect 27896 6996 27948 7002
rect 27896 6938 27948 6944
rect 27528 6860 27580 6866
rect 27528 6802 27580 6808
rect 27620 6860 27672 6866
rect 27620 6802 27672 6808
rect 27540 6746 27568 6802
rect 27540 6718 27660 6746
rect 26976 6656 27028 6662
rect 26976 6598 27028 6604
rect 26988 6458 27016 6598
rect 26976 6452 27028 6458
rect 26976 6394 27028 6400
rect 27632 6390 27660 6718
rect 27712 6656 27764 6662
rect 27712 6598 27764 6604
rect 27724 6458 27752 6598
rect 27712 6452 27764 6458
rect 27712 6394 27764 6400
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 26792 5908 26844 5914
rect 26792 5850 26844 5856
rect 25744 4924 26052 4933
rect 25744 4922 25750 4924
rect 25806 4922 25830 4924
rect 25886 4922 25910 4924
rect 25966 4922 25990 4924
rect 26046 4922 26052 4924
rect 25806 4870 25808 4922
rect 25988 4870 25990 4922
rect 25744 4868 25750 4870
rect 25806 4868 25830 4870
rect 25886 4868 25910 4870
rect 25966 4868 25990 4870
rect 26046 4868 26052 4870
rect 25744 4859 26052 4868
rect 25744 3836 26052 3845
rect 25744 3834 25750 3836
rect 25806 3834 25830 3836
rect 25886 3834 25910 3836
rect 25966 3834 25990 3836
rect 26046 3834 26052 3836
rect 25806 3782 25808 3834
rect 25988 3782 25990 3834
rect 25744 3780 25750 3782
rect 25806 3780 25830 3782
rect 25886 3780 25910 3782
rect 25966 3780 25990 3782
rect 26046 3780 26052 3782
rect 25744 3771 26052 3780
rect 27436 3392 27488 3398
rect 27436 3334 27488 3340
rect 24044 2746 24164 2774
rect 25744 2748 26052 2757
rect 25744 2746 25750 2748
rect 25806 2746 25830 2748
rect 25886 2746 25910 2748
rect 25966 2746 25990 2748
rect 26046 2746 26052 2748
rect 24044 2582 24072 2746
rect 25806 2694 25808 2746
rect 25988 2694 25990 2746
rect 25744 2692 25750 2694
rect 25806 2692 25830 2694
rect 25886 2692 25910 2694
rect 25966 2692 25990 2694
rect 26046 2692 26052 2694
rect 25744 2683 26052 2692
rect 22928 2576 22980 2582
rect 22928 2518 22980 2524
rect 24032 2576 24084 2582
rect 24032 2518 24084 2524
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 19892 2372 19944 2378
rect 19892 2314 19944 2320
rect 23204 2372 23256 2378
rect 23204 2314 23256 2320
rect 25136 2372 25188 2378
rect 25136 2314 25188 2320
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 21284 800 21312 2246
rect 22202 2204 22510 2213
rect 22202 2202 22208 2204
rect 22264 2202 22288 2204
rect 22344 2202 22368 2204
rect 22424 2202 22448 2204
rect 22504 2202 22510 2204
rect 22264 2150 22266 2202
rect 22446 2150 22448 2202
rect 22202 2148 22208 2150
rect 22264 2148 22288 2150
rect 22344 2148 22368 2150
rect 22424 2148 22448 2150
rect 22504 2148 22510 2150
rect 22202 2139 22510 2148
rect 23216 800 23244 2314
rect 25148 800 25176 2314
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 5814 0 5870 800
rect 8390 0 8446 800
rect 10322 0 10378 800
rect 12254 0 12310 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 18694 0 18750 800
rect 21270 0 21326 800
rect 23202 0 23258 800
rect 25134 0 25190 800
rect 27448 785 27476 3334
rect 28000 2650 28028 12407
rect 28092 12306 28120 12566
rect 28184 12374 28212 12702
rect 28172 12368 28224 12374
rect 28172 12310 28224 12316
rect 28080 12300 28132 12306
rect 28080 12242 28132 12248
rect 28092 11898 28120 12242
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 28092 9518 28120 11834
rect 28184 11218 28212 12310
rect 28276 11694 28304 12718
rect 28368 12481 28396 13790
rect 28460 13530 28488 13874
rect 28448 13524 28500 13530
rect 28448 13466 28500 13472
rect 28632 12640 28684 12646
rect 28632 12582 28684 12588
rect 28354 12472 28410 12481
rect 28354 12407 28410 12416
rect 28644 12345 28672 12582
rect 28630 12336 28686 12345
rect 28630 12271 28686 12280
rect 28356 12164 28408 12170
rect 28356 12106 28408 12112
rect 28264 11688 28316 11694
rect 28264 11630 28316 11636
rect 28172 11212 28224 11218
rect 28172 11154 28224 11160
rect 28276 10742 28304 11630
rect 28264 10736 28316 10742
rect 28264 10678 28316 10684
rect 28172 10532 28224 10538
rect 28172 10474 28224 10480
rect 28184 10130 28212 10474
rect 28276 10130 28304 10678
rect 28172 10124 28224 10130
rect 28172 10066 28224 10072
rect 28264 10124 28316 10130
rect 28264 10066 28316 10072
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 28092 9178 28120 9454
rect 28368 9330 28396 12106
rect 28722 9616 28778 9625
rect 28722 9551 28724 9560
rect 28776 9551 28778 9560
rect 28724 9522 28776 9528
rect 28276 9302 28396 9330
rect 28540 9376 28592 9382
rect 28540 9318 28592 9324
rect 28080 9172 28132 9178
rect 28080 9114 28132 9120
rect 28172 9104 28224 9110
rect 28172 9046 28224 9052
rect 28080 6860 28132 6866
rect 28080 6802 28132 6808
rect 28092 6458 28120 6802
rect 28184 6730 28212 9046
rect 28172 6724 28224 6730
rect 28172 6666 28224 6672
rect 28080 6452 28132 6458
rect 28080 6394 28132 6400
rect 28184 5846 28212 6666
rect 28276 6662 28304 9302
rect 28356 9172 28408 9178
rect 28356 9114 28408 9120
rect 28368 6866 28396 9114
rect 28552 9110 28580 9318
rect 28736 9178 28764 9522
rect 28828 9450 28856 29446
rect 29286 29404 29594 29413
rect 29286 29402 29292 29404
rect 29348 29402 29372 29404
rect 29428 29402 29452 29404
rect 29508 29402 29532 29404
rect 29588 29402 29594 29404
rect 29348 29350 29350 29402
rect 29530 29350 29532 29402
rect 29286 29348 29292 29350
rect 29348 29348 29372 29350
rect 29428 29348 29452 29350
rect 29508 29348 29532 29350
rect 29588 29348 29594 29350
rect 29286 29339 29594 29348
rect 29286 28316 29594 28325
rect 29286 28314 29292 28316
rect 29348 28314 29372 28316
rect 29428 28314 29452 28316
rect 29508 28314 29532 28316
rect 29588 28314 29594 28316
rect 29348 28262 29350 28314
rect 29530 28262 29532 28314
rect 29286 28260 29292 28262
rect 29348 28260 29372 28262
rect 29428 28260 29452 28262
rect 29508 28260 29532 28262
rect 29588 28260 29594 28262
rect 29286 28251 29594 28260
rect 29286 27228 29594 27237
rect 29286 27226 29292 27228
rect 29348 27226 29372 27228
rect 29428 27226 29452 27228
rect 29508 27226 29532 27228
rect 29588 27226 29594 27228
rect 29348 27174 29350 27226
rect 29530 27174 29532 27226
rect 29286 27172 29292 27174
rect 29348 27172 29372 27174
rect 29428 27172 29452 27174
rect 29508 27172 29532 27174
rect 29588 27172 29594 27174
rect 29286 27163 29594 27172
rect 29286 26140 29594 26149
rect 29286 26138 29292 26140
rect 29348 26138 29372 26140
rect 29428 26138 29452 26140
rect 29508 26138 29532 26140
rect 29588 26138 29594 26140
rect 29348 26086 29350 26138
rect 29530 26086 29532 26138
rect 29286 26084 29292 26086
rect 29348 26084 29372 26086
rect 29428 26084 29452 26086
rect 29508 26084 29532 26086
rect 29588 26084 29594 26086
rect 29286 26075 29594 26084
rect 29286 25052 29594 25061
rect 29286 25050 29292 25052
rect 29348 25050 29372 25052
rect 29428 25050 29452 25052
rect 29508 25050 29532 25052
rect 29588 25050 29594 25052
rect 29348 24998 29350 25050
rect 29530 24998 29532 25050
rect 29286 24996 29292 24998
rect 29348 24996 29372 24998
rect 29428 24996 29452 24998
rect 29508 24996 29532 24998
rect 29588 24996 29594 24998
rect 29286 24987 29594 24996
rect 29286 23964 29594 23973
rect 29286 23962 29292 23964
rect 29348 23962 29372 23964
rect 29428 23962 29452 23964
rect 29508 23962 29532 23964
rect 29588 23962 29594 23964
rect 29348 23910 29350 23962
rect 29530 23910 29532 23962
rect 29286 23908 29292 23910
rect 29348 23908 29372 23910
rect 29428 23908 29452 23910
rect 29508 23908 29532 23910
rect 29588 23908 29594 23910
rect 29286 23899 29594 23908
rect 29286 22876 29594 22885
rect 29286 22874 29292 22876
rect 29348 22874 29372 22876
rect 29428 22874 29452 22876
rect 29508 22874 29532 22876
rect 29588 22874 29594 22876
rect 29348 22822 29350 22874
rect 29530 22822 29532 22874
rect 29286 22820 29292 22822
rect 29348 22820 29372 22822
rect 29428 22820 29452 22822
rect 29508 22820 29532 22822
rect 29588 22820 29594 22822
rect 29286 22811 29594 22820
rect 29286 21788 29594 21797
rect 29286 21786 29292 21788
rect 29348 21786 29372 21788
rect 29428 21786 29452 21788
rect 29508 21786 29532 21788
rect 29588 21786 29594 21788
rect 29348 21734 29350 21786
rect 29530 21734 29532 21786
rect 29286 21732 29292 21734
rect 29348 21732 29372 21734
rect 29428 21732 29452 21734
rect 29508 21732 29532 21734
rect 29588 21732 29594 21734
rect 29286 21723 29594 21732
rect 29286 20700 29594 20709
rect 29286 20698 29292 20700
rect 29348 20698 29372 20700
rect 29428 20698 29452 20700
rect 29508 20698 29532 20700
rect 29588 20698 29594 20700
rect 29348 20646 29350 20698
rect 29530 20646 29532 20698
rect 29286 20644 29292 20646
rect 29348 20644 29372 20646
rect 29428 20644 29452 20646
rect 29508 20644 29532 20646
rect 29588 20644 29594 20646
rect 29286 20635 29594 20644
rect 29286 19612 29594 19621
rect 29286 19610 29292 19612
rect 29348 19610 29372 19612
rect 29428 19610 29452 19612
rect 29508 19610 29532 19612
rect 29588 19610 29594 19612
rect 29348 19558 29350 19610
rect 29530 19558 29532 19610
rect 29286 19556 29292 19558
rect 29348 19556 29372 19558
rect 29428 19556 29452 19558
rect 29508 19556 29532 19558
rect 29588 19556 29594 19558
rect 29286 19547 29594 19556
rect 29286 18524 29594 18533
rect 29286 18522 29292 18524
rect 29348 18522 29372 18524
rect 29428 18522 29452 18524
rect 29508 18522 29532 18524
rect 29588 18522 29594 18524
rect 29348 18470 29350 18522
rect 29530 18470 29532 18522
rect 29286 18468 29292 18470
rect 29348 18468 29372 18470
rect 29428 18468 29452 18470
rect 29508 18468 29532 18470
rect 29588 18468 29594 18470
rect 29286 18459 29594 18468
rect 29286 17436 29594 17445
rect 29286 17434 29292 17436
rect 29348 17434 29372 17436
rect 29428 17434 29452 17436
rect 29508 17434 29532 17436
rect 29588 17434 29594 17436
rect 29348 17382 29350 17434
rect 29530 17382 29532 17434
rect 29286 17380 29292 17382
rect 29348 17380 29372 17382
rect 29428 17380 29452 17382
rect 29508 17380 29532 17382
rect 29588 17380 29594 17382
rect 29286 17371 29594 17380
rect 29286 16348 29594 16357
rect 29286 16346 29292 16348
rect 29348 16346 29372 16348
rect 29428 16346 29452 16348
rect 29508 16346 29532 16348
rect 29588 16346 29594 16348
rect 29348 16294 29350 16346
rect 29530 16294 29532 16346
rect 29286 16292 29292 16294
rect 29348 16292 29372 16294
rect 29428 16292 29452 16294
rect 29508 16292 29532 16294
rect 29588 16292 29594 16294
rect 29286 16283 29594 16292
rect 29286 15260 29594 15269
rect 29286 15258 29292 15260
rect 29348 15258 29372 15260
rect 29428 15258 29452 15260
rect 29508 15258 29532 15260
rect 29588 15258 29594 15260
rect 29348 15206 29350 15258
rect 29530 15206 29532 15258
rect 29286 15204 29292 15206
rect 29348 15204 29372 15206
rect 29428 15204 29452 15206
rect 29508 15204 29532 15206
rect 29588 15204 29594 15206
rect 29286 15195 29594 15204
rect 29286 14172 29594 14181
rect 29286 14170 29292 14172
rect 29348 14170 29372 14172
rect 29428 14170 29452 14172
rect 29508 14170 29532 14172
rect 29588 14170 29594 14172
rect 29348 14118 29350 14170
rect 29530 14118 29532 14170
rect 29286 14116 29292 14118
rect 29348 14116 29372 14118
rect 29428 14116 29452 14118
rect 29508 14116 29532 14118
rect 29588 14116 29594 14118
rect 29286 14107 29594 14116
rect 29286 13084 29594 13093
rect 29286 13082 29292 13084
rect 29348 13082 29372 13084
rect 29428 13082 29452 13084
rect 29508 13082 29532 13084
rect 29588 13082 29594 13084
rect 29348 13030 29350 13082
rect 29530 13030 29532 13082
rect 29286 13028 29292 13030
rect 29348 13028 29372 13030
rect 29428 13028 29452 13030
rect 29508 13028 29532 13030
rect 29588 13028 29594 13030
rect 29286 13019 29594 13028
rect 29286 11996 29594 12005
rect 29286 11994 29292 11996
rect 29348 11994 29372 11996
rect 29428 11994 29452 11996
rect 29508 11994 29532 11996
rect 29588 11994 29594 11996
rect 29348 11942 29350 11994
rect 29530 11942 29532 11994
rect 29286 11940 29292 11942
rect 29348 11940 29372 11942
rect 29428 11940 29452 11942
rect 29508 11940 29532 11942
rect 29588 11940 29594 11942
rect 29286 11931 29594 11940
rect 29286 10908 29594 10917
rect 29286 10906 29292 10908
rect 29348 10906 29372 10908
rect 29428 10906 29452 10908
rect 29508 10906 29532 10908
rect 29588 10906 29594 10908
rect 29348 10854 29350 10906
rect 29530 10854 29532 10906
rect 29286 10852 29292 10854
rect 29348 10852 29372 10854
rect 29428 10852 29452 10854
rect 29508 10852 29532 10854
rect 29588 10852 29594 10854
rect 29286 10843 29594 10852
rect 29286 9820 29594 9829
rect 29286 9818 29292 9820
rect 29348 9818 29372 9820
rect 29428 9818 29452 9820
rect 29508 9818 29532 9820
rect 29588 9818 29594 9820
rect 29348 9766 29350 9818
rect 29530 9766 29532 9818
rect 29286 9764 29292 9766
rect 29348 9764 29372 9766
rect 29428 9764 29452 9766
rect 29508 9764 29532 9766
rect 29588 9764 29594 9766
rect 29286 9755 29594 9764
rect 28816 9444 28868 9450
rect 28816 9386 28868 9392
rect 28724 9172 28776 9178
rect 28724 9114 28776 9120
rect 28540 9104 28592 9110
rect 28540 9046 28592 9052
rect 29286 8732 29594 8741
rect 29286 8730 29292 8732
rect 29348 8730 29372 8732
rect 29428 8730 29452 8732
rect 29508 8730 29532 8732
rect 29588 8730 29594 8732
rect 29348 8678 29350 8730
rect 29530 8678 29532 8730
rect 29286 8676 29292 8678
rect 29348 8676 29372 8678
rect 29428 8676 29452 8678
rect 29508 8676 29532 8678
rect 29588 8676 29594 8678
rect 29286 8667 29594 8676
rect 28448 7812 28500 7818
rect 28448 7754 28500 7760
rect 28724 7812 28776 7818
rect 28724 7754 28776 7760
rect 28356 6860 28408 6866
rect 28356 6802 28408 6808
rect 28264 6656 28316 6662
rect 28264 6598 28316 6604
rect 28368 6390 28396 6802
rect 28460 6798 28488 7754
rect 28736 7478 28764 7754
rect 29286 7644 29594 7653
rect 29286 7642 29292 7644
rect 29348 7642 29372 7644
rect 29428 7642 29452 7644
rect 29508 7642 29532 7644
rect 29588 7642 29594 7644
rect 29348 7590 29350 7642
rect 29530 7590 29532 7642
rect 29286 7588 29292 7590
rect 29348 7588 29372 7590
rect 29428 7588 29452 7590
rect 29508 7588 29532 7590
rect 29588 7588 29594 7590
rect 29286 7579 29594 7588
rect 28724 7472 28776 7478
rect 28722 7440 28724 7449
rect 28776 7440 28778 7449
rect 28722 7375 28778 7384
rect 28448 6792 28500 6798
rect 28448 6734 28500 6740
rect 29286 6556 29594 6565
rect 29286 6554 29292 6556
rect 29348 6554 29372 6556
rect 29428 6554 29452 6556
rect 29508 6554 29532 6556
rect 29588 6554 29594 6556
rect 29348 6502 29350 6554
rect 29530 6502 29532 6554
rect 29286 6500 29292 6502
rect 29348 6500 29372 6502
rect 29428 6500 29452 6502
rect 29508 6500 29532 6502
rect 29588 6500 29594 6502
rect 29286 6491 29594 6500
rect 28356 6384 28408 6390
rect 28356 6326 28408 6332
rect 28172 5840 28224 5846
rect 28172 5782 28224 5788
rect 28724 5704 28776 5710
rect 28724 5646 28776 5652
rect 28736 5370 28764 5646
rect 29286 5468 29594 5477
rect 29286 5466 29292 5468
rect 29348 5466 29372 5468
rect 29428 5466 29452 5468
rect 29508 5466 29532 5468
rect 29588 5466 29594 5468
rect 29348 5414 29350 5466
rect 29530 5414 29532 5466
rect 29286 5412 29292 5414
rect 29348 5412 29372 5414
rect 29428 5412 29452 5414
rect 29508 5412 29532 5414
rect 29588 5412 29594 5414
rect 29286 5403 29594 5412
rect 28724 5364 28776 5370
rect 28724 5306 28776 5312
rect 28736 5273 28764 5306
rect 28722 5264 28778 5273
rect 28722 5199 28778 5208
rect 29286 4380 29594 4389
rect 29286 4378 29292 4380
rect 29348 4378 29372 4380
rect 29428 4378 29452 4380
rect 29508 4378 29532 4380
rect 29588 4378 29594 4380
rect 29348 4326 29350 4378
rect 29530 4326 29532 4378
rect 29286 4324 29292 4326
rect 29348 4324 29372 4326
rect 29428 4324 29452 4326
rect 29508 4324 29532 4326
rect 29588 4324 29594 4326
rect 29286 4315 29594 4324
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28644 3058 28672 3878
rect 29286 3292 29594 3301
rect 29286 3290 29292 3292
rect 29348 3290 29372 3292
rect 29428 3290 29452 3292
rect 29508 3290 29532 3292
rect 29588 3290 29594 3292
rect 29348 3238 29350 3290
rect 29530 3238 29532 3290
rect 29286 3236 29292 3238
rect 29348 3236 29372 3238
rect 29428 3236 29452 3238
rect 29508 3236 29532 3238
rect 29588 3236 29594 3238
rect 29286 3227 29594 3236
rect 28632 3052 28684 3058
rect 28632 2994 28684 3000
rect 28644 2825 28672 2994
rect 29644 2916 29696 2922
rect 29644 2858 29696 2864
rect 28630 2816 28686 2825
rect 28630 2751 28686 2760
rect 27988 2644 28040 2650
rect 27988 2586 28040 2592
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 27724 800 27752 2314
rect 29286 2204 29594 2213
rect 29286 2202 29292 2204
rect 29348 2202 29372 2204
rect 29428 2202 29452 2204
rect 29508 2202 29532 2204
rect 29588 2202 29594 2204
rect 29348 2150 29350 2202
rect 29530 2150 29532 2202
rect 29286 2148 29292 2150
rect 29348 2148 29372 2150
rect 29428 2148 29452 2150
rect 29508 2148 29532 2150
rect 29588 2148 29594 2150
rect 29286 2139 29594 2148
rect 29656 800 29684 2858
rect 27434 776 27490 785
rect 27434 711 27490 720
rect 27710 0 27766 800
rect 29642 0 29698 800
<< via2 >>
rect 1858 31320 1914 31376
rect 1490 29280 1546 29336
rect 1582 26580 1638 26616
rect 1582 26560 1584 26580
rect 1584 26560 1636 26580
rect 1636 26560 1638 26580
rect 1398 24520 1454 24576
rect 1582 22480 1638 22536
rect 1766 22500 1822 22536
rect 1766 22480 1768 22500
rect 1768 22480 1820 22500
rect 1820 22480 1822 22500
rect 8040 30490 8096 30492
rect 8120 30490 8176 30492
rect 8200 30490 8256 30492
rect 8280 30490 8336 30492
rect 8040 30438 8086 30490
rect 8086 30438 8096 30490
rect 8120 30438 8150 30490
rect 8150 30438 8162 30490
rect 8162 30438 8176 30490
rect 8200 30438 8214 30490
rect 8214 30438 8226 30490
rect 8226 30438 8256 30490
rect 8280 30438 8290 30490
rect 8290 30438 8336 30490
rect 8040 30436 8096 30438
rect 8120 30436 8176 30438
rect 8200 30436 8256 30438
rect 8280 30436 8336 30438
rect 4498 29946 4554 29948
rect 4578 29946 4634 29948
rect 4658 29946 4714 29948
rect 4738 29946 4794 29948
rect 4498 29894 4544 29946
rect 4544 29894 4554 29946
rect 4578 29894 4608 29946
rect 4608 29894 4620 29946
rect 4620 29894 4634 29946
rect 4658 29894 4672 29946
rect 4672 29894 4684 29946
rect 4684 29894 4714 29946
rect 4738 29894 4748 29946
rect 4748 29894 4794 29946
rect 4498 29892 4554 29894
rect 4578 29892 4634 29894
rect 4658 29892 4714 29894
rect 4738 29892 4794 29894
rect 1490 19760 1546 19816
rect 1398 15680 1454 15736
rect 1582 17756 1584 17776
rect 1584 17756 1636 17776
rect 1636 17756 1638 17776
rect 1582 17720 1638 17756
rect 1490 12960 1546 13016
rect 1490 10920 1546 10976
rect 1582 8880 1638 8936
rect 4498 28858 4554 28860
rect 4578 28858 4634 28860
rect 4658 28858 4714 28860
rect 4738 28858 4794 28860
rect 4498 28806 4544 28858
rect 4544 28806 4554 28858
rect 4578 28806 4608 28858
rect 4608 28806 4620 28858
rect 4620 28806 4634 28858
rect 4658 28806 4672 28858
rect 4672 28806 4684 28858
rect 4684 28806 4714 28858
rect 4738 28806 4748 28858
rect 4748 28806 4794 28858
rect 4498 28804 4554 28806
rect 4578 28804 4634 28806
rect 4658 28804 4714 28806
rect 4738 28804 4794 28806
rect 4498 27770 4554 27772
rect 4578 27770 4634 27772
rect 4658 27770 4714 27772
rect 4738 27770 4794 27772
rect 4498 27718 4544 27770
rect 4544 27718 4554 27770
rect 4578 27718 4608 27770
rect 4608 27718 4620 27770
rect 4620 27718 4634 27770
rect 4658 27718 4672 27770
rect 4672 27718 4684 27770
rect 4684 27718 4714 27770
rect 4738 27718 4748 27770
rect 4748 27718 4794 27770
rect 4498 27716 4554 27718
rect 4578 27716 4634 27718
rect 4658 27716 4714 27718
rect 4738 27716 4794 27718
rect 4498 26682 4554 26684
rect 4578 26682 4634 26684
rect 4658 26682 4714 26684
rect 4738 26682 4794 26684
rect 4498 26630 4544 26682
rect 4544 26630 4554 26682
rect 4578 26630 4608 26682
rect 4608 26630 4620 26682
rect 4620 26630 4634 26682
rect 4658 26630 4672 26682
rect 4672 26630 4684 26682
rect 4684 26630 4714 26682
rect 4738 26630 4748 26682
rect 4748 26630 4794 26682
rect 4498 26628 4554 26630
rect 4578 26628 4634 26630
rect 4658 26628 4714 26630
rect 4738 26628 4794 26630
rect 4498 25594 4554 25596
rect 4578 25594 4634 25596
rect 4658 25594 4714 25596
rect 4738 25594 4794 25596
rect 4498 25542 4544 25594
rect 4544 25542 4554 25594
rect 4578 25542 4608 25594
rect 4608 25542 4620 25594
rect 4620 25542 4634 25594
rect 4658 25542 4672 25594
rect 4672 25542 4684 25594
rect 4684 25542 4714 25594
rect 4738 25542 4748 25594
rect 4748 25542 4794 25594
rect 4498 25540 4554 25542
rect 4578 25540 4634 25542
rect 4658 25540 4714 25542
rect 4738 25540 4794 25542
rect 5354 26424 5410 26480
rect 4498 24506 4554 24508
rect 4578 24506 4634 24508
rect 4658 24506 4714 24508
rect 4738 24506 4794 24508
rect 4498 24454 4544 24506
rect 4544 24454 4554 24506
rect 4578 24454 4608 24506
rect 4608 24454 4620 24506
rect 4620 24454 4634 24506
rect 4658 24454 4672 24506
rect 4672 24454 4684 24506
rect 4684 24454 4714 24506
rect 4738 24454 4748 24506
rect 4748 24454 4794 24506
rect 4498 24452 4554 24454
rect 4578 24452 4634 24454
rect 4658 24452 4714 24454
rect 4738 24452 4794 24454
rect 3330 22652 3332 22672
rect 3332 22652 3384 22672
rect 3384 22652 3386 22672
rect 3330 22616 3386 22652
rect 1398 6160 1454 6216
rect 1674 6160 1730 6216
rect 1582 4156 1584 4176
rect 1584 4156 1636 4176
rect 1636 4156 1638 4176
rect 1582 4120 1638 4156
rect 2686 8472 2742 8528
rect 4498 23418 4554 23420
rect 4578 23418 4634 23420
rect 4658 23418 4714 23420
rect 4738 23418 4794 23420
rect 4498 23366 4544 23418
rect 4544 23366 4554 23418
rect 4578 23366 4608 23418
rect 4608 23366 4620 23418
rect 4620 23366 4634 23418
rect 4658 23366 4672 23418
rect 4672 23366 4684 23418
rect 4684 23366 4714 23418
rect 4738 23366 4748 23418
rect 4748 23366 4794 23418
rect 4498 23364 4554 23366
rect 4578 23364 4634 23366
rect 4658 23364 4714 23366
rect 4738 23364 4794 23366
rect 4498 22330 4554 22332
rect 4578 22330 4634 22332
rect 4658 22330 4714 22332
rect 4738 22330 4794 22332
rect 4498 22278 4544 22330
rect 4544 22278 4554 22330
rect 4578 22278 4608 22330
rect 4608 22278 4620 22330
rect 4620 22278 4634 22330
rect 4658 22278 4672 22330
rect 4672 22278 4684 22330
rect 4684 22278 4714 22330
rect 4738 22278 4748 22330
rect 4748 22278 4794 22330
rect 4498 22276 4554 22278
rect 4578 22276 4634 22278
rect 4658 22276 4714 22278
rect 4738 22276 4794 22278
rect 4498 21242 4554 21244
rect 4578 21242 4634 21244
rect 4658 21242 4714 21244
rect 4738 21242 4794 21244
rect 4498 21190 4544 21242
rect 4544 21190 4554 21242
rect 4578 21190 4608 21242
rect 4608 21190 4620 21242
rect 4620 21190 4634 21242
rect 4658 21190 4672 21242
rect 4672 21190 4684 21242
rect 4684 21190 4714 21242
rect 4738 21190 4748 21242
rect 4748 21190 4794 21242
rect 4498 21188 4554 21190
rect 4578 21188 4634 21190
rect 4658 21188 4714 21190
rect 4738 21188 4794 21190
rect 4498 20154 4554 20156
rect 4578 20154 4634 20156
rect 4658 20154 4714 20156
rect 4738 20154 4794 20156
rect 4498 20102 4544 20154
rect 4544 20102 4554 20154
rect 4578 20102 4608 20154
rect 4608 20102 4620 20154
rect 4620 20102 4634 20154
rect 4658 20102 4672 20154
rect 4672 20102 4684 20154
rect 4684 20102 4714 20154
rect 4738 20102 4748 20154
rect 4748 20102 4794 20154
rect 4498 20100 4554 20102
rect 4578 20100 4634 20102
rect 4658 20100 4714 20102
rect 4738 20100 4794 20102
rect 4498 19066 4554 19068
rect 4578 19066 4634 19068
rect 4658 19066 4714 19068
rect 4738 19066 4794 19068
rect 4498 19014 4544 19066
rect 4544 19014 4554 19066
rect 4578 19014 4608 19066
rect 4608 19014 4620 19066
rect 4620 19014 4634 19066
rect 4658 19014 4672 19066
rect 4672 19014 4684 19066
rect 4684 19014 4714 19066
rect 4738 19014 4748 19066
rect 4748 19014 4794 19066
rect 4498 19012 4554 19014
rect 4578 19012 4634 19014
rect 4658 19012 4714 19014
rect 4738 19012 4794 19014
rect 4498 17978 4554 17980
rect 4578 17978 4634 17980
rect 4658 17978 4714 17980
rect 4738 17978 4794 17980
rect 4498 17926 4544 17978
rect 4544 17926 4554 17978
rect 4578 17926 4608 17978
rect 4608 17926 4620 17978
rect 4620 17926 4634 17978
rect 4658 17926 4672 17978
rect 4672 17926 4684 17978
rect 4684 17926 4714 17978
rect 4738 17926 4748 17978
rect 4748 17926 4794 17978
rect 4498 17924 4554 17926
rect 4578 17924 4634 17926
rect 4658 17924 4714 17926
rect 4738 17924 4794 17926
rect 4498 16890 4554 16892
rect 4578 16890 4634 16892
rect 4658 16890 4714 16892
rect 4738 16890 4794 16892
rect 4498 16838 4544 16890
rect 4544 16838 4554 16890
rect 4578 16838 4608 16890
rect 4608 16838 4620 16890
rect 4620 16838 4634 16890
rect 4658 16838 4672 16890
rect 4672 16838 4684 16890
rect 4684 16838 4714 16890
rect 4738 16838 4748 16890
rect 4748 16838 4794 16890
rect 4498 16836 4554 16838
rect 4578 16836 4634 16838
rect 4658 16836 4714 16838
rect 4738 16836 4794 16838
rect 4498 15802 4554 15804
rect 4578 15802 4634 15804
rect 4658 15802 4714 15804
rect 4738 15802 4794 15804
rect 4498 15750 4544 15802
rect 4544 15750 4554 15802
rect 4578 15750 4608 15802
rect 4608 15750 4620 15802
rect 4620 15750 4634 15802
rect 4658 15750 4672 15802
rect 4672 15750 4684 15802
rect 4684 15750 4714 15802
rect 4738 15750 4748 15802
rect 4748 15750 4794 15802
rect 4498 15748 4554 15750
rect 4578 15748 4634 15750
rect 4658 15748 4714 15750
rect 4738 15748 4794 15750
rect 4498 14714 4554 14716
rect 4578 14714 4634 14716
rect 4658 14714 4714 14716
rect 4738 14714 4794 14716
rect 4498 14662 4544 14714
rect 4544 14662 4554 14714
rect 4578 14662 4608 14714
rect 4608 14662 4620 14714
rect 4620 14662 4634 14714
rect 4658 14662 4672 14714
rect 4672 14662 4684 14714
rect 4684 14662 4714 14714
rect 4738 14662 4748 14714
rect 4748 14662 4794 14714
rect 4498 14660 4554 14662
rect 4578 14660 4634 14662
rect 4658 14660 4714 14662
rect 4738 14660 4794 14662
rect 4498 13626 4554 13628
rect 4578 13626 4634 13628
rect 4658 13626 4714 13628
rect 4738 13626 4794 13628
rect 4498 13574 4544 13626
rect 4544 13574 4554 13626
rect 4578 13574 4608 13626
rect 4608 13574 4620 13626
rect 4620 13574 4634 13626
rect 4658 13574 4672 13626
rect 4672 13574 4684 13626
rect 4684 13574 4714 13626
rect 4738 13574 4748 13626
rect 4748 13574 4794 13626
rect 4498 13572 4554 13574
rect 4578 13572 4634 13574
rect 4658 13572 4714 13574
rect 4738 13572 4794 13574
rect 4498 12538 4554 12540
rect 4578 12538 4634 12540
rect 4658 12538 4714 12540
rect 4738 12538 4794 12540
rect 4498 12486 4544 12538
rect 4544 12486 4554 12538
rect 4578 12486 4608 12538
rect 4608 12486 4620 12538
rect 4620 12486 4634 12538
rect 4658 12486 4672 12538
rect 4672 12486 4684 12538
rect 4684 12486 4714 12538
rect 4738 12486 4748 12538
rect 4748 12486 4794 12538
rect 4498 12484 4554 12486
rect 4578 12484 4634 12486
rect 4658 12484 4714 12486
rect 4738 12484 4794 12486
rect 3422 7248 3478 7304
rect 2962 4020 2964 4040
rect 2964 4020 3016 4040
rect 3016 4020 3018 4040
rect 2962 3984 3018 4020
rect 4498 11450 4554 11452
rect 4578 11450 4634 11452
rect 4658 11450 4714 11452
rect 4738 11450 4794 11452
rect 4498 11398 4544 11450
rect 4544 11398 4554 11450
rect 4578 11398 4608 11450
rect 4608 11398 4620 11450
rect 4620 11398 4634 11450
rect 4658 11398 4672 11450
rect 4672 11398 4684 11450
rect 4684 11398 4714 11450
rect 4738 11398 4748 11450
rect 4748 11398 4794 11450
rect 4498 11396 4554 11398
rect 4578 11396 4634 11398
rect 4658 11396 4714 11398
rect 4738 11396 4794 11398
rect 8040 29402 8096 29404
rect 8120 29402 8176 29404
rect 8200 29402 8256 29404
rect 8280 29402 8336 29404
rect 8040 29350 8086 29402
rect 8086 29350 8096 29402
rect 8120 29350 8150 29402
rect 8150 29350 8162 29402
rect 8162 29350 8176 29402
rect 8200 29350 8214 29402
rect 8214 29350 8226 29402
rect 8226 29350 8256 29402
rect 8280 29350 8290 29402
rect 8290 29350 8336 29402
rect 8040 29348 8096 29350
rect 8120 29348 8176 29350
rect 8200 29348 8256 29350
rect 8280 29348 8336 29350
rect 8040 28314 8096 28316
rect 8120 28314 8176 28316
rect 8200 28314 8256 28316
rect 8280 28314 8336 28316
rect 8040 28262 8086 28314
rect 8086 28262 8096 28314
rect 8120 28262 8150 28314
rect 8150 28262 8162 28314
rect 8162 28262 8176 28314
rect 8200 28262 8214 28314
rect 8214 28262 8226 28314
rect 8226 28262 8256 28314
rect 8280 28262 8290 28314
rect 8290 28262 8336 28314
rect 8040 28260 8096 28262
rect 8120 28260 8176 28262
rect 8200 28260 8256 28262
rect 8280 28260 8336 28262
rect 15124 30490 15180 30492
rect 15204 30490 15260 30492
rect 15284 30490 15340 30492
rect 15364 30490 15420 30492
rect 15124 30438 15170 30490
rect 15170 30438 15180 30490
rect 15204 30438 15234 30490
rect 15234 30438 15246 30490
rect 15246 30438 15260 30490
rect 15284 30438 15298 30490
rect 15298 30438 15310 30490
rect 15310 30438 15340 30490
rect 15364 30438 15374 30490
rect 15374 30438 15420 30490
rect 15124 30436 15180 30438
rect 15204 30436 15260 30438
rect 15284 30436 15340 30438
rect 15364 30436 15420 30438
rect 22208 30490 22264 30492
rect 22288 30490 22344 30492
rect 22368 30490 22424 30492
rect 22448 30490 22504 30492
rect 22208 30438 22254 30490
rect 22254 30438 22264 30490
rect 22288 30438 22318 30490
rect 22318 30438 22330 30490
rect 22330 30438 22344 30490
rect 22368 30438 22382 30490
rect 22382 30438 22394 30490
rect 22394 30438 22424 30490
rect 22448 30438 22458 30490
rect 22458 30438 22504 30490
rect 22208 30436 22264 30438
rect 22288 30436 22344 30438
rect 22368 30436 22424 30438
rect 22448 30436 22504 30438
rect 11582 29946 11638 29948
rect 11662 29946 11718 29948
rect 11742 29946 11798 29948
rect 11822 29946 11878 29948
rect 11582 29894 11628 29946
rect 11628 29894 11638 29946
rect 11662 29894 11692 29946
rect 11692 29894 11704 29946
rect 11704 29894 11718 29946
rect 11742 29894 11756 29946
rect 11756 29894 11768 29946
rect 11768 29894 11798 29946
rect 11822 29894 11832 29946
rect 11832 29894 11878 29946
rect 11582 29892 11638 29894
rect 11662 29892 11718 29894
rect 11742 29892 11798 29894
rect 11822 29892 11878 29894
rect 8040 27226 8096 27228
rect 8120 27226 8176 27228
rect 8200 27226 8256 27228
rect 8280 27226 8336 27228
rect 8040 27174 8086 27226
rect 8086 27174 8096 27226
rect 8120 27174 8150 27226
rect 8150 27174 8162 27226
rect 8162 27174 8176 27226
rect 8200 27174 8214 27226
rect 8214 27174 8226 27226
rect 8226 27174 8256 27226
rect 8280 27174 8290 27226
rect 8290 27174 8336 27226
rect 8040 27172 8096 27174
rect 8120 27172 8176 27174
rect 8200 27172 8256 27174
rect 8280 27172 8336 27174
rect 8298 26288 8354 26344
rect 8040 26138 8096 26140
rect 8120 26138 8176 26140
rect 8200 26138 8256 26140
rect 8280 26138 8336 26140
rect 8040 26086 8086 26138
rect 8086 26086 8096 26138
rect 8120 26086 8150 26138
rect 8150 26086 8162 26138
rect 8162 26086 8176 26138
rect 8200 26086 8214 26138
rect 8214 26086 8226 26138
rect 8226 26086 8256 26138
rect 8280 26086 8290 26138
rect 8290 26086 8336 26138
rect 8040 26084 8096 26086
rect 8120 26084 8176 26086
rect 8200 26084 8256 26086
rect 8280 26084 8336 26086
rect 8040 25050 8096 25052
rect 8120 25050 8176 25052
rect 8200 25050 8256 25052
rect 8280 25050 8336 25052
rect 8040 24998 8086 25050
rect 8086 24998 8096 25050
rect 8120 24998 8150 25050
rect 8150 24998 8162 25050
rect 8162 24998 8176 25050
rect 8200 24998 8214 25050
rect 8214 24998 8226 25050
rect 8226 24998 8256 25050
rect 8280 24998 8290 25050
rect 8290 24998 8336 25050
rect 8040 24996 8096 24998
rect 8120 24996 8176 24998
rect 8200 24996 8256 24998
rect 8280 24996 8336 24998
rect 8040 23962 8096 23964
rect 8120 23962 8176 23964
rect 8200 23962 8256 23964
rect 8280 23962 8336 23964
rect 8040 23910 8086 23962
rect 8086 23910 8096 23962
rect 8120 23910 8150 23962
rect 8150 23910 8162 23962
rect 8162 23910 8176 23962
rect 8200 23910 8214 23962
rect 8214 23910 8226 23962
rect 8226 23910 8256 23962
rect 8280 23910 8290 23962
rect 8290 23910 8336 23962
rect 8040 23908 8096 23910
rect 8120 23908 8176 23910
rect 8200 23908 8256 23910
rect 8280 23908 8336 23910
rect 8040 22874 8096 22876
rect 8120 22874 8176 22876
rect 8200 22874 8256 22876
rect 8280 22874 8336 22876
rect 8040 22822 8086 22874
rect 8086 22822 8096 22874
rect 8120 22822 8150 22874
rect 8150 22822 8162 22874
rect 8162 22822 8176 22874
rect 8200 22822 8214 22874
rect 8214 22822 8226 22874
rect 8226 22822 8256 22874
rect 8280 22822 8290 22874
rect 8290 22822 8336 22874
rect 8040 22820 8096 22822
rect 8120 22820 8176 22822
rect 8200 22820 8256 22822
rect 8280 22820 8336 22822
rect 8040 21786 8096 21788
rect 8120 21786 8176 21788
rect 8200 21786 8256 21788
rect 8280 21786 8336 21788
rect 8040 21734 8086 21786
rect 8086 21734 8096 21786
rect 8120 21734 8150 21786
rect 8150 21734 8162 21786
rect 8162 21734 8176 21786
rect 8200 21734 8214 21786
rect 8214 21734 8226 21786
rect 8226 21734 8256 21786
rect 8280 21734 8290 21786
rect 8290 21734 8336 21786
rect 8040 21732 8096 21734
rect 8120 21732 8176 21734
rect 8200 21732 8256 21734
rect 8280 21732 8336 21734
rect 8040 20698 8096 20700
rect 8120 20698 8176 20700
rect 8200 20698 8256 20700
rect 8280 20698 8336 20700
rect 8040 20646 8086 20698
rect 8086 20646 8096 20698
rect 8120 20646 8150 20698
rect 8150 20646 8162 20698
rect 8162 20646 8176 20698
rect 8200 20646 8214 20698
rect 8214 20646 8226 20698
rect 8226 20646 8256 20698
rect 8280 20646 8290 20698
rect 8290 20646 8336 20698
rect 8040 20644 8096 20646
rect 8120 20644 8176 20646
rect 8200 20644 8256 20646
rect 8280 20644 8336 20646
rect 4498 10362 4554 10364
rect 4578 10362 4634 10364
rect 4658 10362 4714 10364
rect 4738 10362 4794 10364
rect 4498 10310 4544 10362
rect 4544 10310 4554 10362
rect 4578 10310 4608 10362
rect 4608 10310 4620 10362
rect 4620 10310 4634 10362
rect 4658 10310 4672 10362
rect 4672 10310 4684 10362
rect 4684 10310 4714 10362
rect 4738 10310 4748 10362
rect 4748 10310 4794 10362
rect 4498 10308 4554 10310
rect 4578 10308 4634 10310
rect 4658 10308 4714 10310
rect 4738 10308 4794 10310
rect 4498 9274 4554 9276
rect 4578 9274 4634 9276
rect 4658 9274 4714 9276
rect 4738 9274 4794 9276
rect 4498 9222 4544 9274
rect 4544 9222 4554 9274
rect 4578 9222 4608 9274
rect 4608 9222 4620 9274
rect 4620 9222 4634 9274
rect 4658 9222 4672 9274
rect 4672 9222 4684 9274
rect 4684 9222 4714 9274
rect 4738 9222 4748 9274
rect 4748 9222 4794 9274
rect 4498 9220 4554 9222
rect 4578 9220 4634 9222
rect 4658 9220 4714 9222
rect 4738 9220 4794 9222
rect 4498 8186 4554 8188
rect 4578 8186 4634 8188
rect 4658 8186 4714 8188
rect 4738 8186 4794 8188
rect 4498 8134 4544 8186
rect 4544 8134 4554 8186
rect 4578 8134 4608 8186
rect 4608 8134 4620 8186
rect 4620 8134 4634 8186
rect 4658 8134 4672 8186
rect 4672 8134 4684 8186
rect 4684 8134 4714 8186
rect 4738 8134 4748 8186
rect 4748 8134 4794 8186
rect 4498 8132 4554 8134
rect 4578 8132 4634 8134
rect 4658 8132 4714 8134
rect 4738 8132 4794 8134
rect 4498 7098 4554 7100
rect 4578 7098 4634 7100
rect 4658 7098 4714 7100
rect 4738 7098 4794 7100
rect 4498 7046 4544 7098
rect 4544 7046 4554 7098
rect 4578 7046 4608 7098
rect 4608 7046 4620 7098
rect 4620 7046 4634 7098
rect 4658 7046 4672 7098
rect 4672 7046 4684 7098
rect 4684 7046 4714 7098
rect 4738 7046 4748 7098
rect 4748 7046 4794 7098
rect 4498 7044 4554 7046
rect 4578 7044 4634 7046
rect 4658 7044 4714 7046
rect 4738 7044 4794 7046
rect 4498 6010 4554 6012
rect 4578 6010 4634 6012
rect 4658 6010 4714 6012
rect 4738 6010 4794 6012
rect 4498 5958 4544 6010
rect 4544 5958 4554 6010
rect 4578 5958 4608 6010
rect 4608 5958 4620 6010
rect 4620 5958 4634 6010
rect 4658 5958 4672 6010
rect 4672 5958 4684 6010
rect 4684 5958 4714 6010
rect 4738 5958 4748 6010
rect 4748 5958 4794 6010
rect 4498 5956 4554 5958
rect 4578 5956 4634 5958
rect 4658 5956 4714 5958
rect 4738 5956 4794 5958
rect 7654 15972 7710 16008
rect 8040 19610 8096 19612
rect 8120 19610 8176 19612
rect 8200 19610 8256 19612
rect 8280 19610 8336 19612
rect 8040 19558 8086 19610
rect 8086 19558 8096 19610
rect 8120 19558 8150 19610
rect 8150 19558 8162 19610
rect 8162 19558 8176 19610
rect 8200 19558 8214 19610
rect 8214 19558 8226 19610
rect 8226 19558 8256 19610
rect 8280 19558 8290 19610
rect 8290 19558 8336 19610
rect 8040 19556 8096 19558
rect 8120 19556 8176 19558
rect 8200 19556 8256 19558
rect 8280 19556 8336 19558
rect 8040 18522 8096 18524
rect 8120 18522 8176 18524
rect 8200 18522 8256 18524
rect 8280 18522 8336 18524
rect 8040 18470 8086 18522
rect 8086 18470 8096 18522
rect 8120 18470 8150 18522
rect 8150 18470 8162 18522
rect 8162 18470 8176 18522
rect 8200 18470 8214 18522
rect 8214 18470 8226 18522
rect 8226 18470 8256 18522
rect 8280 18470 8290 18522
rect 8290 18470 8336 18522
rect 8040 18468 8096 18470
rect 8120 18468 8176 18470
rect 8200 18468 8256 18470
rect 8280 18468 8336 18470
rect 8040 17434 8096 17436
rect 8120 17434 8176 17436
rect 8200 17434 8256 17436
rect 8280 17434 8336 17436
rect 8040 17382 8086 17434
rect 8086 17382 8096 17434
rect 8120 17382 8150 17434
rect 8150 17382 8162 17434
rect 8162 17382 8176 17434
rect 8200 17382 8214 17434
rect 8214 17382 8226 17434
rect 8226 17382 8256 17434
rect 8280 17382 8290 17434
rect 8290 17382 8336 17434
rect 8040 17380 8096 17382
rect 8120 17380 8176 17382
rect 8200 17380 8256 17382
rect 8280 17380 8336 17382
rect 8040 16346 8096 16348
rect 8120 16346 8176 16348
rect 8200 16346 8256 16348
rect 8280 16346 8336 16348
rect 8040 16294 8086 16346
rect 8086 16294 8096 16346
rect 8120 16294 8150 16346
rect 8150 16294 8162 16346
rect 8162 16294 8176 16346
rect 8200 16294 8214 16346
rect 8214 16294 8226 16346
rect 8226 16294 8256 16346
rect 8280 16294 8290 16346
rect 8290 16294 8336 16346
rect 8040 16292 8096 16294
rect 8120 16292 8176 16294
rect 8200 16292 8256 16294
rect 8280 16292 8336 16294
rect 7654 15952 7656 15972
rect 7656 15952 7708 15972
rect 7708 15952 7710 15972
rect 7838 15952 7894 16008
rect 8040 15258 8096 15260
rect 8120 15258 8176 15260
rect 8200 15258 8256 15260
rect 8280 15258 8336 15260
rect 8040 15206 8086 15258
rect 8086 15206 8096 15258
rect 8120 15206 8150 15258
rect 8150 15206 8162 15258
rect 8162 15206 8176 15258
rect 8200 15206 8214 15258
rect 8214 15206 8226 15258
rect 8226 15206 8256 15258
rect 8280 15206 8290 15258
rect 8290 15206 8336 15258
rect 8040 15204 8096 15206
rect 8120 15204 8176 15206
rect 8200 15204 8256 15206
rect 8280 15204 8336 15206
rect 7562 13948 7564 13968
rect 7564 13948 7616 13968
rect 7616 13948 7618 13968
rect 7562 13912 7618 13948
rect 8040 14170 8096 14172
rect 8120 14170 8176 14172
rect 8200 14170 8256 14172
rect 8280 14170 8336 14172
rect 8040 14118 8086 14170
rect 8086 14118 8096 14170
rect 8120 14118 8150 14170
rect 8150 14118 8162 14170
rect 8162 14118 8176 14170
rect 8200 14118 8214 14170
rect 8214 14118 8226 14170
rect 8226 14118 8256 14170
rect 8280 14118 8290 14170
rect 8290 14118 8336 14170
rect 8040 14116 8096 14118
rect 8120 14116 8176 14118
rect 8200 14116 8256 14118
rect 8280 14116 8336 14118
rect 8040 13082 8096 13084
rect 8120 13082 8176 13084
rect 8200 13082 8256 13084
rect 8280 13082 8336 13084
rect 8040 13030 8086 13082
rect 8086 13030 8096 13082
rect 8120 13030 8150 13082
rect 8150 13030 8162 13082
rect 8162 13030 8176 13082
rect 8200 13030 8214 13082
rect 8214 13030 8226 13082
rect 8226 13030 8256 13082
rect 8280 13030 8290 13082
rect 8290 13030 8336 13082
rect 8040 13028 8096 13030
rect 8120 13028 8176 13030
rect 8200 13028 8256 13030
rect 8280 13028 8336 13030
rect 10414 25900 10470 25936
rect 10414 25880 10416 25900
rect 10416 25880 10468 25900
rect 10468 25880 10470 25900
rect 8040 11994 8096 11996
rect 8120 11994 8176 11996
rect 8200 11994 8256 11996
rect 8280 11994 8336 11996
rect 8040 11942 8086 11994
rect 8086 11942 8096 11994
rect 8120 11942 8150 11994
rect 8150 11942 8162 11994
rect 8162 11942 8176 11994
rect 8200 11942 8214 11994
rect 8214 11942 8226 11994
rect 8226 11942 8256 11994
rect 8280 11942 8290 11994
rect 8290 11942 8336 11994
rect 8040 11940 8096 11942
rect 8120 11940 8176 11942
rect 8200 11940 8256 11942
rect 8280 11940 8336 11942
rect 8040 10906 8096 10908
rect 8120 10906 8176 10908
rect 8200 10906 8256 10908
rect 8280 10906 8336 10908
rect 8040 10854 8086 10906
rect 8086 10854 8096 10906
rect 8120 10854 8150 10906
rect 8150 10854 8162 10906
rect 8162 10854 8176 10906
rect 8200 10854 8214 10906
rect 8214 10854 8226 10906
rect 8226 10854 8256 10906
rect 8280 10854 8290 10906
rect 8290 10854 8336 10906
rect 8040 10852 8096 10854
rect 8120 10852 8176 10854
rect 8200 10852 8256 10854
rect 8280 10852 8336 10854
rect 7286 9596 7288 9616
rect 7288 9596 7340 9616
rect 7340 9596 7342 9616
rect 7286 9560 7342 9596
rect 8040 9818 8096 9820
rect 8120 9818 8176 9820
rect 8200 9818 8256 9820
rect 8280 9818 8336 9820
rect 8040 9766 8086 9818
rect 8086 9766 8096 9818
rect 8120 9766 8150 9818
rect 8150 9766 8162 9818
rect 8162 9766 8176 9818
rect 8200 9766 8214 9818
rect 8214 9766 8226 9818
rect 8226 9766 8256 9818
rect 8280 9766 8290 9818
rect 8290 9766 8336 9818
rect 8040 9764 8096 9766
rect 8120 9764 8176 9766
rect 8200 9764 8256 9766
rect 8280 9764 8336 9766
rect 7930 8880 7986 8936
rect 8040 8730 8096 8732
rect 8120 8730 8176 8732
rect 8200 8730 8256 8732
rect 8280 8730 8336 8732
rect 8040 8678 8086 8730
rect 8086 8678 8096 8730
rect 8120 8678 8150 8730
rect 8150 8678 8162 8730
rect 8162 8678 8176 8730
rect 8200 8678 8214 8730
rect 8214 8678 8226 8730
rect 8226 8678 8256 8730
rect 8280 8678 8290 8730
rect 8290 8678 8336 8730
rect 8040 8676 8096 8678
rect 8120 8676 8176 8678
rect 8200 8676 8256 8678
rect 8280 8676 8336 8678
rect 8040 7642 8096 7644
rect 8120 7642 8176 7644
rect 8200 7642 8256 7644
rect 8280 7642 8336 7644
rect 8040 7590 8086 7642
rect 8086 7590 8096 7642
rect 8120 7590 8150 7642
rect 8150 7590 8162 7642
rect 8162 7590 8176 7642
rect 8200 7590 8214 7642
rect 8214 7590 8226 7642
rect 8226 7590 8256 7642
rect 8280 7590 8290 7642
rect 8290 7590 8336 7642
rect 8040 7588 8096 7590
rect 8120 7588 8176 7590
rect 8200 7588 8256 7590
rect 8280 7588 8336 7590
rect 8040 6554 8096 6556
rect 8120 6554 8176 6556
rect 8200 6554 8256 6556
rect 8280 6554 8336 6556
rect 8040 6502 8086 6554
rect 8086 6502 8096 6554
rect 8120 6502 8150 6554
rect 8150 6502 8162 6554
rect 8162 6502 8176 6554
rect 8200 6502 8214 6554
rect 8214 6502 8226 6554
rect 8226 6502 8256 6554
rect 8280 6502 8290 6554
rect 8290 6502 8336 6554
rect 8040 6500 8096 6502
rect 8120 6500 8176 6502
rect 8200 6500 8256 6502
rect 8280 6500 8336 6502
rect 4498 4922 4554 4924
rect 4578 4922 4634 4924
rect 4658 4922 4714 4924
rect 4738 4922 4794 4924
rect 4498 4870 4544 4922
rect 4544 4870 4554 4922
rect 4578 4870 4608 4922
rect 4608 4870 4620 4922
rect 4620 4870 4634 4922
rect 4658 4870 4672 4922
rect 4672 4870 4684 4922
rect 4684 4870 4714 4922
rect 4738 4870 4748 4922
rect 4748 4870 4794 4922
rect 4498 4868 4554 4870
rect 4578 4868 4634 4870
rect 4658 4868 4714 4870
rect 4738 4868 4794 4870
rect 4498 3834 4554 3836
rect 4578 3834 4634 3836
rect 4658 3834 4714 3836
rect 4738 3834 4794 3836
rect 4498 3782 4544 3834
rect 4544 3782 4554 3834
rect 4578 3782 4608 3834
rect 4608 3782 4620 3834
rect 4620 3782 4634 3834
rect 4658 3782 4672 3834
rect 4672 3782 4684 3834
rect 4684 3782 4714 3834
rect 4738 3782 4748 3834
rect 4748 3782 4794 3834
rect 4498 3780 4554 3782
rect 4578 3780 4634 3782
rect 4658 3780 4714 3782
rect 4738 3780 4794 3782
rect 4498 2746 4554 2748
rect 4578 2746 4634 2748
rect 4658 2746 4714 2748
rect 4738 2746 4794 2748
rect 4498 2694 4544 2746
rect 4544 2694 4554 2746
rect 4578 2694 4608 2746
rect 4608 2694 4620 2746
rect 4620 2694 4634 2746
rect 4658 2694 4672 2746
rect 4672 2694 4684 2746
rect 4684 2694 4714 2746
rect 4738 2694 4748 2746
rect 4748 2694 4794 2746
rect 4498 2692 4554 2694
rect 4578 2692 4634 2694
rect 4658 2692 4714 2694
rect 4738 2692 4794 2694
rect 8040 5466 8096 5468
rect 8120 5466 8176 5468
rect 8200 5466 8256 5468
rect 8280 5466 8336 5468
rect 8040 5414 8086 5466
rect 8086 5414 8096 5466
rect 8120 5414 8150 5466
rect 8150 5414 8162 5466
rect 8162 5414 8176 5466
rect 8200 5414 8214 5466
rect 8214 5414 8226 5466
rect 8226 5414 8256 5466
rect 8280 5414 8290 5466
rect 8290 5414 8336 5466
rect 8040 5412 8096 5414
rect 8120 5412 8176 5414
rect 8200 5412 8256 5414
rect 8280 5412 8336 5414
rect 8040 4378 8096 4380
rect 8120 4378 8176 4380
rect 8200 4378 8256 4380
rect 8280 4378 8336 4380
rect 8040 4326 8086 4378
rect 8086 4326 8096 4378
rect 8120 4326 8150 4378
rect 8150 4326 8162 4378
rect 8162 4326 8176 4378
rect 8200 4326 8214 4378
rect 8214 4326 8226 4378
rect 8226 4326 8256 4378
rect 8280 4326 8290 4378
rect 8290 4326 8336 4378
rect 8040 4324 8096 4326
rect 8120 4324 8176 4326
rect 8200 4324 8256 4326
rect 8280 4324 8336 4326
rect 8040 3290 8096 3292
rect 8120 3290 8176 3292
rect 8200 3290 8256 3292
rect 8280 3290 8336 3292
rect 8040 3238 8086 3290
rect 8086 3238 8096 3290
rect 8120 3238 8150 3290
rect 8150 3238 8162 3290
rect 8162 3238 8176 3290
rect 8200 3238 8214 3290
rect 8214 3238 8226 3290
rect 8226 3238 8256 3290
rect 8280 3238 8290 3290
rect 8290 3238 8336 3290
rect 8040 3236 8096 3238
rect 8120 3236 8176 3238
rect 8200 3236 8256 3238
rect 8280 3236 8336 3238
rect 9402 14864 9458 14920
rect 11582 28858 11638 28860
rect 11662 28858 11718 28860
rect 11742 28858 11798 28860
rect 11822 28858 11878 28860
rect 11582 28806 11628 28858
rect 11628 28806 11638 28858
rect 11662 28806 11692 28858
rect 11692 28806 11704 28858
rect 11704 28806 11718 28858
rect 11742 28806 11756 28858
rect 11756 28806 11768 28858
rect 11768 28806 11798 28858
rect 11822 28806 11832 28858
rect 11832 28806 11878 28858
rect 11582 28804 11638 28806
rect 11662 28804 11718 28806
rect 11742 28804 11798 28806
rect 11822 28804 11878 28806
rect 11582 27770 11638 27772
rect 11662 27770 11718 27772
rect 11742 27770 11798 27772
rect 11822 27770 11878 27772
rect 11582 27718 11628 27770
rect 11628 27718 11638 27770
rect 11662 27718 11692 27770
rect 11692 27718 11704 27770
rect 11704 27718 11718 27770
rect 11742 27718 11756 27770
rect 11756 27718 11768 27770
rect 11768 27718 11798 27770
rect 11822 27718 11832 27770
rect 11832 27718 11878 27770
rect 11582 27716 11638 27718
rect 11662 27716 11718 27718
rect 11742 27716 11798 27718
rect 11822 27716 11878 27718
rect 11582 26682 11638 26684
rect 11662 26682 11718 26684
rect 11742 26682 11798 26684
rect 11822 26682 11878 26684
rect 11582 26630 11628 26682
rect 11628 26630 11638 26682
rect 11662 26630 11692 26682
rect 11692 26630 11704 26682
rect 11704 26630 11718 26682
rect 11742 26630 11756 26682
rect 11756 26630 11768 26682
rect 11768 26630 11798 26682
rect 11822 26630 11832 26682
rect 11832 26630 11878 26682
rect 11582 26628 11638 26630
rect 11662 26628 11718 26630
rect 11742 26628 11798 26630
rect 11822 26628 11878 26630
rect 11978 25880 12034 25936
rect 11582 25594 11638 25596
rect 11662 25594 11718 25596
rect 11742 25594 11798 25596
rect 11822 25594 11878 25596
rect 11582 25542 11628 25594
rect 11628 25542 11638 25594
rect 11662 25542 11692 25594
rect 11692 25542 11704 25594
rect 11704 25542 11718 25594
rect 11742 25542 11756 25594
rect 11756 25542 11768 25594
rect 11768 25542 11798 25594
rect 11822 25542 11832 25594
rect 11832 25542 11878 25594
rect 11582 25540 11638 25542
rect 11662 25540 11718 25542
rect 11742 25540 11798 25542
rect 11822 25540 11878 25542
rect 11582 24506 11638 24508
rect 11662 24506 11718 24508
rect 11742 24506 11798 24508
rect 11822 24506 11878 24508
rect 11582 24454 11628 24506
rect 11628 24454 11638 24506
rect 11662 24454 11692 24506
rect 11692 24454 11704 24506
rect 11704 24454 11718 24506
rect 11742 24454 11756 24506
rect 11756 24454 11768 24506
rect 11768 24454 11798 24506
rect 11822 24454 11832 24506
rect 11832 24454 11878 24506
rect 11582 24452 11638 24454
rect 11662 24452 11718 24454
rect 11742 24452 11798 24454
rect 11822 24452 11878 24454
rect 11582 23418 11638 23420
rect 11662 23418 11718 23420
rect 11742 23418 11798 23420
rect 11822 23418 11878 23420
rect 11582 23366 11628 23418
rect 11628 23366 11638 23418
rect 11662 23366 11692 23418
rect 11692 23366 11704 23418
rect 11704 23366 11718 23418
rect 11742 23366 11756 23418
rect 11756 23366 11768 23418
rect 11768 23366 11798 23418
rect 11822 23366 11832 23418
rect 11832 23366 11878 23418
rect 11582 23364 11638 23366
rect 11662 23364 11718 23366
rect 11742 23364 11798 23366
rect 11822 23364 11878 23366
rect 11582 22330 11638 22332
rect 11662 22330 11718 22332
rect 11742 22330 11798 22332
rect 11822 22330 11878 22332
rect 11582 22278 11628 22330
rect 11628 22278 11638 22330
rect 11662 22278 11692 22330
rect 11692 22278 11704 22330
rect 11704 22278 11718 22330
rect 11742 22278 11756 22330
rect 11756 22278 11768 22330
rect 11768 22278 11798 22330
rect 11822 22278 11832 22330
rect 11832 22278 11878 22330
rect 11582 22276 11638 22278
rect 11662 22276 11718 22278
rect 11742 22276 11798 22278
rect 11822 22276 11878 22278
rect 11582 21242 11638 21244
rect 11662 21242 11718 21244
rect 11742 21242 11798 21244
rect 11822 21242 11878 21244
rect 11582 21190 11628 21242
rect 11628 21190 11638 21242
rect 11662 21190 11692 21242
rect 11692 21190 11704 21242
rect 11704 21190 11718 21242
rect 11742 21190 11756 21242
rect 11756 21190 11768 21242
rect 11768 21190 11798 21242
rect 11822 21190 11832 21242
rect 11832 21190 11878 21242
rect 11582 21188 11638 21190
rect 11662 21188 11718 21190
rect 11742 21188 11798 21190
rect 11822 21188 11878 21190
rect 11582 20154 11638 20156
rect 11662 20154 11718 20156
rect 11742 20154 11798 20156
rect 11822 20154 11878 20156
rect 11582 20102 11628 20154
rect 11628 20102 11638 20154
rect 11662 20102 11692 20154
rect 11692 20102 11704 20154
rect 11704 20102 11718 20154
rect 11742 20102 11756 20154
rect 11756 20102 11768 20154
rect 11768 20102 11798 20154
rect 11822 20102 11832 20154
rect 11832 20102 11878 20154
rect 11582 20100 11638 20102
rect 11662 20100 11718 20102
rect 11742 20100 11798 20102
rect 11822 20100 11878 20102
rect 11518 19780 11574 19816
rect 11518 19760 11520 19780
rect 11520 19760 11572 19780
rect 11572 19760 11574 19780
rect 10874 15408 10930 15464
rect 11582 19066 11638 19068
rect 11662 19066 11718 19068
rect 11742 19066 11798 19068
rect 11822 19066 11878 19068
rect 11582 19014 11628 19066
rect 11628 19014 11638 19066
rect 11662 19014 11692 19066
rect 11692 19014 11704 19066
rect 11704 19014 11718 19066
rect 11742 19014 11756 19066
rect 11756 19014 11768 19066
rect 11768 19014 11798 19066
rect 11822 19014 11832 19066
rect 11832 19014 11878 19066
rect 11582 19012 11638 19014
rect 11662 19012 11718 19014
rect 11742 19012 11798 19014
rect 11822 19012 11878 19014
rect 11582 17978 11638 17980
rect 11662 17978 11718 17980
rect 11742 17978 11798 17980
rect 11822 17978 11878 17980
rect 11582 17926 11628 17978
rect 11628 17926 11638 17978
rect 11662 17926 11692 17978
rect 11692 17926 11704 17978
rect 11704 17926 11718 17978
rect 11742 17926 11756 17978
rect 11756 17926 11768 17978
rect 11768 17926 11798 17978
rect 11822 17926 11832 17978
rect 11832 17926 11878 17978
rect 11582 17924 11638 17926
rect 11662 17924 11718 17926
rect 11742 17924 11798 17926
rect 11822 17924 11878 17926
rect 11582 16890 11638 16892
rect 11662 16890 11718 16892
rect 11742 16890 11798 16892
rect 11822 16890 11878 16892
rect 11582 16838 11628 16890
rect 11628 16838 11638 16890
rect 11662 16838 11692 16890
rect 11692 16838 11704 16890
rect 11704 16838 11718 16890
rect 11742 16838 11756 16890
rect 11756 16838 11768 16890
rect 11768 16838 11798 16890
rect 11822 16838 11832 16890
rect 11832 16838 11878 16890
rect 11582 16836 11638 16838
rect 11662 16836 11718 16838
rect 11742 16836 11798 16838
rect 11822 16836 11878 16838
rect 11886 16532 11888 16552
rect 11888 16532 11940 16552
rect 11940 16532 11942 16552
rect 11886 16496 11942 16532
rect 11582 15802 11638 15804
rect 11662 15802 11718 15804
rect 11742 15802 11798 15804
rect 11822 15802 11878 15804
rect 11582 15750 11628 15802
rect 11628 15750 11638 15802
rect 11662 15750 11692 15802
rect 11692 15750 11704 15802
rect 11704 15750 11718 15802
rect 11742 15750 11756 15802
rect 11756 15750 11768 15802
rect 11768 15750 11798 15802
rect 11822 15750 11832 15802
rect 11832 15750 11878 15802
rect 11582 15748 11638 15750
rect 11662 15748 11718 15750
rect 11742 15748 11798 15750
rect 11822 15748 11878 15750
rect 11334 12280 11390 12336
rect 11242 9560 11298 9616
rect 11582 14714 11638 14716
rect 11662 14714 11718 14716
rect 11742 14714 11798 14716
rect 11822 14714 11878 14716
rect 11582 14662 11628 14714
rect 11628 14662 11638 14714
rect 11662 14662 11692 14714
rect 11692 14662 11704 14714
rect 11704 14662 11718 14714
rect 11742 14662 11756 14714
rect 11756 14662 11768 14714
rect 11768 14662 11798 14714
rect 11822 14662 11832 14714
rect 11832 14662 11878 14714
rect 11582 14660 11638 14662
rect 11662 14660 11718 14662
rect 11742 14660 11798 14662
rect 11822 14660 11878 14662
rect 11610 14456 11666 14512
rect 11582 13626 11638 13628
rect 11662 13626 11718 13628
rect 11742 13626 11798 13628
rect 11822 13626 11878 13628
rect 11582 13574 11628 13626
rect 11628 13574 11638 13626
rect 11662 13574 11692 13626
rect 11692 13574 11704 13626
rect 11704 13574 11718 13626
rect 11742 13574 11756 13626
rect 11756 13574 11768 13626
rect 11768 13574 11798 13626
rect 11822 13574 11832 13626
rect 11832 13574 11878 13626
rect 11582 13572 11638 13574
rect 11662 13572 11718 13574
rect 11742 13572 11798 13574
rect 11822 13572 11878 13574
rect 13358 16632 13414 16688
rect 11582 12538 11638 12540
rect 11662 12538 11718 12540
rect 11742 12538 11798 12540
rect 11822 12538 11878 12540
rect 11582 12486 11628 12538
rect 11628 12486 11638 12538
rect 11662 12486 11692 12538
rect 11692 12486 11704 12538
rect 11704 12486 11718 12538
rect 11742 12486 11756 12538
rect 11756 12486 11768 12538
rect 11768 12486 11798 12538
rect 11822 12486 11832 12538
rect 11832 12486 11878 12538
rect 11582 12484 11638 12486
rect 11662 12484 11718 12486
rect 11742 12484 11798 12486
rect 11822 12484 11878 12486
rect 11582 11450 11638 11452
rect 11662 11450 11718 11452
rect 11742 11450 11798 11452
rect 11822 11450 11878 11452
rect 11582 11398 11628 11450
rect 11628 11398 11638 11450
rect 11662 11398 11692 11450
rect 11692 11398 11704 11450
rect 11704 11398 11718 11450
rect 11742 11398 11756 11450
rect 11756 11398 11768 11450
rect 11768 11398 11798 11450
rect 11822 11398 11832 11450
rect 11832 11398 11878 11450
rect 11582 11396 11638 11398
rect 11662 11396 11718 11398
rect 11742 11396 11798 11398
rect 11822 11396 11878 11398
rect 11582 10362 11638 10364
rect 11662 10362 11718 10364
rect 11742 10362 11798 10364
rect 11822 10362 11878 10364
rect 11582 10310 11628 10362
rect 11628 10310 11638 10362
rect 11662 10310 11692 10362
rect 11692 10310 11704 10362
rect 11704 10310 11718 10362
rect 11742 10310 11756 10362
rect 11756 10310 11768 10362
rect 11768 10310 11798 10362
rect 11822 10310 11832 10362
rect 11832 10310 11878 10362
rect 11582 10308 11638 10310
rect 11662 10308 11718 10310
rect 11742 10308 11798 10310
rect 11822 10308 11878 10310
rect 11582 9274 11638 9276
rect 11662 9274 11718 9276
rect 11742 9274 11798 9276
rect 11822 9274 11878 9276
rect 11582 9222 11628 9274
rect 11628 9222 11638 9274
rect 11662 9222 11692 9274
rect 11692 9222 11704 9274
rect 11704 9222 11718 9274
rect 11742 9222 11756 9274
rect 11756 9222 11768 9274
rect 11768 9222 11798 9274
rect 11822 9222 11832 9274
rect 11832 9222 11878 9274
rect 11582 9220 11638 9222
rect 11662 9220 11718 9222
rect 11742 9220 11798 9222
rect 11822 9220 11878 9222
rect 11582 8186 11638 8188
rect 11662 8186 11718 8188
rect 11742 8186 11798 8188
rect 11822 8186 11878 8188
rect 11582 8134 11628 8186
rect 11628 8134 11638 8186
rect 11662 8134 11692 8186
rect 11692 8134 11704 8186
rect 11704 8134 11718 8186
rect 11742 8134 11756 8186
rect 11756 8134 11768 8186
rect 11768 8134 11798 8186
rect 11822 8134 11832 8186
rect 11832 8134 11878 8186
rect 11582 8132 11638 8134
rect 11662 8132 11718 8134
rect 11742 8132 11798 8134
rect 11822 8132 11878 8134
rect 12898 11212 12954 11248
rect 12898 11192 12900 11212
rect 12900 11192 12952 11212
rect 12952 11192 12954 11212
rect 11582 7098 11638 7100
rect 11662 7098 11718 7100
rect 11742 7098 11798 7100
rect 11822 7098 11878 7100
rect 11582 7046 11628 7098
rect 11628 7046 11638 7098
rect 11662 7046 11692 7098
rect 11692 7046 11704 7098
rect 11704 7046 11718 7098
rect 11742 7046 11756 7098
rect 11756 7046 11768 7098
rect 11768 7046 11798 7098
rect 11822 7046 11832 7098
rect 11832 7046 11878 7098
rect 11582 7044 11638 7046
rect 11662 7044 11718 7046
rect 11742 7044 11798 7046
rect 11822 7044 11878 7046
rect 11582 6010 11638 6012
rect 11662 6010 11718 6012
rect 11742 6010 11798 6012
rect 11822 6010 11878 6012
rect 11582 5958 11628 6010
rect 11628 5958 11638 6010
rect 11662 5958 11692 6010
rect 11692 5958 11704 6010
rect 11704 5958 11718 6010
rect 11742 5958 11756 6010
rect 11756 5958 11768 6010
rect 11768 5958 11798 6010
rect 11822 5958 11832 6010
rect 11832 5958 11878 6010
rect 11582 5956 11638 5958
rect 11662 5956 11718 5958
rect 11742 5956 11798 5958
rect 11822 5956 11878 5958
rect 11582 4922 11638 4924
rect 11662 4922 11718 4924
rect 11742 4922 11798 4924
rect 11822 4922 11878 4924
rect 11582 4870 11628 4922
rect 11628 4870 11638 4922
rect 11662 4870 11692 4922
rect 11692 4870 11704 4922
rect 11704 4870 11718 4922
rect 11742 4870 11756 4922
rect 11756 4870 11768 4922
rect 11768 4870 11798 4922
rect 11822 4870 11832 4922
rect 11832 4870 11878 4922
rect 11582 4868 11638 4870
rect 11662 4868 11718 4870
rect 11742 4868 11798 4870
rect 11822 4868 11878 4870
rect 11582 3834 11638 3836
rect 11662 3834 11718 3836
rect 11742 3834 11798 3836
rect 11822 3834 11878 3836
rect 11582 3782 11628 3834
rect 11628 3782 11638 3834
rect 11662 3782 11692 3834
rect 11692 3782 11704 3834
rect 11704 3782 11718 3834
rect 11742 3782 11756 3834
rect 11756 3782 11768 3834
rect 11768 3782 11798 3834
rect 11822 3782 11832 3834
rect 11832 3782 11878 3834
rect 11582 3780 11638 3782
rect 11662 3780 11718 3782
rect 11742 3780 11798 3782
rect 11822 3780 11878 3782
rect 15124 29402 15180 29404
rect 15204 29402 15260 29404
rect 15284 29402 15340 29404
rect 15364 29402 15420 29404
rect 15124 29350 15170 29402
rect 15170 29350 15180 29402
rect 15204 29350 15234 29402
rect 15234 29350 15246 29402
rect 15246 29350 15260 29402
rect 15284 29350 15298 29402
rect 15298 29350 15310 29402
rect 15310 29350 15340 29402
rect 15364 29350 15374 29402
rect 15374 29350 15420 29402
rect 15124 29348 15180 29350
rect 15204 29348 15260 29350
rect 15284 29348 15340 29350
rect 15364 29348 15420 29350
rect 14830 28620 14886 28656
rect 14830 28600 14832 28620
rect 14832 28600 14884 28620
rect 14884 28600 14886 28620
rect 15124 28314 15180 28316
rect 15204 28314 15260 28316
rect 15284 28314 15340 28316
rect 15364 28314 15420 28316
rect 15124 28262 15170 28314
rect 15170 28262 15180 28314
rect 15204 28262 15234 28314
rect 15234 28262 15246 28314
rect 15246 28262 15260 28314
rect 15284 28262 15298 28314
rect 15298 28262 15310 28314
rect 15310 28262 15340 28314
rect 15364 28262 15374 28314
rect 15374 28262 15420 28314
rect 15124 28260 15180 28262
rect 15204 28260 15260 28262
rect 15284 28260 15340 28262
rect 15364 28260 15420 28262
rect 15124 27226 15180 27228
rect 15204 27226 15260 27228
rect 15284 27226 15340 27228
rect 15364 27226 15420 27228
rect 15124 27174 15170 27226
rect 15170 27174 15180 27226
rect 15204 27174 15234 27226
rect 15234 27174 15246 27226
rect 15246 27174 15260 27226
rect 15284 27174 15298 27226
rect 15298 27174 15310 27226
rect 15310 27174 15340 27226
rect 15364 27174 15374 27226
rect 15374 27174 15420 27226
rect 15124 27172 15180 27174
rect 15204 27172 15260 27174
rect 15284 27172 15340 27174
rect 15364 27172 15420 27174
rect 15124 26138 15180 26140
rect 15204 26138 15260 26140
rect 15284 26138 15340 26140
rect 15364 26138 15420 26140
rect 15124 26086 15170 26138
rect 15170 26086 15180 26138
rect 15204 26086 15234 26138
rect 15234 26086 15246 26138
rect 15246 26086 15260 26138
rect 15284 26086 15298 26138
rect 15298 26086 15310 26138
rect 15310 26086 15340 26138
rect 15364 26086 15374 26138
rect 15374 26086 15420 26138
rect 15124 26084 15180 26086
rect 15204 26084 15260 26086
rect 15284 26084 15340 26086
rect 15364 26084 15420 26086
rect 15842 25880 15898 25936
rect 15124 25050 15180 25052
rect 15204 25050 15260 25052
rect 15284 25050 15340 25052
rect 15364 25050 15420 25052
rect 15124 24998 15170 25050
rect 15170 24998 15180 25050
rect 15204 24998 15234 25050
rect 15234 24998 15246 25050
rect 15246 24998 15260 25050
rect 15284 24998 15298 25050
rect 15298 24998 15310 25050
rect 15310 24998 15340 25050
rect 15364 24998 15374 25050
rect 15374 24998 15420 25050
rect 15124 24996 15180 24998
rect 15204 24996 15260 24998
rect 15284 24996 15340 24998
rect 15364 24996 15420 24998
rect 15124 23962 15180 23964
rect 15204 23962 15260 23964
rect 15284 23962 15340 23964
rect 15364 23962 15420 23964
rect 15124 23910 15170 23962
rect 15170 23910 15180 23962
rect 15204 23910 15234 23962
rect 15234 23910 15246 23962
rect 15246 23910 15260 23962
rect 15284 23910 15298 23962
rect 15298 23910 15310 23962
rect 15310 23910 15340 23962
rect 15364 23910 15374 23962
rect 15374 23910 15420 23962
rect 15124 23908 15180 23910
rect 15204 23908 15260 23910
rect 15284 23908 15340 23910
rect 15364 23908 15420 23910
rect 15124 22874 15180 22876
rect 15204 22874 15260 22876
rect 15284 22874 15340 22876
rect 15364 22874 15420 22876
rect 15124 22822 15170 22874
rect 15170 22822 15180 22874
rect 15204 22822 15234 22874
rect 15234 22822 15246 22874
rect 15246 22822 15260 22874
rect 15284 22822 15298 22874
rect 15298 22822 15310 22874
rect 15310 22822 15340 22874
rect 15364 22822 15374 22874
rect 15374 22822 15420 22874
rect 15124 22820 15180 22822
rect 15204 22820 15260 22822
rect 15284 22820 15340 22822
rect 15364 22820 15420 22822
rect 14002 19352 14058 19408
rect 11582 2746 11638 2748
rect 11662 2746 11718 2748
rect 11742 2746 11798 2748
rect 11822 2746 11878 2748
rect 11582 2694 11628 2746
rect 11628 2694 11638 2746
rect 11662 2694 11692 2746
rect 11692 2694 11704 2746
rect 11704 2694 11718 2746
rect 11742 2694 11756 2746
rect 11756 2694 11768 2746
rect 11768 2694 11798 2746
rect 11822 2694 11832 2746
rect 11832 2694 11878 2746
rect 11582 2692 11638 2694
rect 11662 2692 11718 2694
rect 11742 2692 11798 2694
rect 11822 2692 11878 2694
rect 15124 21786 15180 21788
rect 15204 21786 15260 21788
rect 15284 21786 15340 21788
rect 15364 21786 15420 21788
rect 15124 21734 15170 21786
rect 15170 21734 15180 21786
rect 15204 21734 15234 21786
rect 15234 21734 15246 21786
rect 15246 21734 15260 21786
rect 15284 21734 15298 21786
rect 15298 21734 15310 21786
rect 15310 21734 15340 21786
rect 15364 21734 15374 21786
rect 15374 21734 15420 21786
rect 15124 21732 15180 21734
rect 15204 21732 15260 21734
rect 15284 21732 15340 21734
rect 15364 21732 15420 21734
rect 15124 20698 15180 20700
rect 15204 20698 15260 20700
rect 15284 20698 15340 20700
rect 15364 20698 15420 20700
rect 15124 20646 15170 20698
rect 15170 20646 15180 20698
rect 15204 20646 15234 20698
rect 15234 20646 15246 20698
rect 15246 20646 15260 20698
rect 15284 20646 15298 20698
rect 15298 20646 15310 20698
rect 15310 20646 15340 20698
rect 15364 20646 15374 20698
rect 15374 20646 15420 20698
rect 15124 20644 15180 20646
rect 15204 20644 15260 20646
rect 15284 20644 15340 20646
rect 15364 20644 15420 20646
rect 15124 19610 15180 19612
rect 15204 19610 15260 19612
rect 15284 19610 15340 19612
rect 15364 19610 15420 19612
rect 15124 19558 15170 19610
rect 15170 19558 15180 19610
rect 15204 19558 15234 19610
rect 15234 19558 15246 19610
rect 15246 19558 15260 19610
rect 15284 19558 15298 19610
rect 15298 19558 15310 19610
rect 15310 19558 15340 19610
rect 15364 19558 15374 19610
rect 15374 19558 15420 19610
rect 15124 19556 15180 19558
rect 15204 19556 15260 19558
rect 15284 19556 15340 19558
rect 15364 19556 15420 19558
rect 15124 18522 15180 18524
rect 15204 18522 15260 18524
rect 15284 18522 15340 18524
rect 15364 18522 15420 18524
rect 15124 18470 15170 18522
rect 15170 18470 15180 18522
rect 15204 18470 15234 18522
rect 15234 18470 15246 18522
rect 15246 18470 15260 18522
rect 15284 18470 15298 18522
rect 15298 18470 15310 18522
rect 15310 18470 15340 18522
rect 15364 18470 15374 18522
rect 15374 18470 15420 18522
rect 15124 18468 15180 18470
rect 15204 18468 15260 18470
rect 15284 18468 15340 18470
rect 15364 18468 15420 18470
rect 18666 29946 18722 29948
rect 18746 29946 18802 29948
rect 18826 29946 18882 29948
rect 18906 29946 18962 29948
rect 18666 29894 18712 29946
rect 18712 29894 18722 29946
rect 18746 29894 18776 29946
rect 18776 29894 18788 29946
rect 18788 29894 18802 29946
rect 18826 29894 18840 29946
rect 18840 29894 18852 29946
rect 18852 29894 18882 29946
rect 18906 29894 18916 29946
rect 18916 29894 18962 29946
rect 18666 29892 18722 29894
rect 18746 29892 18802 29894
rect 18826 29892 18882 29894
rect 18906 29892 18962 29894
rect 16210 28484 16266 28520
rect 16210 28464 16212 28484
rect 16212 28464 16264 28484
rect 16264 28464 16266 28484
rect 18666 28858 18722 28860
rect 18746 28858 18802 28860
rect 18826 28858 18882 28860
rect 18906 28858 18962 28860
rect 18666 28806 18712 28858
rect 18712 28806 18722 28858
rect 18746 28806 18776 28858
rect 18776 28806 18788 28858
rect 18788 28806 18802 28858
rect 18826 28806 18840 28858
rect 18840 28806 18852 28858
rect 18852 28806 18882 28858
rect 18906 28806 18916 28858
rect 18916 28806 18962 28858
rect 18666 28804 18722 28806
rect 18746 28804 18802 28806
rect 18826 28804 18882 28806
rect 18906 28804 18962 28806
rect 16670 27956 16672 27976
rect 16672 27956 16724 27976
rect 16724 27956 16726 27976
rect 16670 27920 16726 27956
rect 16946 26324 16948 26344
rect 16948 26324 17000 26344
rect 17000 26324 17002 26344
rect 16946 26288 17002 26324
rect 16302 23160 16358 23216
rect 18050 26288 18106 26344
rect 17498 21836 17500 21856
rect 17500 21836 17552 21856
rect 17552 21836 17554 21856
rect 17498 21800 17554 21836
rect 15124 17434 15180 17436
rect 15204 17434 15260 17436
rect 15284 17434 15340 17436
rect 15364 17434 15420 17436
rect 15124 17382 15170 17434
rect 15170 17382 15180 17434
rect 15204 17382 15234 17434
rect 15234 17382 15246 17434
rect 15246 17382 15260 17434
rect 15284 17382 15298 17434
rect 15298 17382 15310 17434
rect 15310 17382 15340 17434
rect 15364 17382 15374 17434
rect 15374 17382 15420 17434
rect 15124 17380 15180 17382
rect 15204 17380 15260 17382
rect 15284 17380 15340 17382
rect 15364 17380 15420 17382
rect 15124 16346 15180 16348
rect 15204 16346 15260 16348
rect 15284 16346 15340 16348
rect 15364 16346 15420 16348
rect 15124 16294 15170 16346
rect 15170 16294 15180 16346
rect 15204 16294 15234 16346
rect 15234 16294 15246 16346
rect 15246 16294 15260 16346
rect 15284 16294 15298 16346
rect 15298 16294 15310 16346
rect 15310 16294 15340 16346
rect 15364 16294 15374 16346
rect 15374 16294 15420 16346
rect 15124 16292 15180 16294
rect 15204 16292 15260 16294
rect 15284 16292 15340 16294
rect 15364 16292 15420 16294
rect 15124 15258 15180 15260
rect 15204 15258 15260 15260
rect 15284 15258 15340 15260
rect 15364 15258 15420 15260
rect 15124 15206 15170 15258
rect 15170 15206 15180 15258
rect 15204 15206 15234 15258
rect 15234 15206 15246 15258
rect 15246 15206 15260 15258
rect 15284 15206 15298 15258
rect 15298 15206 15310 15258
rect 15310 15206 15340 15258
rect 15364 15206 15374 15258
rect 15374 15206 15420 15258
rect 15124 15204 15180 15206
rect 15204 15204 15260 15206
rect 15284 15204 15340 15206
rect 15364 15204 15420 15206
rect 16394 15408 16450 15464
rect 15124 14170 15180 14172
rect 15204 14170 15260 14172
rect 15284 14170 15340 14172
rect 15364 14170 15420 14172
rect 15124 14118 15170 14170
rect 15170 14118 15180 14170
rect 15204 14118 15234 14170
rect 15234 14118 15246 14170
rect 15246 14118 15260 14170
rect 15284 14118 15298 14170
rect 15298 14118 15310 14170
rect 15310 14118 15340 14170
rect 15364 14118 15374 14170
rect 15374 14118 15420 14170
rect 15124 14116 15180 14118
rect 15204 14116 15260 14118
rect 15284 14116 15340 14118
rect 15364 14116 15420 14118
rect 15124 13082 15180 13084
rect 15204 13082 15260 13084
rect 15284 13082 15340 13084
rect 15364 13082 15420 13084
rect 15124 13030 15170 13082
rect 15170 13030 15180 13082
rect 15204 13030 15234 13082
rect 15234 13030 15246 13082
rect 15246 13030 15260 13082
rect 15284 13030 15298 13082
rect 15298 13030 15310 13082
rect 15310 13030 15340 13082
rect 15364 13030 15374 13082
rect 15374 13030 15420 13082
rect 15124 13028 15180 13030
rect 15204 13028 15260 13030
rect 15284 13028 15340 13030
rect 15364 13028 15420 13030
rect 14554 10668 14610 10704
rect 14554 10648 14556 10668
rect 14556 10648 14608 10668
rect 14608 10648 14610 10668
rect 14370 10512 14426 10568
rect 17130 17740 17186 17776
rect 17130 17720 17132 17740
rect 17132 17720 17184 17740
rect 17184 17720 17186 17740
rect 15382 12164 15438 12200
rect 15382 12144 15384 12164
rect 15384 12144 15436 12164
rect 15436 12144 15438 12164
rect 15124 11994 15180 11996
rect 15204 11994 15260 11996
rect 15284 11994 15340 11996
rect 15364 11994 15420 11996
rect 15124 11942 15170 11994
rect 15170 11942 15180 11994
rect 15204 11942 15234 11994
rect 15234 11942 15246 11994
rect 15246 11942 15260 11994
rect 15284 11942 15298 11994
rect 15298 11942 15310 11994
rect 15310 11942 15340 11994
rect 15364 11942 15374 11994
rect 15374 11942 15420 11994
rect 15124 11940 15180 11942
rect 15204 11940 15260 11942
rect 15284 11940 15340 11942
rect 15364 11940 15420 11942
rect 15124 10906 15180 10908
rect 15204 10906 15260 10908
rect 15284 10906 15340 10908
rect 15364 10906 15420 10908
rect 15124 10854 15170 10906
rect 15170 10854 15180 10906
rect 15204 10854 15234 10906
rect 15234 10854 15246 10906
rect 15246 10854 15260 10906
rect 15284 10854 15298 10906
rect 15298 10854 15310 10906
rect 15310 10854 15340 10906
rect 15364 10854 15374 10906
rect 15374 10854 15420 10906
rect 15124 10852 15180 10854
rect 15204 10852 15260 10854
rect 15284 10852 15340 10854
rect 15364 10852 15420 10854
rect 15124 9818 15180 9820
rect 15204 9818 15260 9820
rect 15284 9818 15340 9820
rect 15364 9818 15420 9820
rect 15124 9766 15170 9818
rect 15170 9766 15180 9818
rect 15204 9766 15234 9818
rect 15234 9766 15246 9818
rect 15246 9766 15260 9818
rect 15284 9766 15298 9818
rect 15298 9766 15310 9818
rect 15310 9766 15340 9818
rect 15364 9766 15374 9818
rect 15374 9766 15420 9818
rect 15124 9764 15180 9766
rect 15204 9764 15260 9766
rect 15284 9764 15340 9766
rect 15364 9764 15420 9766
rect 15290 9580 15346 9616
rect 15290 9560 15292 9580
rect 15292 9560 15344 9580
rect 15344 9560 15346 9580
rect 15124 8730 15180 8732
rect 15204 8730 15260 8732
rect 15284 8730 15340 8732
rect 15364 8730 15420 8732
rect 15124 8678 15170 8730
rect 15170 8678 15180 8730
rect 15204 8678 15234 8730
rect 15234 8678 15246 8730
rect 15246 8678 15260 8730
rect 15284 8678 15298 8730
rect 15298 8678 15310 8730
rect 15310 8678 15340 8730
rect 15364 8678 15374 8730
rect 15374 8678 15420 8730
rect 15124 8676 15180 8678
rect 15204 8676 15260 8678
rect 15284 8676 15340 8678
rect 15364 8676 15420 8678
rect 15124 7642 15180 7644
rect 15204 7642 15260 7644
rect 15284 7642 15340 7644
rect 15364 7642 15420 7644
rect 15124 7590 15170 7642
rect 15170 7590 15180 7642
rect 15204 7590 15234 7642
rect 15234 7590 15246 7642
rect 15246 7590 15260 7642
rect 15284 7590 15298 7642
rect 15298 7590 15310 7642
rect 15310 7590 15340 7642
rect 15364 7590 15374 7642
rect 15374 7590 15420 7642
rect 15124 7588 15180 7590
rect 15204 7588 15260 7590
rect 15284 7588 15340 7590
rect 15364 7588 15420 7590
rect 15124 6554 15180 6556
rect 15204 6554 15260 6556
rect 15284 6554 15340 6556
rect 15364 6554 15420 6556
rect 15124 6502 15170 6554
rect 15170 6502 15180 6554
rect 15204 6502 15234 6554
rect 15234 6502 15246 6554
rect 15246 6502 15260 6554
rect 15284 6502 15298 6554
rect 15298 6502 15310 6554
rect 15310 6502 15340 6554
rect 15364 6502 15374 6554
rect 15374 6502 15420 6554
rect 15124 6500 15180 6502
rect 15204 6500 15260 6502
rect 15284 6500 15340 6502
rect 15364 6500 15420 6502
rect 18050 19352 18106 19408
rect 18666 27770 18722 27772
rect 18746 27770 18802 27772
rect 18826 27770 18882 27772
rect 18906 27770 18962 27772
rect 18666 27718 18712 27770
rect 18712 27718 18722 27770
rect 18746 27718 18776 27770
rect 18776 27718 18788 27770
rect 18788 27718 18802 27770
rect 18826 27718 18840 27770
rect 18840 27718 18852 27770
rect 18852 27718 18882 27770
rect 18906 27718 18916 27770
rect 18916 27718 18962 27770
rect 18666 27716 18722 27718
rect 18746 27716 18802 27718
rect 18826 27716 18882 27718
rect 18906 27716 18962 27718
rect 18666 26682 18722 26684
rect 18746 26682 18802 26684
rect 18826 26682 18882 26684
rect 18906 26682 18962 26684
rect 18666 26630 18712 26682
rect 18712 26630 18722 26682
rect 18746 26630 18776 26682
rect 18776 26630 18788 26682
rect 18788 26630 18802 26682
rect 18826 26630 18840 26682
rect 18840 26630 18852 26682
rect 18852 26630 18882 26682
rect 18906 26630 18916 26682
rect 18916 26630 18962 26682
rect 18666 26628 18722 26630
rect 18746 26628 18802 26630
rect 18826 26628 18882 26630
rect 18906 26628 18962 26630
rect 18666 25594 18722 25596
rect 18746 25594 18802 25596
rect 18826 25594 18882 25596
rect 18906 25594 18962 25596
rect 18666 25542 18712 25594
rect 18712 25542 18722 25594
rect 18746 25542 18776 25594
rect 18776 25542 18788 25594
rect 18788 25542 18802 25594
rect 18826 25542 18840 25594
rect 18840 25542 18852 25594
rect 18852 25542 18882 25594
rect 18906 25542 18916 25594
rect 18916 25542 18962 25594
rect 18666 25540 18722 25542
rect 18746 25540 18802 25542
rect 18826 25540 18882 25542
rect 18906 25540 18962 25542
rect 19890 26968 19946 27024
rect 18666 24506 18722 24508
rect 18746 24506 18802 24508
rect 18826 24506 18882 24508
rect 18906 24506 18962 24508
rect 18666 24454 18712 24506
rect 18712 24454 18722 24506
rect 18746 24454 18776 24506
rect 18776 24454 18788 24506
rect 18788 24454 18802 24506
rect 18826 24454 18840 24506
rect 18840 24454 18852 24506
rect 18852 24454 18882 24506
rect 18906 24454 18916 24506
rect 18916 24454 18962 24506
rect 18666 24452 18722 24454
rect 18746 24452 18802 24454
rect 18826 24452 18882 24454
rect 18906 24452 18962 24454
rect 18666 23418 18722 23420
rect 18746 23418 18802 23420
rect 18826 23418 18882 23420
rect 18906 23418 18962 23420
rect 18666 23366 18712 23418
rect 18712 23366 18722 23418
rect 18746 23366 18776 23418
rect 18776 23366 18788 23418
rect 18788 23366 18802 23418
rect 18826 23366 18840 23418
rect 18840 23366 18852 23418
rect 18852 23366 18882 23418
rect 18906 23366 18916 23418
rect 18916 23366 18962 23418
rect 18666 23364 18722 23366
rect 18746 23364 18802 23366
rect 18826 23364 18882 23366
rect 18906 23364 18962 23366
rect 18666 22330 18722 22332
rect 18746 22330 18802 22332
rect 18826 22330 18882 22332
rect 18906 22330 18962 22332
rect 18666 22278 18712 22330
rect 18712 22278 18722 22330
rect 18746 22278 18776 22330
rect 18776 22278 18788 22330
rect 18788 22278 18802 22330
rect 18826 22278 18840 22330
rect 18840 22278 18852 22330
rect 18852 22278 18882 22330
rect 18906 22278 18916 22330
rect 18916 22278 18962 22330
rect 18666 22276 18722 22278
rect 18746 22276 18802 22278
rect 18826 22276 18882 22278
rect 18906 22276 18962 22278
rect 18970 21800 19026 21856
rect 18666 21242 18722 21244
rect 18746 21242 18802 21244
rect 18826 21242 18882 21244
rect 18906 21242 18962 21244
rect 18666 21190 18712 21242
rect 18712 21190 18722 21242
rect 18746 21190 18776 21242
rect 18776 21190 18788 21242
rect 18788 21190 18802 21242
rect 18826 21190 18840 21242
rect 18840 21190 18852 21242
rect 18852 21190 18882 21242
rect 18906 21190 18916 21242
rect 18916 21190 18962 21242
rect 18666 21188 18722 21190
rect 18746 21188 18802 21190
rect 18826 21188 18882 21190
rect 18906 21188 18962 21190
rect 18666 20154 18722 20156
rect 18746 20154 18802 20156
rect 18826 20154 18882 20156
rect 18906 20154 18962 20156
rect 18666 20102 18712 20154
rect 18712 20102 18722 20154
rect 18746 20102 18776 20154
rect 18776 20102 18788 20154
rect 18788 20102 18802 20154
rect 18826 20102 18840 20154
rect 18840 20102 18852 20154
rect 18852 20102 18882 20154
rect 18906 20102 18916 20154
rect 18916 20102 18962 20154
rect 18666 20100 18722 20102
rect 18746 20100 18802 20102
rect 18826 20100 18882 20102
rect 18906 20100 18962 20102
rect 18666 19066 18722 19068
rect 18746 19066 18802 19068
rect 18826 19066 18882 19068
rect 18906 19066 18962 19068
rect 18666 19014 18712 19066
rect 18712 19014 18722 19066
rect 18746 19014 18776 19066
rect 18776 19014 18788 19066
rect 18788 19014 18802 19066
rect 18826 19014 18840 19066
rect 18840 19014 18852 19066
rect 18852 19014 18882 19066
rect 18906 19014 18916 19066
rect 18916 19014 18962 19066
rect 18666 19012 18722 19014
rect 18746 19012 18802 19014
rect 18826 19012 18882 19014
rect 18906 19012 18962 19014
rect 18666 17978 18722 17980
rect 18746 17978 18802 17980
rect 18826 17978 18882 17980
rect 18906 17978 18962 17980
rect 18666 17926 18712 17978
rect 18712 17926 18722 17978
rect 18746 17926 18776 17978
rect 18776 17926 18788 17978
rect 18788 17926 18802 17978
rect 18826 17926 18840 17978
rect 18840 17926 18852 17978
rect 18852 17926 18882 17978
rect 18906 17926 18916 17978
rect 18916 17926 18962 17978
rect 18666 17924 18722 17926
rect 18746 17924 18802 17926
rect 18826 17924 18882 17926
rect 18906 17924 18962 17926
rect 18050 14884 18106 14920
rect 18050 14864 18052 14884
rect 18052 14864 18104 14884
rect 18104 14864 18106 14884
rect 16670 7284 16672 7304
rect 16672 7284 16724 7304
rect 16724 7284 16726 7304
rect 16670 7248 16726 7284
rect 16578 6160 16634 6216
rect 15124 5466 15180 5468
rect 15204 5466 15260 5468
rect 15284 5466 15340 5468
rect 15364 5466 15420 5468
rect 15124 5414 15170 5466
rect 15170 5414 15180 5466
rect 15204 5414 15234 5466
rect 15234 5414 15246 5466
rect 15246 5414 15260 5466
rect 15284 5414 15298 5466
rect 15298 5414 15310 5466
rect 15310 5414 15340 5466
rect 15364 5414 15374 5466
rect 15374 5414 15420 5466
rect 15124 5412 15180 5414
rect 15204 5412 15260 5414
rect 15284 5412 15340 5414
rect 15364 5412 15420 5414
rect 15124 4378 15180 4380
rect 15204 4378 15260 4380
rect 15284 4378 15340 4380
rect 15364 4378 15420 4380
rect 15124 4326 15170 4378
rect 15170 4326 15180 4378
rect 15204 4326 15234 4378
rect 15234 4326 15246 4378
rect 15246 4326 15260 4378
rect 15284 4326 15298 4378
rect 15298 4326 15310 4378
rect 15310 4326 15340 4378
rect 15364 4326 15374 4378
rect 15374 4326 15420 4378
rect 15124 4324 15180 4326
rect 15204 4324 15260 4326
rect 15284 4324 15340 4326
rect 15364 4324 15420 4326
rect 16394 3476 16396 3496
rect 16396 3476 16448 3496
rect 16448 3476 16450 3496
rect 16394 3440 16450 3476
rect 18510 17720 18566 17776
rect 18666 16890 18722 16892
rect 18746 16890 18802 16892
rect 18826 16890 18882 16892
rect 18906 16890 18962 16892
rect 18666 16838 18712 16890
rect 18712 16838 18722 16890
rect 18746 16838 18776 16890
rect 18776 16838 18788 16890
rect 18788 16838 18802 16890
rect 18826 16838 18840 16890
rect 18840 16838 18852 16890
rect 18852 16838 18882 16890
rect 18906 16838 18916 16890
rect 18916 16838 18962 16890
rect 18666 16836 18722 16838
rect 18746 16836 18802 16838
rect 18826 16836 18882 16838
rect 18906 16836 18962 16838
rect 18666 15802 18722 15804
rect 18746 15802 18802 15804
rect 18826 15802 18882 15804
rect 18906 15802 18962 15804
rect 18666 15750 18712 15802
rect 18712 15750 18722 15802
rect 18746 15750 18776 15802
rect 18776 15750 18788 15802
rect 18788 15750 18802 15802
rect 18826 15750 18840 15802
rect 18840 15750 18852 15802
rect 18852 15750 18882 15802
rect 18906 15750 18916 15802
rect 18916 15750 18962 15802
rect 18666 15748 18722 15750
rect 18746 15748 18802 15750
rect 18826 15748 18882 15750
rect 18906 15748 18962 15750
rect 18666 14714 18722 14716
rect 18746 14714 18802 14716
rect 18826 14714 18882 14716
rect 18906 14714 18962 14716
rect 18666 14662 18712 14714
rect 18712 14662 18722 14714
rect 18746 14662 18776 14714
rect 18776 14662 18788 14714
rect 18788 14662 18802 14714
rect 18826 14662 18840 14714
rect 18840 14662 18852 14714
rect 18852 14662 18882 14714
rect 18906 14662 18916 14714
rect 18916 14662 18962 14714
rect 18666 14660 18722 14662
rect 18746 14660 18802 14662
rect 18826 14660 18882 14662
rect 18906 14660 18962 14662
rect 18666 13626 18722 13628
rect 18746 13626 18802 13628
rect 18826 13626 18882 13628
rect 18906 13626 18962 13628
rect 18666 13574 18712 13626
rect 18712 13574 18722 13626
rect 18746 13574 18776 13626
rect 18776 13574 18788 13626
rect 18788 13574 18802 13626
rect 18826 13574 18840 13626
rect 18840 13574 18852 13626
rect 18852 13574 18882 13626
rect 18906 13574 18916 13626
rect 18916 13574 18962 13626
rect 18666 13572 18722 13574
rect 18746 13572 18802 13574
rect 18826 13572 18882 13574
rect 18906 13572 18962 13574
rect 18666 12538 18722 12540
rect 18746 12538 18802 12540
rect 18826 12538 18882 12540
rect 18906 12538 18962 12540
rect 18666 12486 18712 12538
rect 18712 12486 18722 12538
rect 18746 12486 18776 12538
rect 18776 12486 18788 12538
rect 18788 12486 18802 12538
rect 18826 12486 18840 12538
rect 18840 12486 18852 12538
rect 18852 12486 18882 12538
rect 18906 12486 18916 12538
rect 18916 12486 18962 12538
rect 18666 12484 18722 12486
rect 18746 12484 18802 12486
rect 18826 12484 18882 12486
rect 18906 12484 18962 12486
rect 18418 12280 18474 12336
rect 18666 11450 18722 11452
rect 18746 11450 18802 11452
rect 18826 11450 18882 11452
rect 18906 11450 18962 11452
rect 18666 11398 18712 11450
rect 18712 11398 18722 11450
rect 18746 11398 18776 11450
rect 18776 11398 18788 11450
rect 18788 11398 18802 11450
rect 18826 11398 18840 11450
rect 18840 11398 18852 11450
rect 18852 11398 18882 11450
rect 18906 11398 18916 11450
rect 18916 11398 18962 11450
rect 18666 11396 18722 11398
rect 18746 11396 18802 11398
rect 18826 11396 18882 11398
rect 18906 11396 18962 11398
rect 18326 10648 18382 10704
rect 17682 3476 17684 3496
rect 17684 3476 17736 3496
rect 17736 3476 17738 3496
rect 17682 3440 17738 3476
rect 15124 3290 15180 3292
rect 15204 3290 15260 3292
rect 15284 3290 15340 3292
rect 15364 3290 15420 3292
rect 15124 3238 15170 3290
rect 15170 3238 15180 3290
rect 15204 3238 15234 3290
rect 15234 3238 15246 3290
rect 15246 3238 15260 3290
rect 15284 3238 15298 3290
rect 15298 3238 15310 3290
rect 15310 3238 15340 3290
rect 15364 3238 15374 3290
rect 15374 3238 15420 3290
rect 15124 3236 15180 3238
rect 15204 3236 15260 3238
rect 15284 3236 15340 3238
rect 15364 3236 15420 3238
rect 18666 10362 18722 10364
rect 18746 10362 18802 10364
rect 18826 10362 18882 10364
rect 18906 10362 18962 10364
rect 18666 10310 18712 10362
rect 18712 10310 18722 10362
rect 18746 10310 18776 10362
rect 18776 10310 18788 10362
rect 18788 10310 18802 10362
rect 18826 10310 18840 10362
rect 18840 10310 18852 10362
rect 18852 10310 18882 10362
rect 18906 10310 18916 10362
rect 18916 10310 18962 10362
rect 18666 10308 18722 10310
rect 18746 10308 18802 10310
rect 18826 10308 18882 10310
rect 18906 10308 18962 10310
rect 19338 10004 19340 10024
rect 19340 10004 19392 10024
rect 19392 10004 19394 10024
rect 19338 9968 19394 10004
rect 18666 9274 18722 9276
rect 18746 9274 18802 9276
rect 18826 9274 18882 9276
rect 18906 9274 18962 9276
rect 18666 9222 18712 9274
rect 18712 9222 18722 9274
rect 18746 9222 18776 9274
rect 18776 9222 18788 9274
rect 18788 9222 18802 9274
rect 18826 9222 18840 9274
rect 18840 9222 18852 9274
rect 18852 9222 18882 9274
rect 18906 9222 18916 9274
rect 18916 9222 18962 9274
rect 18666 9220 18722 9222
rect 18746 9220 18802 9222
rect 18826 9220 18882 9222
rect 18906 9220 18962 9222
rect 18666 8186 18722 8188
rect 18746 8186 18802 8188
rect 18826 8186 18882 8188
rect 18906 8186 18962 8188
rect 18666 8134 18712 8186
rect 18712 8134 18722 8186
rect 18746 8134 18776 8186
rect 18776 8134 18788 8186
rect 18788 8134 18802 8186
rect 18826 8134 18840 8186
rect 18840 8134 18852 8186
rect 18852 8134 18882 8186
rect 18906 8134 18916 8186
rect 18916 8134 18962 8186
rect 18666 8132 18722 8134
rect 18746 8132 18802 8134
rect 18826 8132 18882 8134
rect 18906 8132 18962 8134
rect 18666 7098 18722 7100
rect 18746 7098 18802 7100
rect 18826 7098 18882 7100
rect 18906 7098 18962 7100
rect 18666 7046 18712 7098
rect 18712 7046 18722 7098
rect 18746 7046 18776 7098
rect 18776 7046 18788 7098
rect 18788 7046 18802 7098
rect 18826 7046 18840 7098
rect 18840 7046 18852 7098
rect 18852 7046 18882 7098
rect 18906 7046 18916 7098
rect 18916 7046 18962 7098
rect 18666 7044 18722 7046
rect 18746 7044 18802 7046
rect 18826 7044 18882 7046
rect 18906 7044 18962 7046
rect 18666 6010 18722 6012
rect 18746 6010 18802 6012
rect 18826 6010 18882 6012
rect 18906 6010 18962 6012
rect 18666 5958 18712 6010
rect 18712 5958 18722 6010
rect 18746 5958 18776 6010
rect 18776 5958 18788 6010
rect 18788 5958 18802 6010
rect 18826 5958 18840 6010
rect 18840 5958 18852 6010
rect 18852 5958 18882 6010
rect 18906 5958 18916 6010
rect 18916 5958 18962 6010
rect 18666 5956 18722 5958
rect 18746 5956 18802 5958
rect 18826 5956 18882 5958
rect 18906 5956 18962 5958
rect 19522 6860 19578 6896
rect 19522 6840 19524 6860
rect 19524 6840 19576 6860
rect 19576 6840 19578 6860
rect 18666 4922 18722 4924
rect 18746 4922 18802 4924
rect 18826 4922 18882 4924
rect 18906 4922 18962 4924
rect 18666 4870 18712 4922
rect 18712 4870 18722 4922
rect 18746 4870 18776 4922
rect 18776 4870 18788 4922
rect 18788 4870 18802 4922
rect 18826 4870 18840 4922
rect 18840 4870 18852 4922
rect 18852 4870 18882 4922
rect 18906 4870 18916 4922
rect 18916 4870 18962 4922
rect 18666 4868 18722 4870
rect 18746 4868 18802 4870
rect 18826 4868 18882 4870
rect 18906 4868 18962 4870
rect 18666 3834 18722 3836
rect 18746 3834 18802 3836
rect 18826 3834 18882 3836
rect 18906 3834 18962 3836
rect 18666 3782 18712 3834
rect 18712 3782 18722 3834
rect 18746 3782 18776 3834
rect 18776 3782 18788 3834
rect 18788 3782 18802 3834
rect 18826 3782 18840 3834
rect 18840 3782 18852 3834
rect 18852 3782 18882 3834
rect 18906 3782 18916 3834
rect 18916 3782 18962 3834
rect 18666 3780 18722 3782
rect 18746 3780 18802 3782
rect 18826 3780 18882 3782
rect 18906 3780 18962 3782
rect 18666 2746 18722 2748
rect 18746 2746 18802 2748
rect 18826 2746 18882 2748
rect 18906 2746 18962 2748
rect 18666 2694 18712 2746
rect 18712 2694 18722 2746
rect 18746 2694 18776 2746
rect 18776 2694 18788 2746
rect 18788 2694 18802 2746
rect 18826 2694 18840 2746
rect 18840 2694 18852 2746
rect 18852 2694 18882 2746
rect 18906 2694 18916 2746
rect 18916 2694 18962 2746
rect 18666 2692 18722 2694
rect 18746 2692 18802 2694
rect 18826 2692 18882 2694
rect 18906 2692 18962 2694
rect 20166 26988 20222 27024
rect 20166 26968 20168 26988
rect 20168 26968 20220 26988
rect 20220 26968 20222 26988
rect 22208 29402 22264 29404
rect 22288 29402 22344 29404
rect 22368 29402 22424 29404
rect 22448 29402 22504 29404
rect 22208 29350 22254 29402
rect 22254 29350 22264 29402
rect 22288 29350 22318 29402
rect 22318 29350 22330 29402
rect 22330 29350 22344 29402
rect 22368 29350 22382 29402
rect 22382 29350 22394 29402
rect 22394 29350 22424 29402
rect 22448 29350 22458 29402
rect 22458 29350 22504 29402
rect 22208 29348 22264 29350
rect 22288 29348 22344 29350
rect 22368 29348 22424 29350
rect 22448 29348 22504 29350
rect 22208 28314 22264 28316
rect 22288 28314 22344 28316
rect 22368 28314 22424 28316
rect 22448 28314 22504 28316
rect 22208 28262 22254 28314
rect 22254 28262 22264 28314
rect 22288 28262 22318 28314
rect 22318 28262 22330 28314
rect 22330 28262 22344 28314
rect 22368 28262 22382 28314
rect 22382 28262 22394 28314
rect 22394 28262 22424 28314
rect 22448 28262 22458 28314
rect 22458 28262 22504 28314
rect 22208 28260 22264 28262
rect 22288 28260 22344 28262
rect 22368 28260 22424 28262
rect 22448 28260 22504 28262
rect 22208 27226 22264 27228
rect 22288 27226 22344 27228
rect 22368 27226 22424 27228
rect 22448 27226 22504 27228
rect 22208 27174 22254 27226
rect 22254 27174 22264 27226
rect 22288 27174 22318 27226
rect 22318 27174 22330 27226
rect 22330 27174 22344 27226
rect 22368 27174 22382 27226
rect 22382 27174 22394 27226
rect 22394 27174 22424 27226
rect 22448 27174 22458 27226
rect 22458 27174 22504 27226
rect 22208 27172 22264 27174
rect 22288 27172 22344 27174
rect 22368 27172 22424 27174
rect 22448 27172 22504 27174
rect 22650 26424 22706 26480
rect 22558 26288 22614 26344
rect 22208 26138 22264 26140
rect 22288 26138 22344 26140
rect 22368 26138 22424 26140
rect 22448 26138 22504 26140
rect 22208 26086 22254 26138
rect 22254 26086 22264 26138
rect 22288 26086 22318 26138
rect 22318 26086 22330 26138
rect 22330 26086 22344 26138
rect 22368 26086 22382 26138
rect 22382 26086 22394 26138
rect 22394 26086 22424 26138
rect 22448 26086 22458 26138
rect 22458 26086 22504 26138
rect 22208 26084 22264 26086
rect 22288 26084 22344 26086
rect 22368 26084 22424 26086
rect 22448 26084 22504 26086
rect 22208 25050 22264 25052
rect 22288 25050 22344 25052
rect 22368 25050 22424 25052
rect 22448 25050 22504 25052
rect 22208 24998 22254 25050
rect 22254 24998 22264 25050
rect 22288 24998 22318 25050
rect 22318 24998 22330 25050
rect 22330 24998 22344 25050
rect 22368 24998 22382 25050
rect 22382 24998 22394 25050
rect 22394 24998 22424 25050
rect 22448 24998 22458 25050
rect 22458 24998 22504 25050
rect 22208 24996 22264 24998
rect 22288 24996 22344 24998
rect 22368 24996 22424 24998
rect 22448 24996 22504 24998
rect 21086 22924 21088 22944
rect 21088 22924 21140 22944
rect 21140 22924 21142 22944
rect 21086 22888 21142 22924
rect 21178 22072 21234 22128
rect 21178 21800 21234 21856
rect 20258 15952 20314 16008
rect 20074 8508 20076 8528
rect 20076 8508 20128 8528
rect 20128 8508 20130 8528
rect 20074 8472 20130 8508
rect 19982 6840 20038 6896
rect 20718 17992 20774 18048
rect 20626 16632 20682 16688
rect 20626 14592 20682 14648
rect 20902 12960 20958 13016
rect 22208 23962 22264 23964
rect 22288 23962 22344 23964
rect 22368 23962 22424 23964
rect 22448 23962 22504 23964
rect 22208 23910 22254 23962
rect 22254 23910 22264 23962
rect 22288 23910 22318 23962
rect 22318 23910 22330 23962
rect 22330 23910 22344 23962
rect 22368 23910 22382 23962
rect 22382 23910 22394 23962
rect 22394 23910 22424 23962
rect 22448 23910 22458 23962
rect 22458 23910 22504 23962
rect 22208 23908 22264 23910
rect 22288 23908 22344 23910
rect 22368 23908 22424 23910
rect 22448 23908 22504 23910
rect 22208 22874 22264 22876
rect 22288 22874 22344 22876
rect 22368 22874 22424 22876
rect 22448 22874 22504 22876
rect 22208 22822 22254 22874
rect 22254 22822 22264 22874
rect 22288 22822 22318 22874
rect 22318 22822 22330 22874
rect 22330 22822 22344 22874
rect 22368 22822 22382 22874
rect 22382 22822 22394 22874
rect 22394 22822 22424 22874
rect 22448 22822 22458 22874
rect 22458 22822 22504 22874
rect 22208 22820 22264 22822
rect 22288 22820 22344 22822
rect 22368 22820 22424 22822
rect 22448 22820 22504 22822
rect 22208 21786 22264 21788
rect 22288 21786 22344 21788
rect 22368 21786 22424 21788
rect 22448 21786 22504 21788
rect 22208 21734 22254 21786
rect 22254 21734 22264 21786
rect 22288 21734 22318 21786
rect 22318 21734 22330 21786
rect 22330 21734 22344 21786
rect 22368 21734 22382 21786
rect 22382 21734 22394 21786
rect 22394 21734 22424 21786
rect 22448 21734 22458 21786
rect 22458 21734 22504 21786
rect 22208 21732 22264 21734
rect 22288 21732 22344 21734
rect 22368 21732 22424 21734
rect 22448 21732 22504 21734
rect 22208 20698 22264 20700
rect 22288 20698 22344 20700
rect 22368 20698 22424 20700
rect 22448 20698 22504 20700
rect 22208 20646 22254 20698
rect 22254 20646 22264 20698
rect 22288 20646 22318 20698
rect 22318 20646 22330 20698
rect 22330 20646 22344 20698
rect 22368 20646 22382 20698
rect 22382 20646 22394 20698
rect 22394 20646 22424 20698
rect 22448 20646 22458 20698
rect 22458 20646 22504 20698
rect 22208 20644 22264 20646
rect 22288 20644 22344 20646
rect 22368 20644 22424 20646
rect 22448 20644 22504 20646
rect 22208 19610 22264 19612
rect 22288 19610 22344 19612
rect 22368 19610 22424 19612
rect 22448 19610 22504 19612
rect 22208 19558 22254 19610
rect 22254 19558 22264 19610
rect 22288 19558 22318 19610
rect 22318 19558 22330 19610
rect 22330 19558 22344 19610
rect 22368 19558 22382 19610
rect 22382 19558 22394 19610
rect 22394 19558 22424 19610
rect 22448 19558 22458 19610
rect 22458 19558 22504 19610
rect 22208 19556 22264 19558
rect 22288 19556 22344 19558
rect 22368 19556 22424 19558
rect 22448 19556 22504 19558
rect 21638 14592 21694 14648
rect 22208 18522 22264 18524
rect 22288 18522 22344 18524
rect 22368 18522 22424 18524
rect 22448 18522 22504 18524
rect 22208 18470 22254 18522
rect 22254 18470 22264 18522
rect 22288 18470 22318 18522
rect 22318 18470 22330 18522
rect 22330 18470 22344 18522
rect 22368 18470 22382 18522
rect 22382 18470 22394 18522
rect 22394 18470 22424 18522
rect 22448 18470 22458 18522
rect 22458 18470 22504 18522
rect 22208 18468 22264 18470
rect 22288 18468 22344 18470
rect 22368 18468 22424 18470
rect 22448 18468 22504 18470
rect 22208 17434 22264 17436
rect 22288 17434 22344 17436
rect 22368 17434 22424 17436
rect 22448 17434 22504 17436
rect 22208 17382 22254 17434
rect 22254 17382 22264 17434
rect 22288 17382 22318 17434
rect 22318 17382 22330 17434
rect 22330 17382 22344 17434
rect 22368 17382 22382 17434
rect 22382 17382 22394 17434
rect 22394 17382 22424 17434
rect 22448 17382 22458 17434
rect 22458 17382 22504 17434
rect 22208 17380 22264 17382
rect 22288 17380 22344 17382
rect 22368 17380 22424 17382
rect 22448 17380 22504 17382
rect 22208 16346 22264 16348
rect 22288 16346 22344 16348
rect 22368 16346 22424 16348
rect 22448 16346 22504 16348
rect 22208 16294 22254 16346
rect 22254 16294 22264 16346
rect 22288 16294 22318 16346
rect 22318 16294 22330 16346
rect 22330 16294 22344 16346
rect 22368 16294 22382 16346
rect 22382 16294 22394 16346
rect 22394 16294 22424 16346
rect 22448 16294 22458 16346
rect 22458 16294 22504 16346
rect 22208 16292 22264 16294
rect 22288 16292 22344 16294
rect 22368 16292 22424 16294
rect 22448 16292 22504 16294
rect 22208 15258 22264 15260
rect 22288 15258 22344 15260
rect 22368 15258 22424 15260
rect 22448 15258 22504 15260
rect 22208 15206 22254 15258
rect 22254 15206 22264 15258
rect 22288 15206 22318 15258
rect 22318 15206 22330 15258
rect 22330 15206 22344 15258
rect 22368 15206 22382 15258
rect 22382 15206 22394 15258
rect 22394 15206 22424 15258
rect 22448 15206 22458 15258
rect 22458 15206 22504 15258
rect 22208 15204 22264 15206
rect 22288 15204 22344 15206
rect 22368 15204 22424 15206
rect 22448 15204 22504 15206
rect 22208 14170 22264 14172
rect 22288 14170 22344 14172
rect 22368 14170 22424 14172
rect 22448 14170 22504 14172
rect 22208 14118 22254 14170
rect 22254 14118 22264 14170
rect 22288 14118 22318 14170
rect 22318 14118 22330 14170
rect 22330 14118 22344 14170
rect 22368 14118 22382 14170
rect 22382 14118 22394 14170
rect 22394 14118 22424 14170
rect 22448 14118 22458 14170
rect 22458 14118 22504 14170
rect 22208 14116 22264 14118
rect 22288 14116 22344 14118
rect 22368 14116 22424 14118
rect 22448 14116 22504 14118
rect 22208 13082 22264 13084
rect 22288 13082 22344 13084
rect 22368 13082 22424 13084
rect 22448 13082 22504 13084
rect 22208 13030 22254 13082
rect 22254 13030 22264 13082
rect 22288 13030 22318 13082
rect 22318 13030 22330 13082
rect 22330 13030 22344 13082
rect 22368 13030 22382 13082
rect 22382 13030 22394 13082
rect 22394 13030 22424 13082
rect 22448 13030 22458 13082
rect 22458 13030 22504 13082
rect 22208 13028 22264 13030
rect 22288 13028 22344 13030
rect 22368 13028 22424 13030
rect 22448 13028 22504 13030
rect 21638 10104 21694 10160
rect 20994 9424 21050 9480
rect 22208 11994 22264 11996
rect 22288 11994 22344 11996
rect 22368 11994 22424 11996
rect 22448 11994 22504 11996
rect 22208 11942 22254 11994
rect 22254 11942 22264 11994
rect 22288 11942 22318 11994
rect 22318 11942 22330 11994
rect 22330 11942 22344 11994
rect 22368 11942 22382 11994
rect 22382 11942 22394 11994
rect 22394 11942 22424 11994
rect 22448 11942 22458 11994
rect 22458 11942 22504 11994
rect 22208 11940 22264 11942
rect 22288 11940 22344 11942
rect 22368 11940 22424 11942
rect 22448 11940 22504 11942
rect 22208 10906 22264 10908
rect 22288 10906 22344 10908
rect 22368 10906 22424 10908
rect 22448 10906 22504 10908
rect 22208 10854 22254 10906
rect 22254 10854 22264 10906
rect 22288 10854 22318 10906
rect 22318 10854 22330 10906
rect 22330 10854 22344 10906
rect 22368 10854 22382 10906
rect 22382 10854 22394 10906
rect 22394 10854 22424 10906
rect 22448 10854 22458 10906
rect 22458 10854 22504 10906
rect 22208 10852 22264 10854
rect 22288 10852 22344 10854
rect 22368 10852 22424 10854
rect 22448 10852 22504 10854
rect 22208 9818 22264 9820
rect 22288 9818 22344 9820
rect 22368 9818 22424 9820
rect 22448 9818 22504 9820
rect 22208 9766 22254 9818
rect 22254 9766 22264 9818
rect 22288 9766 22318 9818
rect 22318 9766 22330 9818
rect 22330 9766 22344 9818
rect 22368 9766 22382 9818
rect 22382 9766 22394 9818
rect 22394 9766 22424 9818
rect 22448 9766 22458 9818
rect 22458 9766 22504 9818
rect 22208 9764 22264 9766
rect 22288 9764 22344 9766
rect 22368 9764 22424 9766
rect 22448 9764 22504 9766
rect 22208 8730 22264 8732
rect 22288 8730 22344 8732
rect 22368 8730 22424 8732
rect 22448 8730 22504 8732
rect 22208 8678 22254 8730
rect 22254 8678 22264 8730
rect 22288 8678 22318 8730
rect 22318 8678 22330 8730
rect 22330 8678 22344 8730
rect 22368 8678 22382 8730
rect 22382 8678 22394 8730
rect 22394 8678 22424 8730
rect 22448 8678 22458 8730
rect 22458 8678 22504 8730
rect 22208 8676 22264 8678
rect 22288 8676 22344 8678
rect 22368 8676 22424 8678
rect 22448 8676 22504 8678
rect 21914 7812 21970 7848
rect 21914 7792 21916 7812
rect 21916 7792 21968 7812
rect 21968 7792 21970 7812
rect 22208 7642 22264 7644
rect 22288 7642 22344 7644
rect 22368 7642 22424 7644
rect 22448 7642 22504 7644
rect 22208 7590 22254 7642
rect 22254 7590 22264 7642
rect 22288 7590 22318 7642
rect 22318 7590 22330 7642
rect 22330 7590 22344 7642
rect 22368 7590 22382 7642
rect 22382 7590 22394 7642
rect 22394 7590 22424 7642
rect 22448 7590 22458 7642
rect 22458 7590 22504 7642
rect 22208 7588 22264 7590
rect 22288 7588 22344 7590
rect 22368 7588 22424 7590
rect 22448 7588 22504 7590
rect 1490 2080 1546 2136
rect 8040 2202 8096 2204
rect 8120 2202 8176 2204
rect 8200 2202 8256 2204
rect 8280 2202 8336 2204
rect 8040 2150 8086 2202
rect 8086 2150 8096 2202
rect 8120 2150 8150 2202
rect 8150 2150 8162 2202
rect 8162 2150 8176 2202
rect 8200 2150 8214 2202
rect 8214 2150 8226 2202
rect 8226 2150 8256 2202
rect 8280 2150 8290 2202
rect 8290 2150 8336 2202
rect 8040 2148 8096 2150
rect 8120 2148 8176 2150
rect 8200 2148 8256 2150
rect 8280 2148 8336 2150
rect 15124 2202 15180 2204
rect 15204 2202 15260 2204
rect 15284 2202 15340 2204
rect 15364 2202 15420 2204
rect 15124 2150 15170 2202
rect 15170 2150 15180 2202
rect 15204 2150 15234 2202
rect 15234 2150 15246 2202
rect 15246 2150 15260 2202
rect 15284 2150 15298 2202
rect 15298 2150 15310 2202
rect 15310 2150 15340 2202
rect 15364 2150 15374 2202
rect 15374 2150 15420 2202
rect 15124 2148 15180 2150
rect 15204 2148 15260 2150
rect 15284 2148 15340 2150
rect 15364 2148 15420 2150
rect 22208 6554 22264 6556
rect 22288 6554 22344 6556
rect 22368 6554 22424 6556
rect 22448 6554 22504 6556
rect 22208 6502 22254 6554
rect 22254 6502 22264 6554
rect 22288 6502 22318 6554
rect 22318 6502 22330 6554
rect 22330 6502 22344 6554
rect 22368 6502 22382 6554
rect 22382 6502 22394 6554
rect 22394 6502 22424 6554
rect 22448 6502 22458 6554
rect 22458 6502 22504 6554
rect 22208 6500 22264 6502
rect 22288 6500 22344 6502
rect 22368 6500 22424 6502
rect 22448 6500 22504 6502
rect 22208 5466 22264 5468
rect 22288 5466 22344 5468
rect 22368 5466 22424 5468
rect 22448 5466 22504 5468
rect 22208 5414 22254 5466
rect 22254 5414 22264 5466
rect 22288 5414 22318 5466
rect 22318 5414 22330 5466
rect 22330 5414 22344 5466
rect 22368 5414 22382 5466
rect 22382 5414 22394 5466
rect 22394 5414 22424 5466
rect 22448 5414 22458 5466
rect 22458 5414 22504 5466
rect 22208 5412 22264 5414
rect 22288 5412 22344 5414
rect 22368 5412 22424 5414
rect 22448 5412 22504 5414
rect 22208 4378 22264 4380
rect 22288 4378 22344 4380
rect 22368 4378 22424 4380
rect 22448 4378 22504 4380
rect 22208 4326 22254 4378
rect 22254 4326 22264 4378
rect 22288 4326 22318 4378
rect 22318 4326 22330 4378
rect 22330 4326 22344 4378
rect 22368 4326 22382 4378
rect 22382 4326 22394 4378
rect 22394 4326 22424 4378
rect 22448 4326 22458 4378
rect 22458 4326 22504 4378
rect 22208 4324 22264 4326
rect 22288 4324 22344 4326
rect 22368 4324 22424 4326
rect 22448 4324 22504 4326
rect 24030 16496 24086 16552
rect 23938 11192 23994 11248
rect 23662 9968 23718 10024
rect 23478 9460 23480 9480
rect 23480 9460 23532 9480
rect 23532 9460 23534 9480
rect 23478 9424 23534 9460
rect 22208 3290 22264 3292
rect 22288 3290 22344 3292
rect 22368 3290 22424 3292
rect 22448 3290 22504 3292
rect 22208 3238 22254 3290
rect 22254 3238 22264 3290
rect 22288 3238 22318 3290
rect 22318 3238 22330 3290
rect 22330 3238 22344 3290
rect 22368 3238 22382 3290
rect 22382 3238 22394 3290
rect 22394 3238 22424 3290
rect 22448 3238 22458 3290
rect 22458 3238 22504 3290
rect 22208 3236 22264 3238
rect 22288 3236 22344 3238
rect 22368 3236 22424 3238
rect 22448 3236 22504 3238
rect 23478 5092 23534 5128
rect 23478 5072 23480 5092
rect 23480 5072 23532 5092
rect 23532 5072 23534 5092
rect 23478 4120 23534 4176
rect 25750 29946 25806 29948
rect 25830 29946 25886 29948
rect 25910 29946 25966 29948
rect 25990 29946 26046 29948
rect 25750 29894 25796 29946
rect 25796 29894 25806 29946
rect 25830 29894 25860 29946
rect 25860 29894 25872 29946
rect 25872 29894 25886 29946
rect 25910 29894 25924 29946
rect 25924 29894 25936 29946
rect 25936 29894 25966 29946
rect 25990 29894 26000 29946
rect 26000 29894 26046 29946
rect 25750 29892 25806 29894
rect 25830 29892 25886 29894
rect 25910 29892 25966 29894
rect 25990 29892 26046 29894
rect 25750 28858 25806 28860
rect 25830 28858 25886 28860
rect 25910 28858 25966 28860
rect 25990 28858 26046 28860
rect 25750 28806 25796 28858
rect 25796 28806 25806 28858
rect 25830 28806 25860 28858
rect 25860 28806 25872 28858
rect 25872 28806 25886 28858
rect 25910 28806 25924 28858
rect 25924 28806 25936 28858
rect 25936 28806 25966 28858
rect 25990 28806 26000 28858
rect 26000 28806 26046 28858
rect 25750 28804 25806 28806
rect 25830 28804 25886 28806
rect 25910 28804 25966 28806
rect 25990 28804 26046 28806
rect 27894 29996 27896 30016
rect 27896 29996 27948 30016
rect 27948 29996 27950 30016
rect 27894 29960 27950 29996
rect 27618 29280 27674 29336
rect 29292 30490 29348 30492
rect 29372 30490 29428 30492
rect 29452 30490 29508 30492
rect 29532 30490 29588 30492
rect 29292 30438 29338 30490
rect 29338 30438 29348 30490
rect 29372 30438 29402 30490
rect 29402 30438 29414 30490
rect 29414 30438 29428 30490
rect 29452 30438 29466 30490
rect 29466 30438 29478 30490
rect 29478 30438 29508 30490
rect 29532 30438 29542 30490
rect 29542 30438 29588 30490
rect 29292 30436 29348 30438
rect 29372 30436 29428 30438
rect 29452 30436 29508 30438
rect 29532 30436 29588 30438
rect 26330 28600 26386 28656
rect 28262 28464 28318 28520
rect 25502 27920 25558 27976
rect 28630 27920 28686 27976
rect 25750 27770 25806 27772
rect 25830 27770 25886 27772
rect 25910 27770 25966 27772
rect 25990 27770 26046 27772
rect 25750 27718 25796 27770
rect 25796 27718 25806 27770
rect 25830 27718 25860 27770
rect 25860 27718 25872 27770
rect 25872 27718 25886 27770
rect 25910 27718 25924 27770
rect 25924 27718 25936 27770
rect 25936 27718 25966 27770
rect 25990 27718 26000 27770
rect 26000 27718 26046 27770
rect 25750 27716 25806 27718
rect 25830 27716 25886 27718
rect 25910 27716 25966 27718
rect 25990 27716 26046 27718
rect 24766 22480 24822 22536
rect 25750 26682 25806 26684
rect 25830 26682 25886 26684
rect 25910 26682 25966 26684
rect 25990 26682 26046 26684
rect 25750 26630 25796 26682
rect 25796 26630 25806 26682
rect 25830 26630 25860 26682
rect 25860 26630 25872 26682
rect 25872 26630 25886 26682
rect 25910 26630 25924 26682
rect 25924 26630 25936 26682
rect 25936 26630 25966 26682
rect 25990 26630 26000 26682
rect 26000 26630 26046 26682
rect 25750 26628 25806 26630
rect 25830 26628 25886 26630
rect 25910 26628 25966 26630
rect 25990 26628 26046 26630
rect 25750 25594 25806 25596
rect 25830 25594 25886 25596
rect 25910 25594 25966 25596
rect 25990 25594 26046 25596
rect 25750 25542 25796 25594
rect 25796 25542 25806 25594
rect 25830 25542 25860 25594
rect 25860 25542 25872 25594
rect 25872 25542 25886 25594
rect 25910 25542 25924 25594
rect 25924 25542 25936 25594
rect 25936 25542 25966 25594
rect 25990 25542 26000 25594
rect 26000 25542 26046 25594
rect 25750 25540 25806 25542
rect 25830 25540 25886 25542
rect 25910 25540 25966 25542
rect 25990 25540 26046 25542
rect 25750 24506 25806 24508
rect 25830 24506 25886 24508
rect 25910 24506 25966 24508
rect 25990 24506 26046 24508
rect 25750 24454 25796 24506
rect 25796 24454 25806 24506
rect 25830 24454 25860 24506
rect 25860 24454 25872 24506
rect 25872 24454 25886 24506
rect 25910 24454 25924 24506
rect 25924 24454 25936 24506
rect 25936 24454 25966 24506
rect 25990 24454 26000 24506
rect 26000 24454 26046 24506
rect 25750 24452 25806 24454
rect 25830 24452 25886 24454
rect 25910 24452 25966 24454
rect 25990 24452 26046 24454
rect 25750 23418 25806 23420
rect 25830 23418 25886 23420
rect 25910 23418 25966 23420
rect 25990 23418 26046 23420
rect 25750 23366 25796 23418
rect 25796 23366 25806 23418
rect 25830 23366 25860 23418
rect 25860 23366 25872 23418
rect 25872 23366 25886 23418
rect 25910 23366 25924 23418
rect 25924 23366 25936 23418
rect 25936 23366 25966 23418
rect 25990 23366 26000 23418
rect 26000 23366 26046 23418
rect 25750 23364 25806 23366
rect 25830 23364 25886 23366
rect 25910 23364 25966 23366
rect 25990 23364 26046 23366
rect 26238 23180 26294 23216
rect 26238 23160 26240 23180
rect 26240 23160 26292 23180
rect 26292 23160 26294 23180
rect 25750 22330 25806 22332
rect 25830 22330 25886 22332
rect 25910 22330 25966 22332
rect 25990 22330 26046 22332
rect 25750 22278 25796 22330
rect 25796 22278 25806 22330
rect 25830 22278 25860 22330
rect 25860 22278 25872 22330
rect 25872 22278 25886 22330
rect 25910 22278 25924 22330
rect 25924 22278 25936 22330
rect 25936 22278 25966 22330
rect 25990 22278 26000 22330
rect 26000 22278 26046 22330
rect 25750 22276 25806 22278
rect 25830 22276 25886 22278
rect 25910 22276 25966 22278
rect 25990 22276 26046 22278
rect 25750 21242 25806 21244
rect 25830 21242 25886 21244
rect 25910 21242 25966 21244
rect 25990 21242 26046 21244
rect 25750 21190 25796 21242
rect 25796 21190 25806 21242
rect 25830 21190 25860 21242
rect 25860 21190 25872 21242
rect 25872 21190 25886 21242
rect 25910 21190 25924 21242
rect 25924 21190 25936 21242
rect 25936 21190 25966 21242
rect 25990 21190 26000 21242
rect 26000 21190 26046 21242
rect 25750 21188 25806 21190
rect 25830 21188 25886 21190
rect 25910 21188 25966 21190
rect 25990 21188 26046 21190
rect 25750 20154 25806 20156
rect 25830 20154 25886 20156
rect 25910 20154 25966 20156
rect 25990 20154 26046 20156
rect 25750 20102 25796 20154
rect 25796 20102 25806 20154
rect 25830 20102 25860 20154
rect 25860 20102 25872 20154
rect 25872 20102 25886 20154
rect 25910 20102 25924 20154
rect 25924 20102 25936 20154
rect 25936 20102 25966 20154
rect 25990 20102 26000 20154
rect 26000 20102 26046 20154
rect 25750 20100 25806 20102
rect 25830 20100 25886 20102
rect 25910 20100 25966 20102
rect 25990 20100 26046 20102
rect 25750 19066 25806 19068
rect 25830 19066 25886 19068
rect 25910 19066 25966 19068
rect 25990 19066 26046 19068
rect 25750 19014 25796 19066
rect 25796 19014 25806 19066
rect 25830 19014 25860 19066
rect 25860 19014 25872 19066
rect 25872 19014 25886 19066
rect 25910 19014 25924 19066
rect 25924 19014 25936 19066
rect 25936 19014 25966 19066
rect 25990 19014 26000 19066
rect 26000 19014 26046 19066
rect 25750 19012 25806 19014
rect 25830 19012 25886 19014
rect 25910 19012 25966 19014
rect 25990 19012 26046 19014
rect 25750 17978 25806 17980
rect 25830 17978 25886 17980
rect 25910 17978 25966 17980
rect 25990 17978 26046 17980
rect 25750 17926 25796 17978
rect 25796 17926 25806 17978
rect 25830 17926 25860 17978
rect 25860 17926 25872 17978
rect 25872 17926 25886 17978
rect 25910 17926 25924 17978
rect 25924 17926 25936 17978
rect 25936 17926 25966 17978
rect 25990 17926 26000 17978
rect 26000 17926 26046 17978
rect 25750 17924 25806 17926
rect 25830 17924 25886 17926
rect 25910 17924 25966 17926
rect 25990 17924 26046 17926
rect 25750 16890 25806 16892
rect 25830 16890 25886 16892
rect 25910 16890 25966 16892
rect 25990 16890 26046 16892
rect 25750 16838 25796 16890
rect 25796 16838 25806 16890
rect 25830 16838 25860 16890
rect 25860 16838 25872 16890
rect 25872 16838 25886 16890
rect 25910 16838 25924 16890
rect 25924 16838 25936 16890
rect 25936 16838 25966 16890
rect 25990 16838 26000 16890
rect 26000 16838 26046 16890
rect 25750 16836 25806 16838
rect 25830 16836 25886 16838
rect 25910 16836 25966 16838
rect 25990 16836 26046 16838
rect 25042 14476 25098 14512
rect 25042 14456 25044 14476
rect 25044 14456 25096 14476
rect 25096 14456 25098 14476
rect 24398 10648 24454 10704
rect 24214 10532 24270 10568
rect 24214 10512 24216 10532
rect 24216 10512 24268 10532
rect 24268 10512 24270 10532
rect 25750 15802 25806 15804
rect 25830 15802 25886 15804
rect 25910 15802 25966 15804
rect 25990 15802 26046 15804
rect 25750 15750 25796 15802
rect 25796 15750 25806 15802
rect 25830 15750 25860 15802
rect 25860 15750 25872 15802
rect 25872 15750 25886 15802
rect 25910 15750 25924 15802
rect 25924 15750 25936 15802
rect 25936 15750 25966 15802
rect 25990 15750 26000 15802
rect 26000 15750 26046 15802
rect 25750 15748 25806 15750
rect 25830 15748 25886 15750
rect 25910 15748 25966 15750
rect 25990 15748 26046 15750
rect 25750 14714 25806 14716
rect 25830 14714 25886 14716
rect 25910 14714 25966 14716
rect 25990 14714 26046 14716
rect 25750 14662 25796 14714
rect 25796 14662 25806 14714
rect 25830 14662 25860 14714
rect 25860 14662 25872 14714
rect 25872 14662 25886 14714
rect 25910 14662 25924 14714
rect 25924 14662 25936 14714
rect 25936 14662 25966 14714
rect 25990 14662 26000 14714
rect 26000 14662 26046 14714
rect 25750 14660 25806 14662
rect 25830 14660 25886 14662
rect 25910 14660 25966 14662
rect 25990 14660 26046 14662
rect 25750 13626 25806 13628
rect 25830 13626 25886 13628
rect 25910 13626 25966 13628
rect 25990 13626 26046 13628
rect 25750 13574 25796 13626
rect 25796 13574 25806 13626
rect 25830 13574 25860 13626
rect 25860 13574 25872 13626
rect 25872 13574 25886 13626
rect 25910 13574 25924 13626
rect 25924 13574 25936 13626
rect 25936 13574 25966 13626
rect 25990 13574 26000 13626
rect 26000 13574 26046 13626
rect 25750 13572 25806 13574
rect 25830 13572 25886 13574
rect 25910 13572 25966 13574
rect 25990 13572 26046 13574
rect 25750 12538 25806 12540
rect 25830 12538 25886 12540
rect 25910 12538 25966 12540
rect 25990 12538 26046 12540
rect 25750 12486 25796 12538
rect 25796 12486 25806 12538
rect 25830 12486 25860 12538
rect 25860 12486 25872 12538
rect 25872 12486 25886 12538
rect 25910 12486 25924 12538
rect 25924 12486 25936 12538
rect 25936 12486 25966 12538
rect 25990 12486 26000 12538
rect 26000 12486 26046 12538
rect 25750 12484 25806 12486
rect 25830 12484 25886 12486
rect 25910 12484 25966 12486
rect 25990 12484 26046 12486
rect 25750 11450 25806 11452
rect 25830 11450 25886 11452
rect 25910 11450 25966 11452
rect 25990 11450 26046 11452
rect 25750 11398 25796 11450
rect 25796 11398 25806 11450
rect 25830 11398 25860 11450
rect 25860 11398 25872 11450
rect 25872 11398 25886 11450
rect 25910 11398 25924 11450
rect 25924 11398 25936 11450
rect 25936 11398 25966 11450
rect 25990 11398 26000 11450
rect 26000 11398 26046 11450
rect 25750 11396 25806 11398
rect 25830 11396 25886 11398
rect 25910 11396 25966 11398
rect 25990 11396 26046 11398
rect 25502 10104 25558 10160
rect 25750 10362 25806 10364
rect 25830 10362 25886 10364
rect 25910 10362 25966 10364
rect 25990 10362 26046 10364
rect 25750 10310 25796 10362
rect 25796 10310 25806 10362
rect 25830 10310 25860 10362
rect 25860 10310 25872 10362
rect 25872 10310 25886 10362
rect 25910 10310 25924 10362
rect 25924 10310 25936 10362
rect 25936 10310 25966 10362
rect 25990 10310 26000 10362
rect 26000 10310 26046 10362
rect 25750 10308 25806 10310
rect 25830 10308 25886 10310
rect 25910 10308 25966 10310
rect 25990 10308 26046 10310
rect 25750 9274 25806 9276
rect 25830 9274 25886 9276
rect 25910 9274 25966 9276
rect 25990 9274 26046 9276
rect 25750 9222 25796 9274
rect 25796 9222 25806 9274
rect 25830 9222 25860 9274
rect 25860 9222 25872 9274
rect 25872 9222 25886 9274
rect 25910 9222 25924 9274
rect 25924 9222 25936 9274
rect 25936 9222 25966 9274
rect 25990 9222 26000 9274
rect 26000 9222 26046 9274
rect 25750 9220 25806 9222
rect 25830 9220 25886 9222
rect 25910 9220 25966 9222
rect 25990 9220 26046 9222
rect 25750 8186 25806 8188
rect 25830 8186 25886 8188
rect 25910 8186 25966 8188
rect 25990 8186 26046 8188
rect 25750 8134 25796 8186
rect 25796 8134 25806 8186
rect 25830 8134 25860 8186
rect 25860 8134 25872 8186
rect 25872 8134 25886 8186
rect 25910 8134 25924 8186
rect 25924 8134 25936 8186
rect 25936 8134 25966 8186
rect 25990 8134 26000 8186
rect 26000 8134 26046 8186
rect 25750 8132 25806 8134
rect 25830 8132 25886 8134
rect 25910 8132 25966 8134
rect 25990 8132 26046 8134
rect 26514 9560 26570 9616
rect 25750 7098 25806 7100
rect 25830 7098 25886 7100
rect 25910 7098 25966 7100
rect 25990 7098 26046 7100
rect 25750 7046 25796 7098
rect 25796 7046 25806 7098
rect 25830 7046 25860 7098
rect 25860 7046 25872 7098
rect 25872 7046 25886 7098
rect 25910 7046 25924 7098
rect 25924 7046 25936 7098
rect 25936 7046 25966 7098
rect 25990 7046 26000 7098
rect 26000 7046 26046 7098
rect 25750 7044 25806 7046
rect 25830 7044 25886 7046
rect 25910 7044 25966 7046
rect 25990 7044 26046 7046
rect 25750 6010 25806 6012
rect 25830 6010 25886 6012
rect 25910 6010 25966 6012
rect 25990 6010 26046 6012
rect 25750 5958 25796 6010
rect 25796 5958 25806 6010
rect 25830 5958 25860 6010
rect 25860 5958 25872 6010
rect 25872 5958 25886 6010
rect 25910 5958 25924 6010
rect 25924 5958 25936 6010
rect 25936 5958 25966 6010
rect 25990 5958 26000 6010
rect 26000 5958 26046 6010
rect 25750 5956 25806 5958
rect 25830 5956 25886 5958
rect 25910 5956 25966 5958
rect 25990 5956 26046 5958
rect 28262 22616 28318 22672
rect 27986 19796 27988 19816
rect 27988 19796 28040 19816
rect 28040 19796 28042 19816
rect 27986 19760 28042 19796
rect 28630 25880 28686 25936
rect 28630 23160 28686 23216
rect 28722 21120 28778 21176
rect 28722 19080 28778 19136
rect 28722 16532 28724 16552
rect 28724 16532 28776 16552
rect 28776 16532 28778 16552
rect 28722 16496 28778 16532
rect 28630 14320 28686 14376
rect 28446 13932 28502 13968
rect 28446 13912 28448 13932
rect 28448 13912 28500 13932
rect 28500 13912 28502 13932
rect 27986 12416 28042 12472
rect 27894 8880 27950 8936
rect 25750 4922 25806 4924
rect 25830 4922 25886 4924
rect 25910 4922 25966 4924
rect 25990 4922 26046 4924
rect 25750 4870 25796 4922
rect 25796 4870 25806 4922
rect 25830 4870 25860 4922
rect 25860 4870 25872 4922
rect 25872 4870 25886 4922
rect 25910 4870 25924 4922
rect 25924 4870 25936 4922
rect 25936 4870 25966 4922
rect 25990 4870 26000 4922
rect 26000 4870 26046 4922
rect 25750 4868 25806 4870
rect 25830 4868 25886 4870
rect 25910 4868 25966 4870
rect 25990 4868 26046 4870
rect 25750 3834 25806 3836
rect 25830 3834 25886 3836
rect 25910 3834 25966 3836
rect 25990 3834 26046 3836
rect 25750 3782 25796 3834
rect 25796 3782 25806 3834
rect 25830 3782 25860 3834
rect 25860 3782 25872 3834
rect 25872 3782 25886 3834
rect 25910 3782 25924 3834
rect 25924 3782 25936 3834
rect 25936 3782 25966 3834
rect 25990 3782 26000 3834
rect 26000 3782 26046 3834
rect 25750 3780 25806 3782
rect 25830 3780 25886 3782
rect 25910 3780 25966 3782
rect 25990 3780 26046 3782
rect 25750 2746 25806 2748
rect 25830 2746 25886 2748
rect 25910 2746 25966 2748
rect 25990 2746 26046 2748
rect 25750 2694 25796 2746
rect 25796 2694 25806 2746
rect 25830 2694 25860 2746
rect 25860 2694 25872 2746
rect 25872 2694 25886 2746
rect 25910 2694 25924 2746
rect 25924 2694 25936 2746
rect 25936 2694 25966 2746
rect 25990 2694 26000 2746
rect 26000 2694 26046 2746
rect 25750 2692 25806 2694
rect 25830 2692 25886 2694
rect 25910 2692 25966 2694
rect 25990 2692 26046 2694
rect 22208 2202 22264 2204
rect 22288 2202 22344 2204
rect 22368 2202 22424 2204
rect 22448 2202 22504 2204
rect 22208 2150 22254 2202
rect 22254 2150 22264 2202
rect 22288 2150 22318 2202
rect 22318 2150 22330 2202
rect 22330 2150 22344 2202
rect 22368 2150 22382 2202
rect 22382 2150 22394 2202
rect 22394 2150 22424 2202
rect 22448 2150 22458 2202
rect 22458 2150 22504 2202
rect 22208 2148 22264 2150
rect 22288 2148 22344 2150
rect 22368 2148 22424 2150
rect 22448 2148 22504 2150
rect 28354 12416 28410 12472
rect 28630 12280 28686 12336
rect 28722 9580 28778 9616
rect 28722 9560 28724 9580
rect 28724 9560 28776 9580
rect 28776 9560 28778 9580
rect 29292 29402 29348 29404
rect 29372 29402 29428 29404
rect 29452 29402 29508 29404
rect 29532 29402 29588 29404
rect 29292 29350 29338 29402
rect 29338 29350 29348 29402
rect 29372 29350 29402 29402
rect 29402 29350 29414 29402
rect 29414 29350 29428 29402
rect 29452 29350 29466 29402
rect 29466 29350 29478 29402
rect 29478 29350 29508 29402
rect 29532 29350 29542 29402
rect 29542 29350 29588 29402
rect 29292 29348 29348 29350
rect 29372 29348 29428 29350
rect 29452 29348 29508 29350
rect 29532 29348 29588 29350
rect 29292 28314 29348 28316
rect 29372 28314 29428 28316
rect 29452 28314 29508 28316
rect 29532 28314 29588 28316
rect 29292 28262 29338 28314
rect 29338 28262 29348 28314
rect 29372 28262 29402 28314
rect 29402 28262 29414 28314
rect 29414 28262 29428 28314
rect 29452 28262 29466 28314
rect 29466 28262 29478 28314
rect 29478 28262 29508 28314
rect 29532 28262 29542 28314
rect 29542 28262 29588 28314
rect 29292 28260 29348 28262
rect 29372 28260 29428 28262
rect 29452 28260 29508 28262
rect 29532 28260 29588 28262
rect 29292 27226 29348 27228
rect 29372 27226 29428 27228
rect 29452 27226 29508 27228
rect 29532 27226 29588 27228
rect 29292 27174 29338 27226
rect 29338 27174 29348 27226
rect 29372 27174 29402 27226
rect 29402 27174 29414 27226
rect 29414 27174 29428 27226
rect 29452 27174 29466 27226
rect 29466 27174 29478 27226
rect 29478 27174 29508 27226
rect 29532 27174 29542 27226
rect 29542 27174 29588 27226
rect 29292 27172 29348 27174
rect 29372 27172 29428 27174
rect 29452 27172 29508 27174
rect 29532 27172 29588 27174
rect 29292 26138 29348 26140
rect 29372 26138 29428 26140
rect 29452 26138 29508 26140
rect 29532 26138 29588 26140
rect 29292 26086 29338 26138
rect 29338 26086 29348 26138
rect 29372 26086 29402 26138
rect 29402 26086 29414 26138
rect 29414 26086 29428 26138
rect 29452 26086 29466 26138
rect 29466 26086 29478 26138
rect 29478 26086 29508 26138
rect 29532 26086 29542 26138
rect 29542 26086 29588 26138
rect 29292 26084 29348 26086
rect 29372 26084 29428 26086
rect 29452 26084 29508 26086
rect 29532 26084 29588 26086
rect 29292 25050 29348 25052
rect 29372 25050 29428 25052
rect 29452 25050 29508 25052
rect 29532 25050 29588 25052
rect 29292 24998 29338 25050
rect 29338 24998 29348 25050
rect 29372 24998 29402 25050
rect 29402 24998 29414 25050
rect 29414 24998 29428 25050
rect 29452 24998 29466 25050
rect 29466 24998 29478 25050
rect 29478 24998 29508 25050
rect 29532 24998 29542 25050
rect 29542 24998 29588 25050
rect 29292 24996 29348 24998
rect 29372 24996 29428 24998
rect 29452 24996 29508 24998
rect 29532 24996 29588 24998
rect 29292 23962 29348 23964
rect 29372 23962 29428 23964
rect 29452 23962 29508 23964
rect 29532 23962 29588 23964
rect 29292 23910 29338 23962
rect 29338 23910 29348 23962
rect 29372 23910 29402 23962
rect 29402 23910 29414 23962
rect 29414 23910 29428 23962
rect 29452 23910 29466 23962
rect 29466 23910 29478 23962
rect 29478 23910 29508 23962
rect 29532 23910 29542 23962
rect 29542 23910 29588 23962
rect 29292 23908 29348 23910
rect 29372 23908 29428 23910
rect 29452 23908 29508 23910
rect 29532 23908 29588 23910
rect 29292 22874 29348 22876
rect 29372 22874 29428 22876
rect 29452 22874 29508 22876
rect 29532 22874 29588 22876
rect 29292 22822 29338 22874
rect 29338 22822 29348 22874
rect 29372 22822 29402 22874
rect 29402 22822 29414 22874
rect 29414 22822 29428 22874
rect 29452 22822 29466 22874
rect 29466 22822 29478 22874
rect 29478 22822 29508 22874
rect 29532 22822 29542 22874
rect 29542 22822 29588 22874
rect 29292 22820 29348 22822
rect 29372 22820 29428 22822
rect 29452 22820 29508 22822
rect 29532 22820 29588 22822
rect 29292 21786 29348 21788
rect 29372 21786 29428 21788
rect 29452 21786 29508 21788
rect 29532 21786 29588 21788
rect 29292 21734 29338 21786
rect 29338 21734 29348 21786
rect 29372 21734 29402 21786
rect 29402 21734 29414 21786
rect 29414 21734 29428 21786
rect 29452 21734 29466 21786
rect 29466 21734 29478 21786
rect 29478 21734 29508 21786
rect 29532 21734 29542 21786
rect 29542 21734 29588 21786
rect 29292 21732 29348 21734
rect 29372 21732 29428 21734
rect 29452 21732 29508 21734
rect 29532 21732 29588 21734
rect 29292 20698 29348 20700
rect 29372 20698 29428 20700
rect 29452 20698 29508 20700
rect 29532 20698 29588 20700
rect 29292 20646 29338 20698
rect 29338 20646 29348 20698
rect 29372 20646 29402 20698
rect 29402 20646 29414 20698
rect 29414 20646 29428 20698
rect 29452 20646 29466 20698
rect 29466 20646 29478 20698
rect 29478 20646 29508 20698
rect 29532 20646 29542 20698
rect 29542 20646 29588 20698
rect 29292 20644 29348 20646
rect 29372 20644 29428 20646
rect 29452 20644 29508 20646
rect 29532 20644 29588 20646
rect 29292 19610 29348 19612
rect 29372 19610 29428 19612
rect 29452 19610 29508 19612
rect 29532 19610 29588 19612
rect 29292 19558 29338 19610
rect 29338 19558 29348 19610
rect 29372 19558 29402 19610
rect 29402 19558 29414 19610
rect 29414 19558 29428 19610
rect 29452 19558 29466 19610
rect 29466 19558 29478 19610
rect 29478 19558 29508 19610
rect 29532 19558 29542 19610
rect 29542 19558 29588 19610
rect 29292 19556 29348 19558
rect 29372 19556 29428 19558
rect 29452 19556 29508 19558
rect 29532 19556 29588 19558
rect 29292 18522 29348 18524
rect 29372 18522 29428 18524
rect 29452 18522 29508 18524
rect 29532 18522 29588 18524
rect 29292 18470 29338 18522
rect 29338 18470 29348 18522
rect 29372 18470 29402 18522
rect 29402 18470 29414 18522
rect 29414 18470 29428 18522
rect 29452 18470 29466 18522
rect 29466 18470 29478 18522
rect 29478 18470 29508 18522
rect 29532 18470 29542 18522
rect 29542 18470 29588 18522
rect 29292 18468 29348 18470
rect 29372 18468 29428 18470
rect 29452 18468 29508 18470
rect 29532 18468 29588 18470
rect 29292 17434 29348 17436
rect 29372 17434 29428 17436
rect 29452 17434 29508 17436
rect 29532 17434 29588 17436
rect 29292 17382 29338 17434
rect 29338 17382 29348 17434
rect 29372 17382 29402 17434
rect 29402 17382 29414 17434
rect 29414 17382 29428 17434
rect 29452 17382 29466 17434
rect 29466 17382 29478 17434
rect 29478 17382 29508 17434
rect 29532 17382 29542 17434
rect 29542 17382 29588 17434
rect 29292 17380 29348 17382
rect 29372 17380 29428 17382
rect 29452 17380 29508 17382
rect 29532 17380 29588 17382
rect 29292 16346 29348 16348
rect 29372 16346 29428 16348
rect 29452 16346 29508 16348
rect 29532 16346 29588 16348
rect 29292 16294 29338 16346
rect 29338 16294 29348 16346
rect 29372 16294 29402 16346
rect 29402 16294 29414 16346
rect 29414 16294 29428 16346
rect 29452 16294 29466 16346
rect 29466 16294 29478 16346
rect 29478 16294 29508 16346
rect 29532 16294 29542 16346
rect 29542 16294 29588 16346
rect 29292 16292 29348 16294
rect 29372 16292 29428 16294
rect 29452 16292 29508 16294
rect 29532 16292 29588 16294
rect 29292 15258 29348 15260
rect 29372 15258 29428 15260
rect 29452 15258 29508 15260
rect 29532 15258 29588 15260
rect 29292 15206 29338 15258
rect 29338 15206 29348 15258
rect 29372 15206 29402 15258
rect 29402 15206 29414 15258
rect 29414 15206 29428 15258
rect 29452 15206 29466 15258
rect 29466 15206 29478 15258
rect 29478 15206 29508 15258
rect 29532 15206 29542 15258
rect 29542 15206 29588 15258
rect 29292 15204 29348 15206
rect 29372 15204 29428 15206
rect 29452 15204 29508 15206
rect 29532 15204 29588 15206
rect 29292 14170 29348 14172
rect 29372 14170 29428 14172
rect 29452 14170 29508 14172
rect 29532 14170 29588 14172
rect 29292 14118 29338 14170
rect 29338 14118 29348 14170
rect 29372 14118 29402 14170
rect 29402 14118 29414 14170
rect 29414 14118 29428 14170
rect 29452 14118 29466 14170
rect 29466 14118 29478 14170
rect 29478 14118 29508 14170
rect 29532 14118 29542 14170
rect 29542 14118 29588 14170
rect 29292 14116 29348 14118
rect 29372 14116 29428 14118
rect 29452 14116 29508 14118
rect 29532 14116 29588 14118
rect 29292 13082 29348 13084
rect 29372 13082 29428 13084
rect 29452 13082 29508 13084
rect 29532 13082 29588 13084
rect 29292 13030 29338 13082
rect 29338 13030 29348 13082
rect 29372 13030 29402 13082
rect 29402 13030 29414 13082
rect 29414 13030 29428 13082
rect 29452 13030 29466 13082
rect 29466 13030 29478 13082
rect 29478 13030 29508 13082
rect 29532 13030 29542 13082
rect 29542 13030 29588 13082
rect 29292 13028 29348 13030
rect 29372 13028 29428 13030
rect 29452 13028 29508 13030
rect 29532 13028 29588 13030
rect 29292 11994 29348 11996
rect 29372 11994 29428 11996
rect 29452 11994 29508 11996
rect 29532 11994 29588 11996
rect 29292 11942 29338 11994
rect 29338 11942 29348 11994
rect 29372 11942 29402 11994
rect 29402 11942 29414 11994
rect 29414 11942 29428 11994
rect 29452 11942 29466 11994
rect 29466 11942 29478 11994
rect 29478 11942 29508 11994
rect 29532 11942 29542 11994
rect 29542 11942 29588 11994
rect 29292 11940 29348 11942
rect 29372 11940 29428 11942
rect 29452 11940 29508 11942
rect 29532 11940 29588 11942
rect 29292 10906 29348 10908
rect 29372 10906 29428 10908
rect 29452 10906 29508 10908
rect 29532 10906 29588 10908
rect 29292 10854 29338 10906
rect 29338 10854 29348 10906
rect 29372 10854 29402 10906
rect 29402 10854 29414 10906
rect 29414 10854 29428 10906
rect 29452 10854 29466 10906
rect 29466 10854 29478 10906
rect 29478 10854 29508 10906
rect 29532 10854 29542 10906
rect 29542 10854 29588 10906
rect 29292 10852 29348 10854
rect 29372 10852 29428 10854
rect 29452 10852 29508 10854
rect 29532 10852 29588 10854
rect 29292 9818 29348 9820
rect 29372 9818 29428 9820
rect 29452 9818 29508 9820
rect 29532 9818 29588 9820
rect 29292 9766 29338 9818
rect 29338 9766 29348 9818
rect 29372 9766 29402 9818
rect 29402 9766 29414 9818
rect 29414 9766 29428 9818
rect 29452 9766 29466 9818
rect 29466 9766 29478 9818
rect 29478 9766 29508 9818
rect 29532 9766 29542 9818
rect 29542 9766 29588 9818
rect 29292 9764 29348 9766
rect 29372 9764 29428 9766
rect 29452 9764 29508 9766
rect 29532 9764 29588 9766
rect 29292 8730 29348 8732
rect 29372 8730 29428 8732
rect 29452 8730 29508 8732
rect 29532 8730 29588 8732
rect 29292 8678 29338 8730
rect 29338 8678 29348 8730
rect 29372 8678 29402 8730
rect 29402 8678 29414 8730
rect 29414 8678 29428 8730
rect 29452 8678 29466 8730
rect 29466 8678 29478 8730
rect 29478 8678 29508 8730
rect 29532 8678 29542 8730
rect 29542 8678 29588 8730
rect 29292 8676 29348 8678
rect 29372 8676 29428 8678
rect 29452 8676 29508 8678
rect 29532 8676 29588 8678
rect 29292 7642 29348 7644
rect 29372 7642 29428 7644
rect 29452 7642 29508 7644
rect 29532 7642 29588 7644
rect 29292 7590 29338 7642
rect 29338 7590 29348 7642
rect 29372 7590 29402 7642
rect 29402 7590 29414 7642
rect 29414 7590 29428 7642
rect 29452 7590 29466 7642
rect 29466 7590 29478 7642
rect 29478 7590 29508 7642
rect 29532 7590 29542 7642
rect 29542 7590 29588 7642
rect 29292 7588 29348 7590
rect 29372 7588 29428 7590
rect 29452 7588 29508 7590
rect 29532 7588 29588 7590
rect 28722 7420 28724 7440
rect 28724 7420 28776 7440
rect 28776 7420 28778 7440
rect 28722 7384 28778 7420
rect 29292 6554 29348 6556
rect 29372 6554 29428 6556
rect 29452 6554 29508 6556
rect 29532 6554 29588 6556
rect 29292 6502 29338 6554
rect 29338 6502 29348 6554
rect 29372 6502 29402 6554
rect 29402 6502 29414 6554
rect 29414 6502 29428 6554
rect 29452 6502 29466 6554
rect 29466 6502 29478 6554
rect 29478 6502 29508 6554
rect 29532 6502 29542 6554
rect 29542 6502 29588 6554
rect 29292 6500 29348 6502
rect 29372 6500 29428 6502
rect 29452 6500 29508 6502
rect 29532 6500 29588 6502
rect 29292 5466 29348 5468
rect 29372 5466 29428 5468
rect 29452 5466 29508 5468
rect 29532 5466 29588 5468
rect 29292 5414 29338 5466
rect 29338 5414 29348 5466
rect 29372 5414 29402 5466
rect 29402 5414 29414 5466
rect 29414 5414 29428 5466
rect 29452 5414 29466 5466
rect 29466 5414 29478 5466
rect 29478 5414 29508 5466
rect 29532 5414 29542 5466
rect 29542 5414 29588 5466
rect 29292 5412 29348 5414
rect 29372 5412 29428 5414
rect 29452 5412 29508 5414
rect 29532 5412 29588 5414
rect 28722 5208 28778 5264
rect 29292 4378 29348 4380
rect 29372 4378 29428 4380
rect 29452 4378 29508 4380
rect 29532 4378 29588 4380
rect 29292 4326 29338 4378
rect 29338 4326 29348 4378
rect 29372 4326 29402 4378
rect 29402 4326 29414 4378
rect 29414 4326 29428 4378
rect 29452 4326 29466 4378
rect 29466 4326 29478 4378
rect 29478 4326 29508 4378
rect 29532 4326 29542 4378
rect 29542 4326 29588 4378
rect 29292 4324 29348 4326
rect 29372 4324 29428 4326
rect 29452 4324 29508 4326
rect 29532 4324 29588 4326
rect 29292 3290 29348 3292
rect 29372 3290 29428 3292
rect 29452 3290 29508 3292
rect 29532 3290 29588 3292
rect 29292 3238 29338 3290
rect 29338 3238 29348 3290
rect 29372 3238 29402 3290
rect 29402 3238 29414 3290
rect 29414 3238 29428 3290
rect 29452 3238 29466 3290
rect 29466 3238 29478 3290
rect 29478 3238 29508 3290
rect 29532 3238 29542 3290
rect 29542 3238 29588 3290
rect 29292 3236 29348 3238
rect 29372 3236 29428 3238
rect 29452 3236 29508 3238
rect 29532 3236 29588 3238
rect 28630 2760 28686 2816
rect 29292 2202 29348 2204
rect 29372 2202 29428 2204
rect 29452 2202 29508 2204
rect 29532 2202 29588 2204
rect 29292 2150 29338 2202
rect 29338 2150 29348 2202
rect 29372 2150 29402 2202
rect 29402 2150 29414 2202
rect 29414 2150 29428 2202
rect 29452 2150 29466 2202
rect 29466 2150 29478 2202
rect 29478 2150 29508 2202
rect 29532 2150 29542 2202
rect 29542 2150 29588 2202
rect 29292 2148 29348 2150
rect 29372 2148 29428 2150
rect 29452 2148 29508 2150
rect 29532 2148 29588 2150
rect 27434 720 27490 776
<< metal3 >>
rect 0 31378 800 31408
rect 1853 31378 1919 31381
rect 0 31376 1919 31378
rect 0 31320 1858 31376
rect 1914 31320 1919 31376
rect 0 31318 1919 31320
rect 0 31288 800 31318
rect 1853 31315 1919 31318
rect 8030 30496 8346 30497
rect 8030 30432 8036 30496
rect 8100 30432 8116 30496
rect 8180 30432 8196 30496
rect 8260 30432 8276 30496
rect 8340 30432 8346 30496
rect 8030 30431 8346 30432
rect 15114 30496 15430 30497
rect 15114 30432 15120 30496
rect 15184 30432 15200 30496
rect 15264 30432 15280 30496
rect 15344 30432 15360 30496
rect 15424 30432 15430 30496
rect 15114 30431 15430 30432
rect 22198 30496 22514 30497
rect 22198 30432 22204 30496
rect 22268 30432 22284 30496
rect 22348 30432 22364 30496
rect 22428 30432 22444 30496
rect 22508 30432 22514 30496
rect 22198 30431 22514 30432
rect 29282 30496 29598 30497
rect 29282 30432 29288 30496
rect 29352 30432 29368 30496
rect 29432 30432 29448 30496
rect 29512 30432 29528 30496
rect 29592 30432 29598 30496
rect 29282 30431 29598 30432
rect 27889 30018 27955 30021
rect 29821 30018 30621 30048
rect 27889 30016 30621 30018
rect 27889 29960 27894 30016
rect 27950 29960 30621 30016
rect 27889 29958 30621 29960
rect 27889 29955 27955 29958
rect 4488 29952 4804 29953
rect 4488 29888 4494 29952
rect 4558 29888 4574 29952
rect 4638 29888 4654 29952
rect 4718 29888 4734 29952
rect 4798 29888 4804 29952
rect 4488 29887 4804 29888
rect 11572 29952 11888 29953
rect 11572 29888 11578 29952
rect 11642 29888 11658 29952
rect 11722 29888 11738 29952
rect 11802 29888 11818 29952
rect 11882 29888 11888 29952
rect 11572 29887 11888 29888
rect 18656 29952 18972 29953
rect 18656 29888 18662 29952
rect 18726 29888 18742 29952
rect 18806 29888 18822 29952
rect 18886 29888 18902 29952
rect 18966 29888 18972 29952
rect 18656 29887 18972 29888
rect 25740 29952 26056 29953
rect 25740 29888 25746 29952
rect 25810 29888 25826 29952
rect 25890 29888 25906 29952
rect 25970 29888 25986 29952
rect 26050 29888 26056 29952
rect 29821 29928 30621 29958
rect 25740 29887 26056 29888
rect 8030 29408 8346 29409
rect 0 29338 800 29368
rect 8030 29344 8036 29408
rect 8100 29344 8116 29408
rect 8180 29344 8196 29408
rect 8260 29344 8276 29408
rect 8340 29344 8346 29408
rect 8030 29343 8346 29344
rect 15114 29408 15430 29409
rect 15114 29344 15120 29408
rect 15184 29344 15200 29408
rect 15264 29344 15280 29408
rect 15344 29344 15360 29408
rect 15424 29344 15430 29408
rect 15114 29343 15430 29344
rect 22198 29408 22514 29409
rect 22198 29344 22204 29408
rect 22268 29344 22284 29408
rect 22348 29344 22364 29408
rect 22428 29344 22444 29408
rect 22508 29344 22514 29408
rect 22198 29343 22514 29344
rect 29282 29408 29598 29409
rect 29282 29344 29288 29408
rect 29352 29344 29368 29408
rect 29432 29344 29448 29408
rect 29512 29344 29528 29408
rect 29592 29344 29598 29408
rect 29282 29343 29598 29344
rect 1485 29338 1551 29341
rect 0 29336 1551 29338
rect 0 29280 1490 29336
rect 1546 29280 1551 29336
rect 0 29278 1551 29280
rect 0 29248 800 29278
rect 1485 29275 1551 29278
rect 27613 29338 27679 29341
rect 27838 29338 27844 29340
rect 27613 29336 27844 29338
rect 27613 29280 27618 29336
rect 27674 29280 27844 29336
rect 27613 29278 27844 29280
rect 27613 29275 27679 29278
rect 27838 29276 27844 29278
rect 27908 29276 27914 29340
rect 4488 28864 4804 28865
rect 4488 28800 4494 28864
rect 4558 28800 4574 28864
rect 4638 28800 4654 28864
rect 4718 28800 4734 28864
rect 4798 28800 4804 28864
rect 4488 28799 4804 28800
rect 11572 28864 11888 28865
rect 11572 28800 11578 28864
rect 11642 28800 11658 28864
rect 11722 28800 11738 28864
rect 11802 28800 11818 28864
rect 11882 28800 11888 28864
rect 11572 28799 11888 28800
rect 18656 28864 18972 28865
rect 18656 28800 18662 28864
rect 18726 28800 18742 28864
rect 18806 28800 18822 28864
rect 18886 28800 18902 28864
rect 18966 28800 18972 28864
rect 18656 28799 18972 28800
rect 25740 28864 26056 28865
rect 25740 28800 25746 28864
rect 25810 28800 25826 28864
rect 25890 28800 25906 28864
rect 25970 28800 25986 28864
rect 26050 28800 26056 28864
rect 25740 28799 26056 28800
rect 14825 28658 14891 28661
rect 26325 28658 26391 28661
rect 14825 28656 26391 28658
rect 14825 28600 14830 28656
rect 14886 28600 26330 28656
rect 26386 28600 26391 28656
rect 14825 28598 26391 28600
rect 14825 28595 14891 28598
rect 26325 28595 26391 28598
rect 16205 28522 16271 28525
rect 28257 28522 28323 28525
rect 16205 28520 28323 28522
rect 16205 28464 16210 28520
rect 16266 28464 28262 28520
rect 28318 28464 28323 28520
rect 16205 28462 28323 28464
rect 16205 28459 16271 28462
rect 28257 28459 28323 28462
rect 8030 28320 8346 28321
rect 8030 28256 8036 28320
rect 8100 28256 8116 28320
rect 8180 28256 8196 28320
rect 8260 28256 8276 28320
rect 8340 28256 8346 28320
rect 8030 28255 8346 28256
rect 15114 28320 15430 28321
rect 15114 28256 15120 28320
rect 15184 28256 15200 28320
rect 15264 28256 15280 28320
rect 15344 28256 15360 28320
rect 15424 28256 15430 28320
rect 15114 28255 15430 28256
rect 22198 28320 22514 28321
rect 22198 28256 22204 28320
rect 22268 28256 22284 28320
rect 22348 28256 22364 28320
rect 22428 28256 22444 28320
rect 22508 28256 22514 28320
rect 22198 28255 22514 28256
rect 29282 28320 29598 28321
rect 29282 28256 29288 28320
rect 29352 28256 29368 28320
rect 29432 28256 29448 28320
rect 29512 28256 29528 28320
rect 29592 28256 29598 28320
rect 29282 28255 29598 28256
rect 16665 27978 16731 27981
rect 25497 27978 25563 27981
rect 16665 27976 25563 27978
rect 16665 27920 16670 27976
rect 16726 27920 25502 27976
rect 25558 27920 25563 27976
rect 16665 27918 25563 27920
rect 16665 27915 16731 27918
rect 25497 27915 25563 27918
rect 28625 27978 28691 27981
rect 29821 27978 30621 28008
rect 28625 27976 30621 27978
rect 28625 27920 28630 27976
rect 28686 27920 30621 27976
rect 28625 27918 30621 27920
rect 28625 27915 28691 27918
rect 29821 27888 30621 27918
rect 4488 27776 4804 27777
rect 4488 27712 4494 27776
rect 4558 27712 4574 27776
rect 4638 27712 4654 27776
rect 4718 27712 4734 27776
rect 4798 27712 4804 27776
rect 4488 27711 4804 27712
rect 11572 27776 11888 27777
rect 11572 27712 11578 27776
rect 11642 27712 11658 27776
rect 11722 27712 11738 27776
rect 11802 27712 11818 27776
rect 11882 27712 11888 27776
rect 11572 27711 11888 27712
rect 18656 27776 18972 27777
rect 18656 27712 18662 27776
rect 18726 27712 18742 27776
rect 18806 27712 18822 27776
rect 18886 27712 18902 27776
rect 18966 27712 18972 27776
rect 18656 27711 18972 27712
rect 25740 27776 26056 27777
rect 25740 27712 25746 27776
rect 25810 27712 25826 27776
rect 25890 27712 25906 27776
rect 25970 27712 25986 27776
rect 26050 27712 26056 27776
rect 25740 27711 26056 27712
rect 8030 27232 8346 27233
rect 8030 27168 8036 27232
rect 8100 27168 8116 27232
rect 8180 27168 8196 27232
rect 8260 27168 8276 27232
rect 8340 27168 8346 27232
rect 8030 27167 8346 27168
rect 15114 27232 15430 27233
rect 15114 27168 15120 27232
rect 15184 27168 15200 27232
rect 15264 27168 15280 27232
rect 15344 27168 15360 27232
rect 15424 27168 15430 27232
rect 15114 27167 15430 27168
rect 22198 27232 22514 27233
rect 22198 27168 22204 27232
rect 22268 27168 22284 27232
rect 22348 27168 22364 27232
rect 22428 27168 22444 27232
rect 22508 27168 22514 27232
rect 22198 27167 22514 27168
rect 29282 27232 29598 27233
rect 29282 27168 29288 27232
rect 29352 27168 29368 27232
rect 29432 27168 29448 27232
rect 29512 27168 29528 27232
rect 29592 27168 29598 27232
rect 29282 27167 29598 27168
rect 19885 27026 19951 27029
rect 20161 27026 20227 27029
rect 19885 27024 20227 27026
rect 19885 26968 19890 27024
rect 19946 26968 20166 27024
rect 20222 26968 20227 27024
rect 19885 26966 20227 26968
rect 19885 26963 19951 26966
rect 20161 26963 20227 26966
rect 4488 26688 4804 26689
rect 0 26618 800 26648
rect 4488 26624 4494 26688
rect 4558 26624 4574 26688
rect 4638 26624 4654 26688
rect 4718 26624 4734 26688
rect 4798 26624 4804 26688
rect 4488 26623 4804 26624
rect 11572 26688 11888 26689
rect 11572 26624 11578 26688
rect 11642 26624 11658 26688
rect 11722 26624 11738 26688
rect 11802 26624 11818 26688
rect 11882 26624 11888 26688
rect 11572 26623 11888 26624
rect 18656 26688 18972 26689
rect 18656 26624 18662 26688
rect 18726 26624 18742 26688
rect 18806 26624 18822 26688
rect 18886 26624 18902 26688
rect 18966 26624 18972 26688
rect 18656 26623 18972 26624
rect 25740 26688 26056 26689
rect 25740 26624 25746 26688
rect 25810 26624 25826 26688
rect 25890 26624 25906 26688
rect 25970 26624 25986 26688
rect 26050 26624 26056 26688
rect 25740 26623 26056 26624
rect 1577 26618 1643 26621
rect 0 26616 1643 26618
rect 0 26560 1582 26616
rect 1638 26560 1643 26616
rect 0 26558 1643 26560
rect 0 26528 800 26558
rect 1577 26555 1643 26558
rect 5349 26482 5415 26485
rect 22645 26482 22711 26485
rect 5349 26480 22711 26482
rect 5349 26424 5354 26480
rect 5410 26424 22650 26480
rect 22706 26424 22711 26480
rect 5349 26422 22711 26424
rect 5349 26419 5415 26422
rect 22645 26419 22711 26422
rect 8293 26346 8359 26349
rect 16941 26346 17007 26349
rect 18045 26346 18111 26349
rect 22553 26346 22619 26349
rect 22686 26346 22692 26348
rect 8293 26344 22692 26346
rect 8293 26288 8298 26344
rect 8354 26288 16946 26344
rect 17002 26288 18050 26344
rect 18106 26288 22558 26344
rect 22614 26288 22692 26344
rect 8293 26286 22692 26288
rect 8293 26283 8359 26286
rect 16941 26283 17007 26286
rect 18045 26283 18111 26286
rect 22553 26283 22619 26286
rect 22686 26284 22692 26286
rect 22756 26284 22762 26348
rect 8030 26144 8346 26145
rect 8030 26080 8036 26144
rect 8100 26080 8116 26144
rect 8180 26080 8196 26144
rect 8260 26080 8276 26144
rect 8340 26080 8346 26144
rect 8030 26079 8346 26080
rect 15114 26144 15430 26145
rect 15114 26080 15120 26144
rect 15184 26080 15200 26144
rect 15264 26080 15280 26144
rect 15344 26080 15360 26144
rect 15424 26080 15430 26144
rect 15114 26079 15430 26080
rect 22198 26144 22514 26145
rect 22198 26080 22204 26144
rect 22268 26080 22284 26144
rect 22348 26080 22364 26144
rect 22428 26080 22444 26144
rect 22508 26080 22514 26144
rect 22198 26079 22514 26080
rect 29282 26144 29598 26145
rect 29282 26080 29288 26144
rect 29352 26080 29368 26144
rect 29432 26080 29448 26144
rect 29512 26080 29528 26144
rect 29592 26080 29598 26144
rect 29282 26079 29598 26080
rect 10409 25938 10475 25941
rect 11973 25938 12039 25941
rect 15837 25938 15903 25941
rect 10409 25936 15903 25938
rect 10409 25880 10414 25936
rect 10470 25880 11978 25936
rect 12034 25880 15842 25936
rect 15898 25880 15903 25936
rect 10409 25878 15903 25880
rect 10409 25875 10475 25878
rect 11973 25875 12039 25878
rect 15837 25875 15903 25878
rect 28625 25938 28691 25941
rect 29821 25938 30621 25968
rect 28625 25936 30621 25938
rect 28625 25880 28630 25936
rect 28686 25880 30621 25936
rect 28625 25878 30621 25880
rect 28625 25875 28691 25878
rect 29821 25848 30621 25878
rect 4488 25600 4804 25601
rect 4488 25536 4494 25600
rect 4558 25536 4574 25600
rect 4638 25536 4654 25600
rect 4718 25536 4734 25600
rect 4798 25536 4804 25600
rect 4488 25535 4804 25536
rect 11572 25600 11888 25601
rect 11572 25536 11578 25600
rect 11642 25536 11658 25600
rect 11722 25536 11738 25600
rect 11802 25536 11818 25600
rect 11882 25536 11888 25600
rect 11572 25535 11888 25536
rect 18656 25600 18972 25601
rect 18656 25536 18662 25600
rect 18726 25536 18742 25600
rect 18806 25536 18822 25600
rect 18886 25536 18902 25600
rect 18966 25536 18972 25600
rect 18656 25535 18972 25536
rect 25740 25600 26056 25601
rect 25740 25536 25746 25600
rect 25810 25536 25826 25600
rect 25890 25536 25906 25600
rect 25970 25536 25986 25600
rect 26050 25536 26056 25600
rect 25740 25535 26056 25536
rect 8030 25056 8346 25057
rect 8030 24992 8036 25056
rect 8100 24992 8116 25056
rect 8180 24992 8196 25056
rect 8260 24992 8276 25056
rect 8340 24992 8346 25056
rect 8030 24991 8346 24992
rect 15114 25056 15430 25057
rect 15114 24992 15120 25056
rect 15184 24992 15200 25056
rect 15264 24992 15280 25056
rect 15344 24992 15360 25056
rect 15424 24992 15430 25056
rect 15114 24991 15430 24992
rect 22198 25056 22514 25057
rect 22198 24992 22204 25056
rect 22268 24992 22284 25056
rect 22348 24992 22364 25056
rect 22428 24992 22444 25056
rect 22508 24992 22514 25056
rect 22198 24991 22514 24992
rect 29282 25056 29598 25057
rect 29282 24992 29288 25056
rect 29352 24992 29368 25056
rect 29432 24992 29448 25056
rect 29512 24992 29528 25056
rect 29592 24992 29598 25056
rect 29282 24991 29598 24992
rect 0 24578 800 24608
rect 1393 24578 1459 24581
rect 0 24576 1459 24578
rect 0 24520 1398 24576
rect 1454 24520 1459 24576
rect 0 24518 1459 24520
rect 0 24488 800 24518
rect 1393 24515 1459 24518
rect 4488 24512 4804 24513
rect 4488 24448 4494 24512
rect 4558 24448 4574 24512
rect 4638 24448 4654 24512
rect 4718 24448 4734 24512
rect 4798 24448 4804 24512
rect 4488 24447 4804 24448
rect 11572 24512 11888 24513
rect 11572 24448 11578 24512
rect 11642 24448 11658 24512
rect 11722 24448 11738 24512
rect 11802 24448 11818 24512
rect 11882 24448 11888 24512
rect 11572 24447 11888 24448
rect 18656 24512 18972 24513
rect 18656 24448 18662 24512
rect 18726 24448 18742 24512
rect 18806 24448 18822 24512
rect 18886 24448 18902 24512
rect 18966 24448 18972 24512
rect 18656 24447 18972 24448
rect 25740 24512 26056 24513
rect 25740 24448 25746 24512
rect 25810 24448 25826 24512
rect 25890 24448 25906 24512
rect 25970 24448 25986 24512
rect 26050 24448 26056 24512
rect 25740 24447 26056 24448
rect 8030 23968 8346 23969
rect 8030 23904 8036 23968
rect 8100 23904 8116 23968
rect 8180 23904 8196 23968
rect 8260 23904 8276 23968
rect 8340 23904 8346 23968
rect 8030 23903 8346 23904
rect 15114 23968 15430 23969
rect 15114 23904 15120 23968
rect 15184 23904 15200 23968
rect 15264 23904 15280 23968
rect 15344 23904 15360 23968
rect 15424 23904 15430 23968
rect 15114 23903 15430 23904
rect 22198 23968 22514 23969
rect 22198 23904 22204 23968
rect 22268 23904 22284 23968
rect 22348 23904 22364 23968
rect 22428 23904 22444 23968
rect 22508 23904 22514 23968
rect 22198 23903 22514 23904
rect 29282 23968 29598 23969
rect 29282 23904 29288 23968
rect 29352 23904 29368 23968
rect 29432 23904 29448 23968
rect 29512 23904 29528 23968
rect 29592 23904 29598 23968
rect 29282 23903 29598 23904
rect 4488 23424 4804 23425
rect 4488 23360 4494 23424
rect 4558 23360 4574 23424
rect 4638 23360 4654 23424
rect 4718 23360 4734 23424
rect 4798 23360 4804 23424
rect 4488 23359 4804 23360
rect 11572 23424 11888 23425
rect 11572 23360 11578 23424
rect 11642 23360 11658 23424
rect 11722 23360 11738 23424
rect 11802 23360 11818 23424
rect 11882 23360 11888 23424
rect 11572 23359 11888 23360
rect 18656 23424 18972 23425
rect 18656 23360 18662 23424
rect 18726 23360 18742 23424
rect 18806 23360 18822 23424
rect 18886 23360 18902 23424
rect 18966 23360 18972 23424
rect 18656 23359 18972 23360
rect 25740 23424 26056 23425
rect 25740 23360 25746 23424
rect 25810 23360 25826 23424
rect 25890 23360 25906 23424
rect 25970 23360 25986 23424
rect 26050 23360 26056 23424
rect 25740 23359 26056 23360
rect 16297 23218 16363 23221
rect 26233 23218 26299 23221
rect 16297 23216 26299 23218
rect 16297 23160 16302 23216
rect 16358 23160 26238 23216
rect 26294 23160 26299 23216
rect 16297 23158 26299 23160
rect 16297 23155 16363 23158
rect 26233 23155 26299 23158
rect 28625 23218 28691 23221
rect 29821 23218 30621 23248
rect 28625 23216 30621 23218
rect 28625 23160 28630 23216
rect 28686 23160 30621 23216
rect 28625 23158 30621 23160
rect 28625 23155 28691 23158
rect 29821 23128 30621 23158
rect 21081 22948 21147 22949
rect 21030 22884 21036 22948
rect 21100 22946 21147 22948
rect 21100 22944 21192 22946
rect 21142 22888 21192 22944
rect 21100 22886 21192 22888
rect 21100 22884 21147 22886
rect 21081 22883 21147 22884
rect 8030 22880 8346 22881
rect 8030 22816 8036 22880
rect 8100 22816 8116 22880
rect 8180 22816 8196 22880
rect 8260 22816 8276 22880
rect 8340 22816 8346 22880
rect 8030 22815 8346 22816
rect 15114 22880 15430 22881
rect 15114 22816 15120 22880
rect 15184 22816 15200 22880
rect 15264 22816 15280 22880
rect 15344 22816 15360 22880
rect 15424 22816 15430 22880
rect 15114 22815 15430 22816
rect 22198 22880 22514 22881
rect 22198 22816 22204 22880
rect 22268 22816 22284 22880
rect 22348 22816 22364 22880
rect 22428 22816 22444 22880
rect 22508 22816 22514 22880
rect 22198 22815 22514 22816
rect 29282 22880 29598 22881
rect 29282 22816 29288 22880
rect 29352 22816 29368 22880
rect 29432 22816 29448 22880
rect 29512 22816 29528 22880
rect 29592 22816 29598 22880
rect 29282 22815 29598 22816
rect 3325 22674 3391 22677
rect 28257 22674 28323 22677
rect 3325 22672 28323 22674
rect 3325 22616 3330 22672
rect 3386 22616 28262 22672
rect 28318 22616 28323 22672
rect 3325 22614 28323 22616
rect 3325 22611 3391 22614
rect 28257 22611 28323 22614
rect 0 22538 800 22568
rect 1577 22538 1643 22541
rect 0 22536 1643 22538
rect 0 22480 1582 22536
rect 1638 22480 1643 22536
rect 0 22478 1643 22480
rect 0 22448 800 22478
rect 1577 22475 1643 22478
rect 1761 22538 1827 22541
rect 24761 22538 24827 22541
rect 1761 22536 24827 22538
rect 1761 22480 1766 22536
rect 1822 22480 24766 22536
rect 24822 22480 24827 22536
rect 1761 22478 24827 22480
rect 1761 22475 1827 22478
rect 24761 22475 24827 22478
rect 4488 22336 4804 22337
rect 4488 22272 4494 22336
rect 4558 22272 4574 22336
rect 4638 22272 4654 22336
rect 4718 22272 4734 22336
rect 4798 22272 4804 22336
rect 4488 22271 4804 22272
rect 11572 22336 11888 22337
rect 11572 22272 11578 22336
rect 11642 22272 11658 22336
rect 11722 22272 11738 22336
rect 11802 22272 11818 22336
rect 11882 22272 11888 22336
rect 11572 22271 11888 22272
rect 18656 22336 18972 22337
rect 18656 22272 18662 22336
rect 18726 22272 18742 22336
rect 18806 22272 18822 22336
rect 18886 22272 18902 22336
rect 18966 22272 18972 22336
rect 18656 22271 18972 22272
rect 25740 22336 26056 22337
rect 25740 22272 25746 22336
rect 25810 22272 25826 22336
rect 25890 22272 25906 22336
rect 25970 22272 25986 22336
rect 26050 22272 26056 22336
rect 25740 22271 26056 22272
rect 21173 22130 21239 22133
rect 21173 22128 21282 22130
rect 21173 22072 21178 22128
rect 21234 22072 21282 22128
rect 21173 22067 21282 22072
rect 21222 21861 21282 22067
rect 17493 21858 17559 21861
rect 18965 21858 19031 21861
rect 17493 21856 19031 21858
rect 17493 21800 17498 21856
rect 17554 21800 18970 21856
rect 19026 21800 19031 21856
rect 17493 21798 19031 21800
rect 17493 21795 17559 21798
rect 18965 21795 19031 21798
rect 21173 21856 21282 21861
rect 21173 21800 21178 21856
rect 21234 21800 21282 21856
rect 21173 21798 21282 21800
rect 21173 21795 21239 21798
rect 8030 21792 8346 21793
rect 8030 21728 8036 21792
rect 8100 21728 8116 21792
rect 8180 21728 8196 21792
rect 8260 21728 8276 21792
rect 8340 21728 8346 21792
rect 8030 21727 8346 21728
rect 15114 21792 15430 21793
rect 15114 21728 15120 21792
rect 15184 21728 15200 21792
rect 15264 21728 15280 21792
rect 15344 21728 15360 21792
rect 15424 21728 15430 21792
rect 15114 21727 15430 21728
rect 22198 21792 22514 21793
rect 22198 21728 22204 21792
rect 22268 21728 22284 21792
rect 22348 21728 22364 21792
rect 22428 21728 22444 21792
rect 22508 21728 22514 21792
rect 22198 21727 22514 21728
rect 29282 21792 29598 21793
rect 29282 21728 29288 21792
rect 29352 21728 29368 21792
rect 29432 21728 29448 21792
rect 29512 21728 29528 21792
rect 29592 21728 29598 21792
rect 29282 21727 29598 21728
rect 4488 21248 4804 21249
rect 4488 21184 4494 21248
rect 4558 21184 4574 21248
rect 4638 21184 4654 21248
rect 4718 21184 4734 21248
rect 4798 21184 4804 21248
rect 4488 21183 4804 21184
rect 11572 21248 11888 21249
rect 11572 21184 11578 21248
rect 11642 21184 11658 21248
rect 11722 21184 11738 21248
rect 11802 21184 11818 21248
rect 11882 21184 11888 21248
rect 11572 21183 11888 21184
rect 18656 21248 18972 21249
rect 18656 21184 18662 21248
rect 18726 21184 18742 21248
rect 18806 21184 18822 21248
rect 18886 21184 18902 21248
rect 18966 21184 18972 21248
rect 18656 21183 18972 21184
rect 25740 21248 26056 21249
rect 25740 21184 25746 21248
rect 25810 21184 25826 21248
rect 25890 21184 25906 21248
rect 25970 21184 25986 21248
rect 26050 21184 26056 21248
rect 25740 21183 26056 21184
rect 28717 21178 28783 21181
rect 29821 21178 30621 21208
rect 28717 21176 30621 21178
rect 28717 21120 28722 21176
rect 28778 21120 30621 21176
rect 28717 21118 30621 21120
rect 28717 21115 28783 21118
rect 29821 21088 30621 21118
rect 8030 20704 8346 20705
rect 8030 20640 8036 20704
rect 8100 20640 8116 20704
rect 8180 20640 8196 20704
rect 8260 20640 8276 20704
rect 8340 20640 8346 20704
rect 8030 20639 8346 20640
rect 15114 20704 15430 20705
rect 15114 20640 15120 20704
rect 15184 20640 15200 20704
rect 15264 20640 15280 20704
rect 15344 20640 15360 20704
rect 15424 20640 15430 20704
rect 15114 20639 15430 20640
rect 22198 20704 22514 20705
rect 22198 20640 22204 20704
rect 22268 20640 22284 20704
rect 22348 20640 22364 20704
rect 22428 20640 22444 20704
rect 22508 20640 22514 20704
rect 22198 20639 22514 20640
rect 29282 20704 29598 20705
rect 29282 20640 29288 20704
rect 29352 20640 29368 20704
rect 29432 20640 29448 20704
rect 29512 20640 29528 20704
rect 29592 20640 29598 20704
rect 29282 20639 29598 20640
rect 4488 20160 4804 20161
rect 4488 20096 4494 20160
rect 4558 20096 4574 20160
rect 4638 20096 4654 20160
rect 4718 20096 4734 20160
rect 4798 20096 4804 20160
rect 4488 20095 4804 20096
rect 11572 20160 11888 20161
rect 11572 20096 11578 20160
rect 11642 20096 11658 20160
rect 11722 20096 11738 20160
rect 11802 20096 11818 20160
rect 11882 20096 11888 20160
rect 11572 20095 11888 20096
rect 18656 20160 18972 20161
rect 18656 20096 18662 20160
rect 18726 20096 18742 20160
rect 18806 20096 18822 20160
rect 18886 20096 18902 20160
rect 18966 20096 18972 20160
rect 18656 20095 18972 20096
rect 25740 20160 26056 20161
rect 25740 20096 25746 20160
rect 25810 20096 25826 20160
rect 25890 20096 25906 20160
rect 25970 20096 25986 20160
rect 26050 20096 26056 20160
rect 25740 20095 26056 20096
rect 0 19818 800 19848
rect 1485 19818 1551 19821
rect 0 19816 1551 19818
rect 0 19760 1490 19816
rect 1546 19760 1551 19816
rect 0 19758 1551 19760
rect 0 19728 800 19758
rect 1485 19755 1551 19758
rect 11513 19818 11579 19821
rect 27981 19818 28047 19821
rect 11513 19816 28047 19818
rect 11513 19760 11518 19816
rect 11574 19760 27986 19816
rect 28042 19760 28047 19816
rect 11513 19758 28047 19760
rect 11513 19755 11579 19758
rect 27981 19755 28047 19758
rect 8030 19616 8346 19617
rect 8030 19552 8036 19616
rect 8100 19552 8116 19616
rect 8180 19552 8196 19616
rect 8260 19552 8276 19616
rect 8340 19552 8346 19616
rect 8030 19551 8346 19552
rect 15114 19616 15430 19617
rect 15114 19552 15120 19616
rect 15184 19552 15200 19616
rect 15264 19552 15280 19616
rect 15344 19552 15360 19616
rect 15424 19552 15430 19616
rect 15114 19551 15430 19552
rect 22198 19616 22514 19617
rect 22198 19552 22204 19616
rect 22268 19552 22284 19616
rect 22348 19552 22364 19616
rect 22428 19552 22444 19616
rect 22508 19552 22514 19616
rect 22198 19551 22514 19552
rect 29282 19616 29598 19617
rect 29282 19552 29288 19616
rect 29352 19552 29368 19616
rect 29432 19552 29448 19616
rect 29512 19552 29528 19616
rect 29592 19552 29598 19616
rect 29282 19551 29598 19552
rect 13997 19410 14063 19413
rect 18045 19410 18111 19413
rect 13997 19408 18111 19410
rect 13997 19352 14002 19408
rect 14058 19352 18050 19408
rect 18106 19352 18111 19408
rect 13997 19350 18111 19352
rect 13997 19347 14063 19350
rect 18045 19347 18111 19350
rect 28717 19138 28783 19141
rect 29821 19138 30621 19168
rect 28717 19136 30621 19138
rect 28717 19080 28722 19136
rect 28778 19080 30621 19136
rect 28717 19078 30621 19080
rect 28717 19075 28783 19078
rect 4488 19072 4804 19073
rect 4488 19008 4494 19072
rect 4558 19008 4574 19072
rect 4638 19008 4654 19072
rect 4718 19008 4734 19072
rect 4798 19008 4804 19072
rect 4488 19007 4804 19008
rect 11572 19072 11888 19073
rect 11572 19008 11578 19072
rect 11642 19008 11658 19072
rect 11722 19008 11738 19072
rect 11802 19008 11818 19072
rect 11882 19008 11888 19072
rect 11572 19007 11888 19008
rect 18656 19072 18972 19073
rect 18656 19008 18662 19072
rect 18726 19008 18742 19072
rect 18806 19008 18822 19072
rect 18886 19008 18902 19072
rect 18966 19008 18972 19072
rect 18656 19007 18972 19008
rect 25740 19072 26056 19073
rect 25740 19008 25746 19072
rect 25810 19008 25826 19072
rect 25890 19008 25906 19072
rect 25970 19008 25986 19072
rect 26050 19008 26056 19072
rect 29821 19048 30621 19078
rect 25740 19007 26056 19008
rect 8030 18528 8346 18529
rect 8030 18464 8036 18528
rect 8100 18464 8116 18528
rect 8180 18464 8196 18528
rect 8260 18464 8276 18528
rect 8340 18464 8346 18528
rect 8030 18463 8346 18464
rect 15114 18528 15430 18529
rect 15114 18464 15120 18528
rect 15184 18464 15200 18528
rect 15264 18464 15280 18528
rect 15344 18464 15360 18528
rect 15424 18464 15430 18528
rect 15114 18463 15430 18464
rect 22198 18528 22514 18529
rect 22198 18464 22204 18528
rect 22268 18464 22284 18528
rect 22348 18464 22364 18528
rect 22428 18464 22444 18528
rect 22508 18464 22514 18528
rect 22198 18463 22514 18464
rect 29282 18528 29598 18529
rect 29282 18464 29288 18528
rect 29352 18464 29368 18528
rect 29432 18464 29448 18528
rect 29512 18464 29528 18528
rect 29592 18464 29598 18528
rect 29282 18463 29598 18464
rect 20713 18050 20779 18053
rect 20670 18048 20779 18050
rect 20670 17992 20718 18048
rect 20774 17992 20779 18048
rect 20670 17987 20779 17992
rect 4488 17984 4804 17985
rect 4488 17920 4494 17984
rect 4558 17920 4574 17984
rect 4638 17920 4654 17984
rect 4718 17920 4734 17984
rect 4798 17920 4804 17984
rect 4488 17919 4804 17920
rect 11572 17984 11888 17985
rect 11572 17920 11578 17984
rect 11642 17920 11658 17984
rect 11722 17920 11738 17984
rect 11802 17920 11818 17984
rect 11882 17920 11888 17984
rect 11572 17919 11888 17920
rect 18656 17984 18972 17985
rect 18656 17920 18662 17984
rect 18726 17920 18742 17984
rect 18806 17920 18822 17984
rect 18886 17920 18902 17984
rect 18966 17920 18972 17984
rect 18656 17919 18972 17920
rect 0 17778 800 17808
rect 1577 17778 1643 17781
rect 0 17776 1643 17778
rect 0 17720 1582 17776
rect 1638 17720 1643 17776
rect 0 17718 1643 17720
rect 0 17688 800 17718
rect 1577 17715 1643 17718
rect 17125 17778 17191 17781
rect 18505 17778 18571 17781
rect 20670 17778 20730 17987
rect 25740 17984 26056 17985
rect 25740 17920 25746 17984
rect 25810 17920 25826 17984
rect 25890 17920 25906 17984
rect 25970 17920 25986 17984
rect 26050 17920 26056 17984
rect 25740 17919 26056 17920
rect 17125 17776 20730 17778
rect 17125 17720 17130 17776
rect 17186 17720 18510 17776
rect 18566 17720 20730 17776
rect 17125 17718 20730 17720
rect 17125 17715 17191 17718
rect 18505 17715 18571 17718
rect 8030 17440 8346 17441
rect 8030 17376 8036 17440
rect 8100 17376 8116 17440
rect 8180 17376 8196 17440
rect 8260 17376 8276 17440
rect 8340 17376 8346 17440
rect 8030 17375 8346 17376
rect 15114 17440 15430 17441
rect 15114 17376 15120 17440
rect 15184 17376 15200 17440
rect 15264 17376 15280 17440
rect 15344 17376 15360 17440
rect 15424 17376 15430 17440
rect 15114 17375 15430 17376
rect 22198 17440 22514 17441
rect 22198 17376 22204 17440
rect 22268 17376 22284 17440
rect 22348 17376 22364 17440
rect 22428 17376 22444 17440
rect 22508 17376 22514 17440
rect 22198 17375 22514 17376
rect 29282 17440 29598 17441
rect 29282 17376 29288 17440
rect 29352 17376 29368 17440
rect 29432 17376 29448 17440
rect 29512 17376 29528 17440
rect 29592 17376 29598 17440
rect 29282 17375 29598 17376
rect 4488 16896 4804 16897
rect 4488 16832 4494 16896
rect 4558 16832 4574 16896
rect 4638 16832 4654 16896
rect 4718 16832 4734 16896
rect 4798 16832 4804 16896
rect 4488 16831 4804 16832
rect 11572 16896 11888 16897
rect 11572 16832 11578 16896
rect 11642 16832 11658 16896
rect 11722 16832 11738 16896
rect 11802 16832 11818 16896
rect 11882 16832 11888 16896
rect 11572 16831 11888 16832
rect 18656 16896 18972 16897
rect 18656 16832 18662 16896
rect 18726 16832 18742 16896
rect 18806 16832 18822 16896
rect 18886 16832 18902 16896
rect 18966 16832 18972 16896
rect 18656 16831 18972 16832
rect 25740 16896 26056 16897
rect 25740 16832 25746 16896
rect 25810 16832 25826 16896
rect 25890 16832 25906 16896
rect 25970 16832 25986 16896
rect 26050 16832 26056 16896
rect 25740 16831 26056 16832
rect 13353 16690 13419 16693
rect 20621 16692 20687 16693
rect 20621 16690 20668 16692
rect 13353 16688 20668 16690
rect 13353 16632 13358 16688
rect 13414 16632 20626 16688
rect 13353 16630 20668 16632
rect 13353 16627 13419 16630
rect 20621 16628 20668 16630
rect 20732 16628 20738 16692
rect 20621 16627 20687 16628
rect 11881 16554 11947 16557
rect 24025 16554 24091 16557
rect 11881 16552 24091 16554
rect 11881 16496 11886 16552
rect 11942 16496 24030 16552
rect 24086 16496 24091 16552
rect 11881 16494 24091 16496
rect 11881 16491 11947 16494
rect 24025 16491 24091 16494
rect 28717 16554 28783 16557
rect 28717 16552 29746 16554
rect 28717 16496 28722 16552
rect 28778 16496 29746 16552
rect 28717 16494 29746 16496
rect 28717 16491 28783 16494
rect 29686 16418 29746 16494
rect 29821 16418 30621 16448
rect 29686 16358 30621 16418
rect 8030 16352 8346 16353
rect 8030 16288 8036 16352
rect 8100 16288 8116 16352
rect 8180 16288 8196 16352
rect 8260 16288 8276 16352
rect 8340 16288 8346 16352
rect 8030 16287 8346 16288
rect 15114 16352 15430 16353
rect 15114 16288 15120 16352
rect 15184 16288 15200 16352
rect 15264 16288 15280 16352
rect 15344 16288 15360 16352
rect 15424 16288 15430 16352
rect 15114 16287 15430 16288
rect 22198 16352 22514 16353
rect 22198 16288 22204 16352
rect 22268 16288 22284 16352
rect 22348 16288 22364 16352
rect 22428 16288 22444 16352
rect 22508 16288 22514 16352
rect 22198 16287 22514 16288
rect 29282 16352 29598 16353
rect 29282 16288 29288 16352
rect 29352 16288 29368 16352
rect 29432 16288 29448 16352
rect 29512 16288 29528 16352
rect 29592 16288 29598 16352
rect 29821 16328 30621 16358
rect 29282 16287 29598 16288
rect 7649 16010 7715 16013
rect 7833 16010 7899 16013
rect 20253 16010 20319 16013
rect 7649 16008 20319 16010
rect 7649 15952 7654 16008
rect 7710 15952 7838 16008
rect 7894 15952 20258 16008
rect 20314 15952 20319 16008
rect 7649 15950 20319 15952
rect 7649 15947 7715 15950
rect 7833 15947 7899 15950
rect 20253 15947 20319 15950
rect 4488 15808 4804 15809
rect 0 15738 800 15768
rect 4488 15744 4494 15808
rect 4558 15744 4574 15808
rect 4638 15744 4654 15808
rect 4718 15744 4734 15808
rect 4798 15744 4804 15808
rect 4488 15743 4804 15744
rect 11572 15808 11888 15809
rect 11572 15744 11578 15808
rect 11642 15744 11658 15808
rect 11722 15744 11738 15808
rect 11802 15744 11818 15808
rect 11882 15744 11888 15808
rect 11572 15743 11888 15744
rect 18656 15808 18972 15809
rect 18656 15744 18662 15808
rect 18726 15744 18742 15808
rect 18806 15744 18822 15808
rect 18886 15744 18902 15808
rect 18966 15744 18972 15808
rect 18656 15743 18972 15744
rect 25740 15808 26056 15809
rect 25740 15744 25746 15808
rect 25810 15744 25826 15808
rect 25890 15744 25906 15808
rect 25970 15744 25986 15808
rect 26050 15744 26056 15808
rect 25740 15743 26056 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 10869 15466 10935 15469
rect 16389 15466 16455 15469
rect 10869 15464 16455 15466
rect 10869 15408 10874 15464
rect 10930 15408 16394 15464
rect 16450 15408 16455 15464
rect 10869 15406 16455 15408
rect 10869 15403 10935 15406
rect 16389 15403 16455 15406
rect 8030 15264 8346 15265
rect 8030 15200 8036 15264
rect 8100 15200 8116 15264
rect 8180 15200 8196 15264
rect 8260 15200 8276 15264
rect 8340 15200 8346 15264
rect 8030 15199 8346 15200
rect 15114 15264 15430 15265
rect 15114 15200 15120 15264
rect 15184 15200 15200 15264
rect 15264 15200 15280 15264
rect 15344 15200 15360 15264
rect 15424 15200 15430 15264
rect 15114 15199 15430 15200
rect 22198 15264 22514 15265
rect 22198 15200 22204 15264
rect 22268 15200 22284 15264
rect 22348 15200 22364 15264
rect 22428 15200 22444 15264
rect 22508 15200 22514 15264
rect 22198 15199 22514 15200
rect 29282 15264 29598 15265
rect 29282 15200 29288 15264
rect 29352 15200 29368 15264
rect 29432 15200 29448 15264
rect 29512 15200 29528 15264
rect 29592 15200 29598 15264
rect 29282 15199 29598 15200
rect 9397 14922 9463 14925
rect 18045 14922 18111 14925
rect 9397 14920 18111 14922
rect 9397 14864 9402 14920
rect 9458 14864 18050 14920
rect 18106 14864 18111 14920
rect 9397 14862 18111 14864
rect 9397 14859 9463 14862
rect 18045 14859 18111 14862
rect 4488 14720 4804 14721
rect 4488 14656 4494 14720
rect 4558 14656 4574 14720
rect 4638 14656 4654 14720
rect 4718 14656 4734 14720
rect 4798 14656 4804 14720
rect 4488 14655 4804 14656
rect 11572 14720 11888 14721
rect 11572 14656 11578 14720
rect 11642 14656 11658 14720
rect 11722 14656 11738 14720
rect 11802 14656 11818 14720
rect 11882 14656 11888 14720
rect 11572 14655 11888 14656
rect 18656 14720 18972 14721
rect 18656 14656 18662 14720
rect 18726 14656 18742 14720
rect 18806 14656 18822 14720
rect 18886 14656 18902 14720
rect 18966 14656 18972 14720
rect 18656 14655 18972 14656
rect 25740 14720 26056 14721
rect 25740 14656 25746 14720
rect 25810 14656 25826 14720
rect 25890 14656 25906 14720
rect 25970 14656 25986 14720
rect 26050 14656 26056 14720
rect 25740 14655 26056 14656
rect 20621 14650 20687 14653
rect 21633 14650 21699 14653
rect 20621 14648 21699 14650
rect 20621 14592 20626 14648
rect 20682 14592 21638 14648
rect 21694 14592 21699 14648
rect 20621 14590 21699 14592
rect 20621 14587 20687 14590
rect 21633 14587 21699 14590
rect 11605 14514 11671 14517
rect 25037 14514 25103 14517
rect 11605 14512 25103 14514
rect 11605 14456 11610 14512
rect 11666 14456 25042 14512
rect 25098 14456 25103 14512
rect 11605 14454 25103 14456
rect 11605 14451 11671 14454
rect 25037 14451 25103 14454
rect 28625 14378 28691 14381
rect 29821 14378 30621 14408
rect 28625 14376 30621 14378
rect 28625 14320 28630 14376
rect 28686 14320 30621 14376
rect 28625 14318 30621 14320
rect 28625 14315 28691 14318
rect 29821 14288 30621 14318
rect 8030 14176 8346 14177
rect 8030 14112 8036 14176
rect 8100 14112 8116 14176
rect 8180 14112 8196 14176
rect 8260 14112 8276 14176
rect 8340 14112 8346 14176
rect 8030 14111 8346 14112
rect 15114 14176 15430 14177
rect 15114 14112 15120 14176
rect 15184 14112 15200 14176
rect 15264 14112 15280 14176
rect 15344 14112 15360 14176
rect 15424 14112 15430 14176
rect 15114 14111 15430 14112
rect 22198 14176 22514 14177
rect 22198 14112 22204 14176
rect 22268 14112 22284 14176
rect 22348 14112 22364 14176
rect 22428 14112 22444 14176
rect 22508 14112 22514 14176
rect 22198 14111 22514 14112
rect 29282 14176 29598 14177
rect 29282 14112 29288 14176
rect 29352 14112 29368 14176
rect 29432 14112 29448 14176
rect 29512 14112 29528 14176
rect 29592 14112 29598 14176
rect 29282 14111 29598 14112
rect 7557 13970 7623 13973
rect 28441 13970 28507 13973
rect 7557 13968 28507 13970
rect 7557 13912 7562 13968
rect 7618 13912 28446 13968
rect 28502 13912 28507 13968
rect 7557 13910 28507 13912
rect 7557 13907 7623 13910
rect 28441 13907 28507 13910
rect 4488 13632 4804 13633
rect 4488 13568 4494 13632
rect 4558 13568 4574 13632
rect 4638 13568 4654 13632
rect 4718 13568 4734 13632
rect 4798 13568 4804 13632
rect 4488 13567 4804 13568
rect 11572 13632 11888 13633
rect 11572 13568 11578 13632
rect 11642 13568 11658 13632
rect 11722 13568 11738 13632
rect 11802 13568 11818 13632
rect 11882 13568 11888 13632
rect 11572 13567 11888 13568
rect 18656 13632 18972 13633
rect 18656 13568 18662 13632
rect 18726 13568 18742 13632
rect 18806 13568 18822 13632
rect 18886 13568 18902 13632
rect 18966 13568 18972 13632
rect 18656 13567 18972 13568
rect 25740 13632 26056 13633
rect 25740 13568 25746 13632
rect 25810 13568 25826 13632
rect 25890 13568 25906 13632
rect 25970 13568 25986 13632
rect 26050 13568 26056 13632
rect 25740 13567 26056 13568
rect 8030 13088 8346 13089
rect 0 13018 800 13048
rect 8030 13024 8036 13088
rect 8100 13024 8116 13088
rect 8180 13024 8196 13088
rect 8260 13024 8276 13088
rect 8340 13024 8346 13088
rect 8030 13023 8346 13024
rect 15114 13088 15430 13089
rect 15114 13024 15120 13088
rect 15184 13024 15200 13088
rect 15264 13024 15280 13088
rect 15344 13024 15360 13088
rect 15424 13024 15430 13088
rect 15114 13023 15430 13024
rect 22198 13088 22514 13089
rect 22198 13024 22204 13088
rect 22268 13024 22284 13088
rect 22348 13024 22364 13088
rect 22428 13024 22444 13088
rect 22508 13024 22514 13088
rect 22198 13023 22514 13024
rect 29282 13088 29598 13089
rect 29282 13024 29288 13088
rect 29352 13024 29368 13088
rect 29432 13024 29448 13088
rect 29512 13024 29528 13088
rect 29592 13024 29598 13088
rect 29282 13023 29598 13024
rect 1485 13018 1551 13021
rect 0 13016 1551 13018
rect 0 12960 1490 13016
rect 1546 12960 1551 13016
rect 0 12958 1551 12960
rect 0 12928 800 12958
rect 1485 12955 1551 12958
rect 20897 13018 20963 13021
rect 21030 13018 21036 13020
rect 20897 13016 21036 13018
rect 20897 12960 20902 13016
rect 20958 12960 21036 13016
rect 20897 12958 21036 12960
rect 20897 12955 20963 12958
rect 21030 12956 21036 12958
rect 21100 12956 21106 13020
rect 4488 12544 4804 12545
rect 4488 12480 4494 12544
rect 4558 12480 4574 12544
rect 4638 12480 4654 12544
rect 4718 12480 4734 12544
rect 4798 12480 4804 12544
rect 4488 12479 4804 12480
rect 11572 12544 11888 12545
rect 11572 12480 11578 12544
rect 11642 12480 11658 12544
rect 11722 12480 11738 12544
rect 11802 12480 11818 12544
rect 11882 12480 11888 12544
rect 11572 12479 11888 12480
rect 18656 12544 18972 12545
rect 18656 12480 18662 12544
rect 18726 12480 18742 12544
rect 18806 12480 18822 12544
rect 18886 12480 18902 12544
rect 18966 12480 18972 12544
rect 18656 12479 18972 12480
rect 25740 12544 26056 12545
rect 25740 12480 25746 12544
rect 25810 12480 25826 12544
rect 25890 12480 25906 12544
rect 25970 12480 25986 12544
rect 26050 12480 26056 12544
rect 25740 12479 26056 12480
rect 27981 12474 28047 12477
rect 28349 12474 28415 12477
rect 27981 12472 28415 12474
rect 27981 12416 27986 12472
rect 28042 12416 28354 12472
rect 28410 12416 28415 12472
rect 27981 12414 28415 12416
rect 27981 12411 28047 12414
rect 28349 12411 28415 12414
rect 11329 12338 11395 12341
rect 18413 12338 18479 12341
rect 11329 12336 18479 12338
rect 11329 12280 11334 12336
rect 11390 12280 18418 12336
rect 18474 12280 18479 12336
rect 11329 12278 18479 12280
rect 11329 12275 11395 12278
rect 18413 12275 18479 12278
rect 28625 12338 28691 12341
rect 29821 12338 30621 12368
rect 28625 12336 30621 12338
rect 28625 12280 28630 12336
rect 28686 12280 30621 12336
rect 28625 12278 30621 12280
rect 28625 12275 28691 12278
rect 29821 12248 30621 12278
rect 15377 12202 15443 12205
rect 20662 12202 20668 12204
rect 15377 12200 20668 12202
rect 15377 12144 15382 12200
rect 15438 12144 20668 12200
rect 15377 12142 20668 12144
rect 15377 12139 15443 12142
rect 20662 12140 20668 12142
rect 20732 12140 20738 12204
rect 8030 12000 8346 12001
rect 8030 11936 8036 12000
rect 8100 11936 8116 12000
rect 8180 11936 8196 12000
rect 8260 11936 8276 12000
rect 8340 11936 8346 12000
rect 8030 11935 8346 11936
rect 15114 12000 15430 12001
rect 15114 11936 15120 12000
rect 15184 11936 15200 12000
rect 15264 11936 15280 12000
rect 15344 11936 15360 12000
rect 15424 11936 15430 12000
rect 15114 11935 15430 11936
rect 22198 12000 22514 12001
rect 22198 11936 22204 12000
rect 22268 11936 22284 12000
rect 22348 11936 22364 12000
rect 22428 11936 22444 12000
rect 22508 11936 22514 12000
rect 22198 11935 22514 11936
rect 29282 12000 29598 12001
rect 29282 11936 29288 12000
rect 29352 11936 29368 12000
rect 29432 11936 29448 12000
rect 29512 11936 29528 12000
rect 29592 11936 29598 12000
rect 29282 11935 29598 11936
rect 4488 11456 4804 11457
rect 4488 11392 4494 11456
rect 4558 11392 4574 11456
rect 4638 11392 4654 11456
rect 4718 11392 4734 11456
rect 4798 11392 4804 11456
rect 4488 11391 4804 11392
rect 11572 11456 11888 11457
rect 11572 11392 11578 11456
rect 11642 11392 11658 11456
rect 11722 11392 11738 11456
rect 11802 11392 11818 11456
rect 11882 11392 11888 11456
rect 11572 11391 11888 11392
rect 18656 11456 18972 11457
rect 18656 11392 18662 11456
rect 18726 11392 18742 11456
rect 18806 11392 18822 11456
rect 18886 11392 18902 11456
rect 18966 11392 18972 11456
rect 18656 11391 18972 11392
rect 25740 11456 26056 11457
rect 25740 11392 25746 11456
rect 25810 11392 25826 11456
rect 25890 11392 25906 11456
rect 25970 11392 25986 11456
rect 26050 11392 26056 11456
rect 25740 11391 26056 11392
rect 12893 11250 12959 11253
rect 23933 11250 23999 11253
rect 12893 11248 23999 11250
rect 12893 11192 12898 11248
rect 12954 11192 23938 11248
rect 23994 11192 23999 11248
rect 12893 11190 23999 11192
rect 12893 11187 12959 11190
rect 23933 11187 23999 11190
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 8030 10912 8346 10913
rect 8030 10848 8036 10912
rect 8100 10848 8116 10912
rect 8180 10848 8196 10912
rect 8260 10848 8276 10912
rect 8340 10848 8346 10912
rect 8030 10847 8346 10848
rect 15114 10912 15430 10913
rect 15114 10848 15120 10912
rect 15184 10848 15200 10912
rect 15264 10848 15280 10912
rect 15344 10848 15360 10912
rect 15424 10848 15430 10912
rect 15114 10847 15430 10848
rect 22198 10912 22514 10913
rect 22198 10848 22204 10912
rect 22268 10848 22284 10912
rect 22348 10848 22364 10912
rect 22428 10848 22444 10912
rect 22508 10848 22514 10912
rect 22198 10847 22514 10848
rect 29282 10912 29598 10913
rect 29282 10848 29288 10912
rect 29352 10848 29368 10912
rect 29432 10848 29448 10912
rect 29512 10848 29528 10912
rect 29592 10848 29598 10912
rect 29282 10847 29598 10848
rect 14549 10706 14615 10709
rect 18321 10706 18387 10709
rect 24393 10706 24459 10709
rect 14549 10704 24459 10706
rect 14549 10648 14554 10704
rect 14610 10648 18326 10704
rect 18382 10648 24398 10704
rect 24454 10648 24459 10704
rect 14549 10646 24459 10648
rect 14549 10643 14615 10646
rect 18321 10643 18387 10646
rect 24393 10643 24459 10646
rect 14365 10570 14431 10573
rect 24209 10570 24275 10573
rect 14365 10568 24275 10570
rect 14365 10512 14370 10568
rect 14426 10512 24214 10568
rect 24270 10512 24275 10568
rect 14365 10510 24275 10512
rect 14365 10507 14431 10510
rect 24209 10507 24275 10510
rect 4488 10368 4804 10369
rect 4488 10304 4494 10368
rect 4558 10304 4574 10368
rect 4638 10304 4654 10368
rect 4718 10304 4734 10368
rect 4798 10304 4804 10368
rect 4488 10303 4804 10304
rect 11572 10368 11888 10369
rect 11572 10304 11578 10368
rect 11642 10304 11658 10368
rect 11722 10304 11738 10368
rect 11802 10304 11818 10368
rect 11882 10304 11888 10368
rect 11572 10303 11888 10304
rect 18656 10368 18972 10369
rect 18656 10304 18662 10368
rect 18726 10304 18742 10368
rect 18806 10304 18822 10368
rect 18886 10304 18902 10368
rect 18966 10304 18972 10368
rect 18656 10303 18972 10304
rect 25740 10368 26056 10369
rect 25740 10304 25746 10368
rect 25810 10304 25826 10368
rect 25890 10304 25906 10368
rect 25970 10304 25986 10368
rect 26050 10304 26056 10368
rect 25740 10303 26056 10304
rect 21633 10162 21699 10165
rect 25497 10162 25563 10165
rect 21633 10160 25563 10162
rect 21633 10104 21638 10160
rect 21694 10104 25502 10160
rect 25558 10104 25563 10160
rect 21633 10102 25563 10104
rect 21633 10099 21699 10102
rect 25497 10099 25563 10102
rect 19333 10026 19399 10029
rect 23657 10026 23723 10029
rect 19333 10024 23723 10026
rect 19333 9968 19338 10024
rect 19394 9968 23662 10024
rect 23718 9968 23723 10024
rect 19333 9966 23723 9968
rect 19333 9963 19399 9966
rect 23657 9963 23723 9966
rect 8030 9824 8346 9825
rect 8030 9760 8036 9824
rect 8100 9760 8116 9824
rect 8180 9760 8196 9824
rect 8260 9760 8276 9824
rect 8340 9760 8346 9824
rect 8030 9759 8346 9760
rect 15114 9824 15430 9825
rect 15114 9760 15120 9824
rect 15184 9760 15200 9824
rect 15264 9760 15280 9824
rect 15344 9760 15360 9824
rect 15424 9760 15430 9824
rect 15114 9759 15430 9760
rect 22198 9824 22514 9825
rect 22198 9760 22204 9824
rect 22268 9760 22284 9824
rect 22348 9760 22364 9824
rect 22428 9760 22444 9824
rect 22508 9760 22514 9824
rect 22198 9759 22514 9760
rect 29282 9824 29598 9825
rect 29282 9760 29288 9824
rect 29352 9760 29368 9824
rect 29432 9760 29448 9824
rect 29512 9760 29528 9824
rect 29592 9760 29598 9824
rect 29282 9759 29598 9760
rect 7281 9618 7347 9621
rect 11237 9618 11303 9621
rect 7281 9616 11303 9618
rect 7281 9560 7286 9616
rect 7342 9560 11242 9616
rect 11298 9560 11303 9616
rect 7281 9558 11303 9560
rect 7281 9555 7347 9558
rect 11237 9555 11303 9558
rect 15285 9618 15351 9621
rect 26509 9618 26575 9621
rect 15285 9616 26575 9618
rect 15285 9560 15290 9616
rect 15346 9560 26514 9616
rect 26570 9560 26575 9616
rect 15285 9558 26575 9560
rect 15285 9555 15351 9558
rect 26509 9555 26575 9558
rect 28717 9618 28783 9621
rect 29821 9618 30621 9648
rect 28717 9616 30621 9618
rect 28717 9560 28722 9616
rect 28778 9560 30621 9616
rect 28717 9558 30621 9560
rect 28717 9555 28783 9558
rect 29821 9528 30621 9558
rect 20989 9482 21055 9485
rect 23473 9482 23539 9485
rect 20989 9480 23539 9482
rect 20989 9424 20994 9480
rect 21050 9424 23478 9480
rect 23534 9424 23539 9480
rect 20989 9422 23539 9424
rect 20989 9419 21055 9422
rect 23473 9419 23539 9422
rect 4488 9280 4804 9281
rect 4488 9216 4494 9280
rect 4558 9216 4574 9280
rect 4638 9216 4654 9280
rect 4718 9216 4734 9280
rect 4798 9216 4804 9280
rect 4488 9215 4804 9216
rect 11572 9280 11888 9281
rect 11572 9216 11578 9280
rect 11642 9216 11658 9280
rect 11722 9216 11738 9280
rect 11802 9216 11818 9280
rect 11882 9216 11888 9280
rect 11572 9215 11888 9216
rect 18656 9280 18972 9281
rect 18656 9216 18662 9280
rect 18726 9216 18742 9280
rect 18806 9216 18822 9280
rect 18886 9216 18902 9280
rect 18966 9216 18972 9280
rect 18656 9215 18972 9216
rect 25740 9280 26056 9281
rect 25740 9216 25746 9280
rect 25810 9216 25826 9280
rect 25890 9216 25906 9280
rect 25970 9216 25986 9280
rect 26050 9216 26056 9280
rect 25740 9215 26056 9216
rect 0 8938 800 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 800 8878
rect 1577 8875 1643 8878
rect 7925 8938 7991 8941
rect 27889 8938 27955 8941
rect 7925 8936 27955 8938
rect 7925 8880 7930 8936
rect 7986 8880 27894 8936
rect 27950 8880 27955 8936
rect 7925 8878 27955 8880
rect 7925 8875 7991 8878
rect 27889 8875 27955 8878
rect 8030 8736 8346 8737
rect 8030 8672 8036 8736
rect 8100 8672 8116 8736
rect 8180 8672 8196 8736
rect 8260 8672 8276 8736
rect 8340 8672 8346 8736
rect 8030 8671 8346 8672
rect 15114 8736 15430 8737
rect 15114 8672 15120 8736
rect 15184 8672 15200 8736
rect 15264 8672 15280 8736
rect 15344 8672 15360 8736
rect 15424 8672 15430 8736
rect 15114 8671 15430 8672
rect 22198 8736 22514 8737
rect 22198 8672 22204 8736
rect 22268 8672 22284 8736
rect 22348 8672 22364 8736
rect 22428 8672 22444 8736
rect 22508 8672 22514 8736
rect 22198 8671 22514 8672
rect 29282 8736 29598 8737
rect 29282 8672 29288 8736
rect 29352 8672 29368 8736
rect 29432 8672 29448 8736
rect 29512 8672 29528 8736
rect 29592 8672 29598 8736
rect 29282 8671 29598 8672
rect 2681 8530 2747 8533
rect 20069 8530 20135 8533
rect 2681 8528 20135 8530
rect 2681 8472 2686 8528
rect 2742 8472 20074 8528
rect 20130 8472 20135 8528
rect 2681 8470 20135 8472
rect 2681 8467 2747 8470
rect 20069 8467 20135 8470
rect 4488 8192 4804 8193
rect 4488 8128 4494 8192
rect 4558 8128 4574 8192
rect 4638 8128 4654 8192
rect 4718 8128 4734 8192
rect 4798 8128 4804 8192
rect 4488 8127 4804 8128
rect 11572 8192 11888 8193
rect 11572 8128 11578 8192
rect 11642 8128 11658 8192
rect 11722 8128 11738 8192
rect 11802 8128 11818 8192
rect 11882 8128 11888 8192
rect 11572 8127 11888 8128
rect 18656 8192 18972 8193
rect 18656 8128 18662 8192
rect 18726 8128 18742 8192
rect 18806 8128 18822 8192
rect 18886 8128 18902 8192
rect 18966 8128 18972 8192
rect 18656 8127 18972 8128
rect 25740 8192 26056 8193
rect 25740 8128 25746 8192
rect 25810 8128 25826 8192
rect 25890 8128 25906 8192
rect 25970 8128 25986 8192
rect 26050 8128 26056 8192
rect 25740 8127 26056 8128
rect 21909 7850 21975 7853
rect 22686 7850 22692 7852
rect 21909 7848 22692 7850
rect 21909 7792 21914 7848
rect 21970 7792 22692 7848
rect 21909 7790 22692 7792
rect 21909 7787 21975 7790
rect 22686 7788 22692 7790
rect 22756 7788 22762 7852
rect 8030 7648 8346 7649
rect 8030 7584 8036 7648
rect 8100 7584 8116 7648
rect 8180 7584 8196 7648
rect 8260 7584 8276 7648
rect 8340 7584 8346 7648
rect 8030 7583 8346 7584
rect 15114 7648 15430 7649
rect 15114 7584 15120 7648
rect 15184 7584 15200 7648
rect 15264 7584 15280 7648
rect 15344 7584 15360 7648
rect 15424 7584 15430 7648
rect 15114 7583 15430 7584
rect 22198 7648 22514 7649
rect 22198 7584 22204 7648
rect 22268 7584 22284 7648
rect 22348 7584 22364 7648
rect 22428 7584 22444 7648
rect 22508 7584 22514 7648
rect 22198 7583 22514 7584
rect 29282 7648 29598 7649
rect 29282 7584 29288 7648
rect 29352 7584 29368 7648
rect 29432 7584 29448 7648
rect 29512 7584 29528 7648
rect 29592 7584 29598 7648
rect 29282 7583 29598 7584
rect 29821 7578 30621 7608
rect 29686 7518 30621 7578
rect 28717 7442 28783 7445
rect 29686 7442 29746 7518
rect 29821 7488 30621 7518
rect 28717 7440 29746 7442
rect 28717 7384 28722 7440
rect 28778 7384 29746 7440
rect 28717 7382 29746 7384
rect 28717 7379 28783 7382
rect 3417 7306 3483 7309
rect 16665 7306 16731 7309
rect 3417 7304 16731 7306
rect 3417 7248 3422 7304
rect 3478 7248 16670 7304
rect 16726 7248 16731 7304
rect 3417 7246 16731 7248
rect 3417 7243 3483 7246
rect 16665 7243 16731 7246
rect 4488 7104 4804 7105
rect 4488 7040 4494 7104
rect 4558 7040 4574 7104
rect 4638 7040 4654 7104
rect 4718 7040 4734 7104
rect 4798 7040 4804 7104
rect 4488 7039 4804 7040
rect 11572 7104 11888 7105
rect 11572 7040 11578 7104
rect 11642 7040 11658 7104
rect 11722 7040 11738 7104
rect 11802 7040 11818 7104
rect 11882 7040 11888 7104
rect 11572 7039 11888 7040
rect 18656 7104 18972 7105
rect 18656 7040 18662 7104
rect 18726 7040 18742 7104
rect 18806 7040 18822 7104
rect 18886 7040 18902 7104
rect 18966 7040 18972 7104
rect 18656 7039 18972 7040
rect 25740 7104 26056 7105
rect 25740 7040 25746 7104
rect 25810 7040 25826 7104
rect 25890 7040 25906 7104
rect 25970 7040 25986 7104
rect 26050 7040 26056 7104
rect 25740 7039 26056 7040
rect 19517 6898 19583 6901
rect 19977 6898 20043 6901
rect 19517 6896 20043 6898
rect 19517 6840 19522 6896
rect 19578 6840 19982 6896
rect 20038 6840 20043 6896
rect 19517 6838 20043 6840
rect 19517 6835 19583 6838
rect 19977 6835 20043 6838
rect 8030 6560 8346 6561
rect 8030 6496 8036 6560
rect 8100 6496 8116 6560
rect 8180 6496 8196 6560
rect 8260 6496 8276 6560
rect 8340 6496 8346 6560
rect 8030 6495 8346 6496
rect 15114 6560 15430 6561
rect 15114 6496 15120 6560
rect 15184 6496 15200 6560
rect 15264 6496 15280 6560
rect 15344 6496 15360 6560
rect 15424 6496 15430 6560
rect 15114 6495 15430 6496
rect 22198 6560 22514 6561
rect 22198 6496 22204 6560
rect 22268 6496 22284 6560
rect 22348 6496 22364 6560
rect 22428 6496 22444 6560
rect 22508 6496 22514 6560
rect 22198 6495 22514 6496
rect 29282 6560 29598 6561
rect 29282 6496 29288 6560
rect 29352 6496 29368 6560
rect 29432 6496 29448 6560
rect 29512 6496 29528 6560
rect 29592 6496 29598 6560
rect 29282 6495 29598 6496
rect 0 6218 800 6248
rect 1393 6218 1459 6221
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 800 6158
rect 1393 6155 1459 6158
rect 1669 6218 1735 6221
rect 16573 6218 16639 6221
rect 1669 6216 16639 6218
rect 1669 6160 1674 6216
rect 1730 6160 16578 6216
rect 16634 6160 16639 6216
rect 1669 6158 16639 6160
rect 1669 6155 1735 6158
rect 16573 6155 16639 6158
rect 4488 6016 4804 6017
rect 4488 5952 4494 6016
rect 4558 5952 4574 6016
rect 4638 5952 4654 6016
rect 4718 5952 4734 6016
rect 4798 5952 4804 6016
rect 4488 5951 4804 5952
rect 11572 6016 11888 6017
rect 11572 5952 11578 6016
rect 11642 5952 11658 6016
rect 11722 5952 11738 6016
rect 11802 5952 11818 6016
rect 11882 5952 11888 6016
rect 11572 5951 11888 5952
rect 18656 6016 18972 6017
rect 18656 5952 18662 6016
rect 18726 5952 18742 6016
rect 18806 5952 18822 6016
rect 18886 5952 18902 6016
rect 18966 5952 18972 6016
rect 18656 5951 18972 5952
rect 25740 6016 26056 6017
rect 25740 5952 25746 6016
rect 25810 5952 25826 6016
rect 25890 5952 25906 6016
rect 25970 5952 25986 6016
rect 26050 5952 26056 6016
rect 25740 5951 26056 5952
rect 29821 5538 30621 5568
rect 29686 5478 30621 5538
rect 8030 5472 8346 5473
rect 8030 5408 8036 5472
rect 8100 5408 8116 5472
rect 8180 5408 8196 5472
rect 8260 5408 8276 5472
rect 8340 5408 8346 5472
rect 8030 5407 8346 5408
rect 15114 5472 15430 5473
rect 15114 5408 15120 5472
rect 15184 5408 15200 5472
rect 15264 5408 15280 5472
rect 15344 5408 15360 5472
rect 15424 5408 15430 5472
rect 15114 5407 15430 5408
rect 22198 5472 22514 5473
rect 22198 5408 22204 5472
rect 22268 5408 22284 5472
rect 22348 5408 22364 5472
rect 22428 5408 22444 5472
rect 22508 5408 22514 5472
rect 22198 5407 22514 5408
rect 29282 5472 29598 5473
rect 29282 5408 29288 5472
rect 29352 5408 29368 5472
rect 29432 5408 29448 5472
rect 29512 5408 29528 5472
rect 29592 5408 29598 5472
rect 29282 5407 29598 5408
rect 28717 5266 28783 5269
rect 29686 5266 29746 5478
rect 29821 5448 30621 5478
rect 28717 5264 29746 5266
rect 28717 5208 28722 5264
rect 28778 5208 29746 5264
rect 28717 5206 29746 5208
rect 28717 5203 28783 5206
rect 23473 5130 23539 5133
rect 27838 5130 27844 5132
rect 23473 5128 27844 5130
rect 23473 5072 23478 5128
rect 23534 5072 27844 5128
rect 23473 5070 27844 5072
rect 23473 5067 23539 5070
rect 27838 5068 27844 5070
rect 27908 5068 27914 5132
rect 4488 4928 4804 4929
rect 4488 4864 4494 4928
rect 4558 4864 4574 4928
rect 4638 4864 4654 4928
rect 4718 4864 4734 4928
rect 4798 4864 4804 4928
rect 4488 4863 4804 4864
rect 11572 4928 11888 4929
rect 11572 4864 11578 4928
rect 11642 4864 11658 4928
rect 11722 4864 11738 4928
rect 11802 4864 11818 4928
rect 11882 4864 11888 4928
rect 11572 4863 11888 4864
rect 18656 4928 18972 4929
rect 18656 4864 18662 4928
rect 18726 4864 18742 4928
rect 18806 4864 18822 4928
rect 18886 4864 18902 4928
rect 18966 4864 18972 4928
rect 18656 4863 18972 4864
rect 25740 4928 26056 4929
rect 25740 4864 25746 4928
rect 25810 4864 25826 4928
rect 25890 4864 25906 4928
rect 25970 4864 25986 4928
rect 26050 4864 26056 4928
rect 25740 4863 26056 4864
rect 8030 4384 8346 4385
rect 8030 4320 8036 4384
rect 8100 4320 8116 4384
rect 8180 4320 8196 4384
rect 8260 4320 8276 4384
rect 8340 4320 8346 4384
rect 8030 4319 8346 4320
rect 15114 4384 15430 4385
rect 15114 4320 15120 4384
rect 15184 4320 15200 4384
rect 15264 4320 15280 4384
rect 15344 4320 15360 4384
rect 15424 4320 15430 4384
rect 15114 4319 15430 4320
rect 22198 4384 22514 4385
rect 22198 4320 22204 4384
rect 22268 4320 22284 4384
rect 22348 4320 22364 4384
rect 22428 4320 22444 4384
rect 22508 4320 22514 4384
rect 22198 4319 22514 4320
rect 29282 4384 29598 4385
rect 29282 4320 29288 4384
rect 29352 4320 29368 4384
rect 29432 4320 29448 4384
rect 29512 4320 29528 4384
rect 29592 4320 29598 4384
rect 29282 4319 29598 4320
rect 0 4178 800 4208
rect 1577 4178 1643 4181
rect 23473 4178 23539 4181
rect 0 4176 1643 4178
rect 0 4120 1582 4176
rect 1638 4120 1643 4176
rect 0 4118 1643 4120
rect 0 4088 800 4118
rect 1577 4115 1643 4118
rect 22050 4176 23539 4178
rect 22050 4120 23478 4176
rect 23534 4120 23539 4176
rect 22050 4118 23539 4120
rect 2957 4042 3023 4045
rect 22050 4042 22110 4118
rect 23473 4115 23539 4118
rect 2957 4040 22110 4042
rect 2957 3984 2962 4040
rect 3018 3984 22110 4040
rect 2957 3982 22110 3984
rect 2957 3979 3023 3982
rect 4488 3840 4804 3841
rect 4488 3776 4494 3840
rect 4558 3776 4574 3840
rect 4638 3776 4654 3840
rect 4718 3776 4734 3840
rect 4798 3776 4804 3840
rect 4488 3775 4804 3776
rect 11572 3840 11888 3841
rect 11572 3776 11578 3840
rect 11642 3776 11658 3840
rect 11722 3776 11738 3840
rect 11802 3776 11818 3840
rect 11882 3776 11888 3840
rect 11572 3775 11888 3776
rect 18656 3840 18972 3841
rect 18656 3776 18662 3840
rect 18726 3776 18742 3840
rect 18806 3776 18822 3840
rect 18886 3776 18902 3840
rect 18966 3776 18972 3840
rect 18656 3775 18972 3776
rect 25740 3840 26056 3841
rect 25740 3776 25746 3840
rect 25810 3776 25826 3840
rect 25890 3776 25906 3840
rect 25970 3776 25986 3840
rect 26050 3776 26056 3840
rect 25740 3775 26056 3776
rect 16389 3498 16455 3501
rect 17677 3498 17743 3501
rect 16389 3496 17743 3498
rect 16389 3440 16394 3496
rect 16450 3440 17682 3496
rect 17738 3440 17743 3496
rect 16389 3438 17743 3440
rect 16389 3435 16455 3438
rect 17677 3435 17743 3438
rect 8030 3296 8346 3297
rect 8030 3232 8036 3296
rect 8100 3232 8116 3296
rect 8180 3232 8196 3296
rect 8260 3232 8276 3296
rect 8340 3232 8346 3296
rect 8030 3231 8346 3232
rect 15114 3296 15430 3297
rect 15114 3232 15120 3296
rect 15184 3232 15200 3296
rect 15264 3232 15280 3296
rect 15344 3232 15360 3296
rect 15424 3232 15430 3296
rect 15114 3231 15430 3232
rect 22198 3296 22514 3297
rect 22198 3232 22204 3296
rect 22268 3232 22284 3296
rect 22348 3232 22364 3296
rect 22428 3232 22444 3296
rect 22508 3232 22514 3296
rect 22198 3231 22514 3232
rect 29282 3296 29598 3297
rect 29282 3232 29288 3296
rect 29352 3232 29368 3296
rect 29432 3232 29448 3296
rect 29512 3232 29528 3296
rect 29592 3232 29598 3296
rect 29282 3231 29598 3232
rect 28625 2818 28691 2821
rect 29821 2818 30621 2848
rect 28625 2816 30621 2818
rect 28625 2760 28630 2816
rect 28686 2760 30621 2816
rect 28625 2758 30621 2760
rect 28625 2755 28691 2758
rect 4488 2752 4804 2753
rect 4488 2688 4494 2752
rect 4558 2688 4574 2752
rect 4638 2688 4654 2752
rect 4718 2688 4734 2752
rect 4798 2688 4804 2752
rect 4488 2687 4804 2688
rect 11572 2752 11888 2753
rect 11572 2688 11578 2752
rect 11642 2688 11658 2752
rect 11722 2688 11738 2752
rect 11802 2688 11818 2752
rect 11882 2688 11888 2752
rect 11572 2687 11888 2688
rect 18656 2752 18972 2753
rect 18656 2688 18662 2752
rect 18726 2688 18742 2752
rect 18806 2688 18822 2752
rect 18886 2688 18902 2752
rect 18966 2688 18972 2752
rect 18656 2687 18972 2688
rect 25740 2752 26056 2753
rect 25740 2688 25746 2752
rect 25810 2688 25826 2752
rect 25890 2688 25906 2752
rect 25970 2688 25986 2752
rect 26050 2688 26056 2752
rect 29821 2728 30621 2758
rect 25740 2687 26056 2688
rect 8030 2208 8346 2209
rect 0 2138 800 2168
rect 8030 2144 8036 2208
rect 8100 2144 8116 2208
rect 8180 2144 8196 2208
rect 8260 2144 8276 2208
rect 8340 2144 8346 2208
rect 8030 2143 8346 2144
rect 15114 2208 15430 2209
rect 15114 2144 15120 2208
rect 15184 2144 15200 2208
rect 15264 2144 15280 2208
rect 15344 2144 15360 2208
rect 15424 2144 15430 2208
rect 15114 2143 15430 2144
rect 22198 2208 22514 2209
rect 22198 2144 22204 2208
rect 22268 2144 22284 2208
rect 22348 2144 22364 2208
rect 22428 2144 22444 2208
rect 22508 2144 22514 2208
rect 22198 2143 22514 2144
rect 29282 2208 29598 2209
rect 29282 2144 29288 2208
rect 29352 2144 29368 2208
rect 29432 2144 29448 2208
rect 29512 2144 29528 2208
rect 29592 2144 29598 2208
rect 29282 2143 29598 2144
rect 1485 2138 1551 2141
rect 0 2136 1551 2138
rect 0 2080 1490 2136
rect 1546 2080 1551 2136
rect 0 2078 1551 2080
rect 0 2048 800 2078
rect 1485 2075 1551 2078
rect 27429 778 27495 781
rect 29821 778 30621 808
rect 27429 776 30621 778
rect 27429 720 27434 776
rect 27490 720 30621 776
rect 27429 718 30621 720
rect 27429 715 27495 718
rect 29821 688 30621 718
<< via3 >>
rect 8036 30492 8100 30496
rect 8036 30436 8040 30492
rect 8040 30436 8096 30492
rect 8096 30436 8100 30492
rect 8036 30432 8100 30436
rect 8116 30492 8180 30496
rect 8116 30436 8120 30492
rect 8120 30436 8176 30492
rect 8176 30436 8180 30492
rect 8116 30432 8180 30436
rect 8196 30492 8260 30496
rect 8196 30436 8200 30492
rect 8200 30436 8256 30492
rect 8256 30436 8260 30492
rect 8196 30432 8260 30436
rect 8276 30492 8340 30496
rect 8276 30436 8280 30492
rect 8280 30436 8336 30492
rect 8336 30436 8340 30492
rect 8276 30432 8340 30436
rect 15120 30492 15184 30496
rect 15120 30436 15124 30492
rect 15124 30436 15180 30492
rect 15180 30436 15184 30492
rect 15120 30432 15184 30436
rect 15200 30492 15264 30496
rect 15200 30436 15204 30492
rect 15204 30436 15260 30492
rect 15260 30436 15264 30492
rect 15200 30432 15264 30436
rect 15280 30492 15344 30496
rect 15280 30436 15284 30492
rect 15284 30436 15340 30492
rect 15340 30436 15344 30492
rect 15280 30432 15344 30436
rect 15360 30492 15424 30496
rect 15360 30436 15364 30492
rect 15364 30436 15420 30492
rect 15420 30436 15424 30492
rect 15360 30432 15424 30436
rect 22204 30492 22268 30496
rect 22204 30436 22208 30492
rect 22208 30436 22264 30492
rect 22264 30436 22268 30492
rect 22204 30432 22268 30436
rect 22284 30492 22348 30496
rect 22284 30436 22288 30492
rect 22288 30436 22344 30492
rect 22344 30436 22348 30492
rect 22284 30432 22348 30436
rect 22364 30492 22428 30496
rect 22364 30436 22368 30492
rect 22368 30436 22424 30492
rect 22424 30436 22428 30492
rect 22364 30432 22428 30436
rect 22444 30492 22508 30496
rect 22444 30436 22448 30492
rect 22448 30436 22504 30492
rect 22504 30436 22508 30492
rect 22444 30432 22508 30436
rect 29288 30492 29352 30496
rect 29288 30436 29292 30492
rect 29292 30436 29348 30492
rect 29348 30436 29352 30492
rect 29288 30432 29352 30436
rect 29368 30492 29432 30496
rect 29368 30436 29372 30492
rect 29372 30436 29428 30492
rect 29428 30436 29432 30492
rect 29368 30432 29432 30436
rect 29448 30492 29512 30496
rect 29448 30436 29452 30492
rect 29452 30436 29508 30492
rect 29508 30436 29512 30492
rect 29448 30432 29512 30436
rect 29528 30492 29592 30496
rect 29528 30436 29532 30492
rect 29532 30436 29588 30492
rect 29588 30436 29592 30492
rect 29528 30432 29592 30436
rect 4494 29948 4558 29952
rect 4494 29892 4498 29948
rect 4498 29892 4554 29948
rect 4554 29892 4558 29948
rect 4494 29888 4558 29892
rect 4574 29948 4638 29952
rect 4574 29892 4578 29948
rect 4578 29892 4634 29948
rect 4634 29892 4638 29948
rect 4574 29888 4638 29892
rect 4654 29948 4718 29952
rect 4654 29892 4658 29948
rect 4658 29892 4714 29948
rect 4714 29892 4718 29948
rect 4654 29888 4718 29892
rect 4734 29948 4798 29952
rect 4734 29892 4738 29948
rect 4738 29892 4794 29948
rect 4794 29892 4798 29948
rect 4734 29888 4798 29892
rect 11578 29948 11642 29952
rect 11578 29892 11582 29948
rect 11582 29892 11638 29948
rect 11638 29892 11642 29948
rect 11578 29888 11642 29892
rect 11658 29948 11722 29952
rect 11658 29892 11662 29948
rect 11662 29892 11718 29948
rect 11718 29892 11722 29948
rect 11658 29888 11722 29892
rect 11738 29948 11802 29952
rect 11738 29892 11742 29948
rect 11742 29892 11798 29948
rect 11798 29892 11802 29948
rect 11738 29888 11802 29892
rect 11818 29948 11882 29952
rect 11818 29892 11822 29948
rect 11822 29892 11878 29948
rect 11878 29892 11882 29948
rect 11818 29888 11882 29892
rect 18662 29948 18726 29952
rect 18662 29892 18666 29948
rect 18666 29892 18722 29948
rect 18722 29892 18726 29948
rect 18662 29888 18726 29892
rect 18742 29948 18806 29952
rect 18742 29892 18746 29948
rect 18746 29892 18802 29948
rect 18802 29892 18806 29948
rect 18742 29888 18806 29892
rect 18822 29948 18886 29952
rect 18822 29892 18826 29948
rect 18826 29892 18882 29948
rect 18882 29892 18886 29948
rect 18822 29888 18886 29892
rect 18902 29948 18966 29952
rect 18902 29892 18906 29948
rect 18906 29892 18962 29948
rect 18962 29892 18966 29948
rect 18902 29888 18966 29892
rect 25746 29948 25810 29952
rect 25746 29892 25750 29948
rect 25750 29892 25806 29948
rect 25806 29892 25810 29948
rect 25746 29888 25810 29892
rect 25826 29948 25890 29952
rect 25826 29892 25830 29948
rect 25830 29892 25886 29948
rect 25886 29892 25890 29948
rect 25826 29888 25890 29892
rect 25906 29948 25970 29952
rect 25906 29892 25910 29948
rect 25910 29892 25966 29948
rect 25966 29892 25970 29948
rect 25906 29888 25970 29892
rect 25986 29948 26050 29952
rect 25986 29892 25990 29948
rect 25990 29892 26046 29948
rect 26046 29892 26050 29948
rect 25986 29888 26050 29892
rect 8036 29404 8100 29408
rect 8036 29348 8040 29404
rect 8040 29348 8096 29404
rect 8096 29348 8100 29404
rect 8036 29344 8100 29348
rect 8116 29404 8180 29408
rect 8116 29348 8120 29404
rect 8120 29348 8176 29404
rect 8176 29348 8180 29404
rect 8116 29344 8180 29348
rect 8196 29404 8260 29408
rect 8196 29348 8200 29404
rect 8200 29348 8256 29404
rect 8256 29348 8260 29404
rect 8196 29344 8260 29348
rect 8276 29404 8340 29408
rect 8276 29348 8280 29404
rect 8280 29348 8336 29404
rect 8336 29348 8340 29404
rect 8276 29344 8340 29348
rect 15120 29404 15184 29408
rect 15120 29348 15124 29404
rect 15124 29348 15180 29404
rect 15180 29348 15184 29404
rect 15120 29344 15184 29348
rect 15200 29404 15264 29408
rect 15200 29348 15204 29404
rect 15204 29348 15260 29404
rect 15260 29348 15264 29404
rect 15200 29344 15264 29348
rect 15280 29404 15344 29408
rect 15280 29348 15284 29404
rect 15284 29348 15340 29404
rect 15340 29348 15344 29404
rect 15280 29344 15344 29348
rect 15360 29404 15424 29408
rect 15360 29348 15364 29404
rect 15364 29348 15420 29404
rect 15420 29348 15424 29404
rect 15360 29344 15424 29348
rect 22204 29404 22268 29408
rect 22204 29348 22208 29404
rect 22208 29348 22264 29404
rect 22264 29348 22268 29404
rect 22204 29344 22268 29348
rect 22284 29404 22348 29408
rect 22284 29348 22288 29404
rect 22288 29348 22344 29404
rect 22344 29348 22348 29404
rect 22284 29344 22348 29348
rect 22364 29404 22428 29408
rect 22364 29348 22368 29404
rect 22368 29348 22424 29404
rect 22424 29348 22428 29404
rect 22364 29344 22428 29348
rect 22444 29404 22508 29408
rect 22444 29348 22448 29404
rect 22448 29348 22504 29404
rect 22504 29348 22508 29404
rect 22444 29344 22508 29348
rect 29288 29404 29352 29408
rect 29288 29348 29292 29404
rect 29292 29348 29348 29404
rect 29348 29348 29352 29404
rect 29288 29344 29352 29348
rect 29368 29404 29432 29408
rect 29368 29348 29372 29404
rect 29372 29348 29428 29404
rect 29428 29348 29432 29404
rect 29368 29344 29432 29348
rect 29448 29404 29512 29408
rect 29448 29348 29452 29404
rect 29452 29348 29508 29404
rect 29508 29348 29512 29404
rect 29448 29344 29512 29348
rect 29528 29404 29592 29408
rect 29528 29348 29532 29404
rect 29532 29348 29588 29404
rect 29588 29348 29592 29404
rect 29528 29344 29592 29348
rect 27844 29276 27908 29340
rect 4494 28860 4558 28864
rect 4494 28804 4498 28860
rect 4498 28804 4554 28860
rect 4554 28804 4558 28860
rect 4494 28800 4558 28804
rect 4574 28860 4638 28864
rect 4574 28804 4578 28860
rect 4578 28804 4634 28860
rect 4634 28804 4638 28860
rect 4574 28800 4638 28804
rect 4654 28860 4718 28864
rect 4654 28804 4658 28860
rect 4658 28804 4714 28860
rect 4714 28804 4718 28860
rect 4654 28800 4718 28804
rect 4734 28860 4798 28864
rect 4734 28804 4738 28860
rect 4738 28804 4794 28860
rect 4794 28804 4798 28860
rect 4734 28800 4798 28804
rect 11578 28860 11642 28864
rect 11578 28804 11582 28860
rect 11582 28804 11638 28860
rect 11638 28804 11642 28860
rect 11578 28800 11642 28804
rect 11658 28860 11722 28864
rect 11658 28804 11662 28860
rect 11662 28804 11718 28860
rect 11718 28804 11722 28860
rect 11658 28800 11722 28804
rect 11738 28860 11802 28864
rect 11738 28804 11742 28860
rect 11742 28804 11798 28860
rect 11798 28804 11802 28860
rect 11738 28800 11802 28804
rect 11818 28860 11882 28864
rect 11818 28804 11822 28860
rect 11822 28804 11878 28860
rect 11878 28804 11882 28860
rect 11818 28800 11882 28804
rect 18662 28860 18726 28864
rect 18662 28804 18666 28860
rect 18666 28804 18722 28860
rect 18722 28804 18726 28860
rect 18662 28800 18726 28804
rect 18742 28860 18806 28864
rect 18742 28804 18746 28860
rect 18746 28804 18802 28860
rect 18802 28804 18806 28860
rect 18742 28800 18806 28804
rect 18822 28860 18886 28864
rect 18822 28804 18826 28860
rect 18826 28804 18882 28860
rect 18882 28804 18886 28860
rect 18822 28800 18886 28804
rect 18902 28860 18966 28864
rect 18902 28804 18906 28860
rect 18906 28804 18962 28860
rect 18962 28804 18966 28860
rect 18902 28800 18966 28804
rect 25746 28860 25810 28864
rect 25746 28804 25750 28860
rect 25750 28804 25806 28860
rect 25806 28804 25810 28860
rect 25746 28800 25810 28804
rect 25826 28860 25890 28864
rect 25826 28804 25830 28860
rect 25830 28804 25886 28860
rect 25886 28804 25890 28860
rect 25826 28800 25890 28804
rect 25906 28860 25970 28864
rect 25906 28804 25910 28860
rect 25910 28804 25966 28860
rect 25966 28804 25970 28860
rect 25906 28800 25970 28804
rect 25986 28860 26050 28864
rect 25986 28804 25990 28860
rect 25990 28804 26046 28860
rect 26046 28804 26050 28860
rect 25986 28800 26050 28804
rect 8036 28316 8100 28320
rect 8036 28260 8040 28316
rect 8040 28260 8096 28316
rect 8096 28260 8100 28316
rect 8036 28256 8100 28260
rect 8116 28316 8180 28320
rect 8116 28260 8120 28316
rect 8120 28260 8176 28316
rect 8176 28260 8180 28316
rect 8116 28256 8180 28260
rect 8196 28316 8260 28320
rect 8196 28260 8200 28316
rect 8200 28260 8256 28316
rect 8256 28260 8260 28316
rect 8196 28256 8260 28260
rect 8276 28316 8340 28320
rect 8276 28260 8280 28316
rect 8280 28260 8336 28316
rect 8336 28260 8340 28316
rect 8276 28256 8340 28260
rect 15120 28316 15184 28320
rect 15120 28260 15124 28316
rect 15124 28260 15180 28316
rect 15180 28260 15184 28316
rect 15120 28256 15184 28260
rect 15200 28316 15264 28320
rect 15200 28260 15204 28316
rect 15204 28260 15260 28316
rect 15260 28260 15264 28316
rect 15200 28256 15264 28260
rect 15280 28316 15344 28320
rect 15280 28260 15284 28316
rect 15284 28260 15340 28316
rect 15340 28260 15344 28316
rect 15280 28256 15344 28260
rect 15360 28316 15424 28320
rect 15360 28260 15364 28316
rect 15364 28260 15420 28316
rect 15420 28260 15424 28316
rect 15360 28256 15424 28260
rect 22204 28316 22268 28320
rect 22204 28260 22208 28316
rect 22208 28260 22264 28316
rect 22264 28260 22268 28316
rect 22204 28256 22268 28260
rect 22284 28316 22348 28320
rect 22284 28260 22288 28316
rect 22288 28260 22344 28316
rect 22344 28260 22348 28316
rect 22284 28256 22348 28260
rect 22364 28316 22428 28320
rect 22364 28260 22368 28316
rect 22368 28260 22424 28316
rect 22424 28260 22428 28316
rect 22364 28256 22428 28260
rect 22444 28316 22508 28320
rect 22444 28260 22448 28316
rect 22448 28260 22504 28316
rect 22504 28260 22508 28316
rect 22444 28256 22508 28260
rect 29288 28316 29352 28320
rect 29288 28260 29292 28316
rect 29292 28260 29348 28316
rect 29348 28260 29352 28316
rect 29288 28256 29352 28260
rect 29368 28316 29432 28320
rect 29368 28260 29372 28316
rect 29372 28260 29428 28316
rect 29428 28260 29432 28316
rect 29368 28256 29432 28260
rect 29448 28316 29512 28320
rect 29448 28260 29452 28316
rect 29452 28260 29508 28316
rect 29508 28260 29512 28316
rect 29448 28256 29512 28260
rect 29528 28316 29592 28320
rect 29528 28260 29532 28316
rect 29532 28260 29588 28316
rect 29588 28260 29592 28316
rect 29528 28256 29592 28260
rect 4494 27772 4558 27776
rect 4494 27716 4498 27772
rect 4498 27716 4554 27772
rect 4554 27716 4558 27772
rect 4494 27712 4558 27716
rect 4574 27772 4638 27776
rect 4574 27716 4578 27772
rect 4578 27716 4634 27772
rect 4634 27716 4638 27772
rect 4574 27712 4638 27716
rect 4654 27772 4718 27776
rect 4654 27716 4658 27772
rect 4658 27716 4714 27772
rect 4714 27716 4718 27772
rect 4654 27712 4718 27716
rect 4734 27772 4798 27776
rect 4734 27716 4738 27772
rect 4738 27716 4794 27772
rect 4794 27716 4798 27772
rect 4734 27712 4798 27716
rect 11578 27772 11642 27776
rect 11578 27716 11582 27772
rect 11582 27716 11638 27772
rect 11638 27716 11642 27772
rect 11578 27712 11642 27716
rect 11658 27772 11722 27776
rect 11658 27716 11662 27772
rect 11662 27716 11718 27772
rect 11718 27716 11722 27772
rect 11658 27712 11722 27716
rect 11738 27772 11802 27776
rect 11738 27716 11742 27772
rect 11742 27716 11798 27772
rect 11798 27716 11802 27772
rect 11738 27712 11802 27716
rect 11818 27772 11882 27776
rect 11818 27716 11822 27772
rect 11822 27716 11878 27772
rect 11878 27716 11882 27772
rect 11818 27712 11882 27716
rect 18662 27772 18726 27776
rect 18662 27716 18666 27772
rect 18666 27716 18722 27772
rect 18722 27716 18726 27772
rect 18662 27712 18726 27716
rect 18742 27772 18806 27776
rect 18742 27716 18746 27772
rect 18746 27716 18802 27772
rect 18802 27716 18806 27772
rect 18742 27712 18806 27716
rect 18822 27772 18886 27776
rect 18822 27716 18826 27772
rect 18826 27716 18882 27772
rect 18882 27716 18886 27772
rect 18822 27712 18886 27716
rect 18902 27772 18966 27776
rect 18902 27716 18906 27772
rect 18906 27716 18962 27772
rect 18962 27716 18966 27772
rect 18902 27712 18966 27716
rect 25746 27772 25810 27776
rect 25746 27716 25750 27772
rect 25750 27716 25806 27772
rect 25806 27716 25810 27772
rect 25746 27712 25810 27716
rect 25826 27772 25890 27776
rect 25826 27716 25830 27772
rect 25830 27716 25886 27772
rect 25886 27716 25890 27772
rect 25826 27712 25890 27716
rect 25906 27772 25970 27776
rect 25906 27716 25910 27772
rect 25910 27716 25966 27772
rect 25966 27716 25970 27772
rect 25906 27712 25970 27716
rect 25986 27772 26050 27776
rect 25986 27716 25990 27772
rect 25990 27716 26046 27772
rect 26046 27716 26050 27772
rect 25986 27712 26050 27716
rect 8036 27228 8100 27232
rect 8036 27172 8040 27228
rect 8040 27172 8096 27228
rect 8096 27172 8100 27228
rect 8036 27168 8100 27172
rect 8116 27228 8180 27232
rect 8116 27172 8120 27228
rect 8120 27172 8176 27228
rect 8176 27172 8180 27228
rect 8116 27168 8180 27172
rect 8196 27228 8260 27232
rect 8196 27172 8200 27228
rect 8200 27172 8256 27228
rect 8256 27172 8260 27228
rect 8196 27168 8260 27172
rect 8276 27228 8340 27232
rect 8276 27172 8280 27228
rect 8280 27172 8336 27228
rect 8336 27172 8340 27228
rect 8276 27168 8340 27172
rect 15120 27228 15184 27232
rect 15120 27172 15124 27228
rect 15124 27172 15180 27228
rect 15180 27172 15184 27228
rect 15120 27168 15184 27172
rect 15200 27228 15264 27232
rect 15200 27172 15204 27228
rect 15204 27172 15260 27228
rect 15260 27172 15264 27228
rect 15200 27168 15264 27172
rect 15280 27228 15344 27232
rect 15280 27172 15284 27228
rect 15284 27172 15340 27228
rect 15340 27172 15344 27228
rect 15280 27168 15344 27172
rect 15360 27228 15424 27232
rect 15360 27172 15364 27228
rect 15364 27172 15420 27228
rect 15420 27172 15424 27228
rect 15360 27168 15424 27172
rect 22204 27228 22268 27232
rect 22204 27172 22208 27228
rect 22208 27172 22264 27228
rect 22264 27172 22268 27228
rect 22204 27168 22268 27172
rect 22284 27228 22348 27232
rect 22284 27172 22288 27228
rect 22288 27172 22344 27228
rect 22344 27172 22348 27228
rect 22284 27168 22348 27172
rect 22364 27228 22428 27232
rect 22364 27172 22368 27228
rect 22368 27172 22424 27228
rect 22424 27172 22428 27228
rect 22364 27168 22428 27172
rect 22444 27228 22508 27232
rect 22444 27172 22448 27228
rect 22448 27172 22504 27228
rect 22504 27172 22508 27228
rect 22444 27168 22508 27172
rect 29288 27228 29352 27232
rect 29288 27172 29292 27228
rect 29292 27172 29348 27228
rect 29348 27172 29352 27228
rect 29288 27168 29352 27172
rect 29368 27228 29432 27232
rect 29368 27172 29372 27228
rect 29372 27172 29428 27228
rect 29428 27172 29432 27228
rect 29368 27168 29432 27172
rect 29448 27228 29512 27232
rect 29448 27172 29452 27228
rect 29452 27172 29508 27228
rect 29508 27172 29512 27228
rect 29448 27168 29512 27172
rect 29528 27228 29592 27232
rect 29528 27172 29532 27228
rect 29532 27172 29588 27228
rect 29588 27172 29592 27228
rect 29528 27168 29592 27172
rect 4494 26684 4558 26688
rect 4494 26628 4498 26684
rect 4498 26628 4554 26684
rect 4554 26628 4558 26684
rect 4494 26624 4558 26628
rect 4574 26684 4638 26688
rect 4574 26628 4578 26684
rect 4578 26628 4634 26684
rect 4634 26628 4638 26684
rect 4574 26624 4638 26628
rect 4654 26684 4718 26688
rect 4654 26628 4658 26684
rect 4658 26628 4714 26684
rect 4714 26628 4718 26684
rect 4654 26624 4718 26628
rect 4734 26684 4798 26688
rect 4734 26628 4738 26684
rect 4738 26628 4794 26684
rect 4794 26628 4798 26684
rect 4734 26624 4798 26628
rect 11578 26684 11642 26688
rect 11578 26628 11582 26684
rect 11582 26628 11638 26684
rect 11638 26628 11642 26684
rect 11578 26624 11642 26628
rect 11658 26684 11722 26688
rect 11658 26628 11662 26684
rect 11662 26628 11718 26684
rect 11718 26628 11722 26684
rect 11658 26624 11722 26628
rect 11738 26684 11802 26688
rect 11738 26628 11742 26684
rect 11742 26628 11798 26684
rect 11798 26628 11802 26684
rect 11738 26624 11802 26628
rect 11818 26684 11882 26688
rect 11818 26628 11822 26684
rect 11822 26628 11878 26684
rect 11878 26628 11882 26684
rect 11818 26624 11882 26628
rect 18662 26684 18726 26688
rect 18662 26628 18666 26684
rect 18666 26628 18722 26684
rect 18722 26628 18726 26684
rect 18662 26624 18726 26628
rect 18742 26684 18806 26688
rect 18742 26628 18746 26684
rect 18746 26628 18802 26684
rect 18802 26628 18806 26684
rect 18742 26624 18806 26628
rect 18822 26684 18886 26688
rect 18822 26628 18826 26684
rect 18826 26628 18882 26684
rect 18882 26628 18886 26684
rect 18822 26624 18886 26628
rect 18902 26684 18966 26688
rect 18902 26628 18906 26684
rect 18906 26628 18962 26684
rect 18962 26628 18966 26684
rect 18902 26624 18966 26628
rect 25746 26684 25810 26688
rect 25746 26628 25750 26684
rect 25750 26628 25806 26684
rect 25806 26628 25810 26684
rect 25746 26624 25810 26628
rect 25826 26684 25890 26688
rect 25826 26628 25830 26684
rect 25830 26628 25886 26684
rect 25886 26628 25890 26684
rect 25826 26624 25890 26628
rect 25906 26684 25970 26688
rect 25906 26628 25910 26684
rect 25910 26628 25966 26684
rect 25966 26628 25970 26684
rect 25906 26624 25970 26628
rect 25986 26684 26050 26688
rect 25986 26628 25990 26684
rect 25990 26628 26046 26684
rect 26046 26628 26050 26684
rect 25986 26624 26050 26628
rect 22692 26284 22756 26348
rect 8036 26140 8100 26144
rect 8036 26084 8040 26140
rect 8040 26084 8096 26140
rect 8096 26084 8100 26140
rect 8036 26080 8100 26084
rect 8116 26140 8180 26144
rect 8116 26084 8120 26140
rect 8120 26084 8176 26140
rect 8176 26084 8180 26140
rect 8116 26080 8180 26084
rect 8196 26140 8260 26144
rect 8196 26084 8200 26140
rect 8200 26084 8256 26140
rect 8256 26084 8260 26140
rect 8196 26080 8260 26084
rect 8276 26140 8340 26144
rect 8276 26084 8280 26140
rect 8280 26084 8336 26140
rect 8336 26084 8340 26140
rect 8276 26080 8340 26084
rect 15120 26140 15184 26144
rect 15120 26084 15124 26140
rect 15124 26084 15180 26140
rect 15180 26084 15184 26140
rect 15120 26080 15184 26084
rect 15200 26140 15264 26144
rect 15200 26084 15204 26140
rect 15204 26084 15260 26140
rect 15260 26084 15264 26140
rect 15200 26080 15264 26084
rect 15280 26140 15344 26144
rect 15280 26084 15284 26140
rect 15284 26084 15340 26140
rect 15340 26084 15344 26140
rect 15280 26080 15344 26084
rect 15360 26140 15424 26144
rect 15360 26084 15364 26140
rect 15364 26084 15420 26140
rect 15420 26084 15424 26140
rect 15360 26080 15424 26084
rect 22204 26140 22268 26144
rect 22204 26084 22208 26140
rect 22208 26084 22264 26140
rect 22264 26084 22268 26140
rect 22204 26080 22268 26084
rect 22284 26140 22348 26144
rect 22284 26084 22288 26140
rect 22288 26084 22344 26140
rect 22344 26084 22348 26140
rect 22284 26080 22348 26084
rect 22364 26140 22428 26144
rect 22364 26084 22368 26140
rect 22368 26084 22424 26140
rect 22424 26084 22428 26140
rect 22364 26080 22428 26084
rect 22444 26140 22508 26144
rect 22444 26084 22448 26140
rect 22448 26084 22504 26140
rect 22504 26084 22508 26140
rect 22444 26080 22508 26084
rect 29288 26140 29352 26144
rect 29288 26084 29292 26140
rect 29292 26084 29348 26140
rect 29348 26084 29352 26140
rect 29288 26080 29352 26084
rect 29368 26140 29432 26144
rect 29368 26084 29372 26140
rect 29372 26084 29428 26140
rect 29428 26084 29432 26140
rect 29368 26080 29432 26084
rect 29448 26140 29512 26144
rect 29448 26084 29452 26140
rect 29452 26084 29508 26140
rect 29508 26084 29512 26140
rect 29448 26080 29512 26084
rect 29528 26140 29592 26144
rect 29528 26084 29532 26140
rect 29532 26084 29588 26140
rect 29588 26084 29592 26140
rect 29528 26080 29592 26084
rect 4494 25596 4558 25600
rect 4494 25540 4498 25596
rect 4498 25540 4554 25596
rect 4554 25540 4558 25596
rect 4494 25536 4558 25540
rect 4574 25596 4638 25600
rect 4574 25540 4578 25596
rect 4578 25540 4634 25596
rect 4634 25540 4638 25596
rect 4574 25536 4638 25540
rect 4654 25596 4718 25600
rect 4654 25540 4658 25596
rect 4658 25540 4714 25596
rect 4714 25540 4718 25596
rect 4654 25536 4718 25540
rect 4734 25596 4798 25600
rect 4734 25540 4738 25596
rect 4738 25540 4794 25596
rect 4794 25540 4798 25596
rect 4734 25536 4798 25540
rect 11578 25596 11642 25600
rect 11578 25540 11582 25596
rect 11582 25540 11638 25596
rect 11638 25540 11642 25596
rect 11578 25536 11642 25540
rect 11658 25596 11722 25600
rect 11658 25540 11662 25596
rect 11662 25540 11718 25596
rect 11718 25540 11722 25596
rect 11658 25536 11722 25540
rect 11738 25596 11802 25600
rect 11738 25540 11742 25596
rect 11742 25540 11798 25596
rect 11798 25540 11802 25596
rect 11738 25536 11802 25540
rect 11818 25596 11882 25600
rect 11818 25540 11822 25596
rect 11822 25540 11878 25596
rect 11878 25540 11882 25596
rect 11818 25536 11882 25540
rect 18662 25596 18726 25600
rect 18662 25540 18666 25596
rect 18666 25540 18722 25596
rect 18722 25540 18726 25596
rect 18662 25536 18726 25540
rect 18742 25596 18806 25600
rect 18742 25540 18746 25596
rect 18746 25540 18802 25596
rect 18802 25540 18806 25596
rect 18742 25536 18806 25540
rect 18822 25596 18886 25600
rect 18822 25540 18826 25596
rect 18826 25540 18882 25596
rect 18882 25540 18886 25596
rect 18822 25536 18886 25540
rect 18902 25596 18966 25600
rect 18902 25540 18906 25596
rect 18906 25540 18962 25596
rect 18962 25540 18966 25596
rect 18902 25536 18966 25540
rect 25746 25596 25810 25600
rect 25746 25540 25750 25596
rect 25750 25540 25806 25596
rect 25806 25540 25810 25596
rect 25746 25536 25810 25540
rect 25826 25596 25890 25600
rect 25826 25540 25830 25596
rect 25830 25540 25886 25596
rect 25886 25540 25890 25596
rect 25826 25536 25890 25540
rect 25906 25596 25970 25600
rect 25906 25540 25910 25596
rect 25910 25540 25966 25596
rect 25966 25540 25970 25596
rect 25906 25536 25970 25540
rect 25986 25596 26050 25600
rect 25986 25540 25990 25596
rect 25990 25540 26046 25596
rect 26046 25540 26050 25596
rect 25986 25536 26050 25540
rect 8036 25052 8100 25056
rect 8036 24996 8040 25052
rect 8040 24996 8096 25052
rect 8096 24996 8100 25052
rect 8036 24992 8100 24996
rect 8116 25052 8180 25056
rect 8116 24996 8120 25052
rect 8120 24996 8176 25052
rect 8176 24996 8180 25052
rect 8116 24992 8180 24996
rect 8196 25052 8260 25056
rect 8196 24996 8200 25052
rect 8200 24996 8256 25052
rect 8256 24996 8260 25052
rect 8196 24992 8260 24996
rect 8276 25052 8340 25056
rect 8276 24996 8280 25052
rect 8280 24996 8336 25052
rect 8336 24996 8340 25052
rect 8276 24992 8340 24996
rect 15120 25052 15184 25056
rect 15120 24996 15124 25052
rect 15124 24996 15180 25052
rect 15180 24996 15184 25052
rect 15120 24992 15184 24996
rect 15200 25052 15264 25056
rect 15200 24996 15204 25052
rect 15204 24996 15260 25052
rect 15260 24996 15264 25052
rect 15200 24992 15264 24996
rect 15280 25052 15344 25056
rect 15280 24996 15284 25052
rect 15284 24996 15340 25052
rect 15340 24996 15344 25052
rect 15280 24992 15344 24996
rect 15360 25052 15424 25056
rect 15360 24996 15364 25052
rect 15364 24996 15420 25052
rect 15420 24996 15424 25052
rect 15360 24992 15424 24996
rect 22204 25052 22268 25056
rect 22204 24996 22208 25052
rect 22208 24996 22264 25052
rect 22264 24996 22268 25052
rect 22204 24992 22268 24996
rect 22284 25052 22348 25056
rect 22284 24996 22288 25052
rect 22288 24996 22344 25052
rect 22344 24996 22348 25052
rect 22284 24992 22348 24996
rect 22364 25052 22428 25056
rect 22364 24996 22368 25052
rect 22368 24996 22424 25052
rect 22424 24996 22428 25052
rect 22364 24992 22428 24996
rect 22444 25052 22508 25056
rect 22444 24996 22448 25052
rect 22448 24996 22504 25052
rect 22504 24996 22508 25052
rect 22444 24992 22508 24996
rect 29288 25052 29352 25056
rect 29288 24996 29292 25052
rect 29292 24996 29348 25052
rect 29348 24996 29352 25052
rect 29288 24992 29352 24996
rect 29368 25052 29432 25056
rect 29368 24996 29372 25052
rect 29372 24996 29428 25052
rect 29428 24996 29432 25052
rect 29368 24992 29432 24996
rect 29448 25052 29512 25056
rect 29448 24996 29452 25052
rect 29452 24996 29508 25052
rect 29508 24996 29512 25052
rect 29448 24992 29512 24996
rect 29528 25052 29592 25056
rect 29528 24996 29532 25052
rect 29532 24996 29588 25052
rect 29588 24996 29592 25052
rect 29528 24992 29592 24996
rect 4494 24508 4558 24512
rect 4494 24452 4498 24508
rect 4498 24452 4554 24508
rect 4554 24452 4558 24508
rect 4494 24448 4558 24452
rect 4574 24508 4638 24512
rect 4574 24452 4578 24508
rect 4578 24452 4634 24508
rect 4634 24452 4638 24508
rect 4574 24448 4638 24452
rect 4654 24508 4718 24512
rect 4654 24452 4658 24508
rect 4658 24452 4714 24508
rect 4714 24452 4718 24508
rect 4654 24448 4718 24452
rect 4734 24508 4798 24512
rect 4734 24452 4738 24508
rect 4738 24452 4794 24508
rect 4794 24452 4798 24508
rect 4734 24448 4798 24452
rect 11578 24508 11642 24512
rect 11578 24452 11582 24508
rect 11582 24452 11638 24508
rect 11638 24452 11642 24508
rect 11578 24448 11642 24452
rect 11658 24508 11722 24512
rect 11658 24452 11662 24508
rect 11662 24452 11718 24508
rect 11718 24452 11722 24508
rect 11658 24448 11722 24452
rect 11738 24508 11802 24512
rect 11738 24452 11742 24508
rect 11742 24452 11798 24508
rect 11798 24452 11802 24508
rect 11738 24448 11802 24452
rect 11818 24508 11882 24512
rect 11818 24452 11822 24508
rect 11822 24452 11878 24508
rect 11878 24452 11882 24508
rect 11818 24448 11882 24452
rect 18662 24508 18726 24512
rect 18662 24452 18666 24508
rect 18666 24452 18722 24508
rect 18722 24452 18726 24508
rect 18662 24448 18726 24452
rect 18742 24508 18806 24512
rect 18742 24452 18746 24508
rect 18746 24452 18802 24508
rect 18802 24452 18806 24508
rect 18742 24448 18806 24452
rect 18822 24508 18886 24512
rect 18822 24452 18826 24508
rect 18826 24452 18882 24508
rect 18882 24452 18886 24508
rect 18822 24448 18886 24452
rect 18902 24508 18966 24512
rect 18902 24452 18906 24508
rect 18906 24452 18962 24508
rect 18962 24452 18966 24508
rect 18902 24448 18966 24452
rect 25746 24508 25810 24512
rect 25746 24452 25750 24508
rect 25750 24452 25806 24508
rect 25806 24452 25810 24508
rect 25746 24448 25810 24452
rect 25826 24508 25890 24512
rect 25826 24452 25830 24508
rect 25830 24452 25886 24508
rect 25886 24452 25890 24508
rect 25826 24448 25890 24452
rect 25906 24508 25970 24512
rect 25906 24452 25910 24508
rect 25910 24452 25966 24508
rect 25966 24452 25970 24508
rect 25906 24448 25970 24452
rect 25986 24508 26050 24512
rect 25986 24452 25990 24508
rect 25990 24452 26046 24508
rect 26046 24452 26050 24508
rect 25986 24448 26050 24452
rect 8036 23964 8100 23968
rect 8036 23908 8040 23964
rect 8040 23908 8096 23964
rect 8096 23908 8100 23964
rect 8036 23904 8100 23908
rect 8116 23964 8180 23968
rect 8116 23908 8120 23964
rect 8120 23908 8176 23964
rect 8176 23908 8180 23964
rect 8116 23904 8180 23908
rect 8196 23964 8260 23968
rect 8196 23908 8200 23964
rect 8200 23908 8256 23964
rect 8256 23908 8260 23964
rect 8196 23904 8260 23908
rect 8276 23964 8340 23968
rect 8276 23908 8280 23964
rect 8280 23908 8336 23964
rect 8336 23908 8340 23964
rect 8276 23904 8340 23908
rect 15120 23964 15184 23968
rect 15120 23908 15124 23964
rect 15124 23908 15180 23964
rect 15180 23908 15184 23964
rect 15120 23904 15184 23908
rect 15200 23964 15264 23968
rect 15200 23908 15204 23964
rect 15204 23908 15260 23964
rect 15260 23908 15264 23964
rect 15200 23904 15264 23908
rect 15280 23964 15344 23968
rect 15280 23908 15284 23964
rect 15284 23908 15340 23964
rect 15340 23908 15344 23964
rect 15280 23904 15344 23908
rect 15360 23964 15424 23968
rect 15360 23908 15364 23964
rect 15364 23908 15420 23964
rect 15420 23908 15424 23964
rect 15360 23904 15424 23908
rect 22204 23964 22268 23968
rect 22204 23908 22208 23964
rect 22208 23908 22264 23964
rect 22264 23908 22268 23964
rect 22204 23904 22268 23908
rect 22284 23964 22348 23968
rect 22284 23908 22288 23964
rect 22288 23908 22344 23964
rect 22344 23908 22348 23964
rect 22284 23904 22348 23908
rect 22364 23964 22428 23968
rect 22364 23908 22368 23964
rect 22368 23908 22424 23964
rect 22424 23908 22428 23964
rect 22364 23904 22428 23908
rect 22444 23964 22508 23968
rect 22444 23908 22448 23964
rect 22448 23908 22504 23964
rect 22504 23908 22508 23964
rect 22444 23904 22508 23908
rect 29288 23964 29352 23968
rect 29288 23908 29292 23964
rect 29292 23908 29348 23964
rect 29348 23908 29352 23964
rect 29288 23904 29352 23908
rect 29368 23964 29432 23968
rect 29368 23908 29372 23964
rect 29372 23908 29428 23964
rect 29428 23908 29432 23964
rect 29368 23904 29432 23908
rect 29448 23964 29512 23968
rect 29448 23908 29452 23964
rect 29452 23908 29508 23964
rect 29508 23908 29512 23964
rect 29448 23904 29512 23908
rect 29528 23964 29592 23968
rect 29528 23908 29532 23964
rect 29532 23908 29588 23964
rect 29588 23908 29592 23964
rect 29528 23904 29592 23908
rect 4494 23420 4558 23424
rect 4494 23364 4498 23420
rect 4498 23364 4554 23420
rect 4554 23364 4558 23420
rect 4494 23360 4558 23364
rect 4574 23420 4638 23424
rect 4574 23364 4578 23420
rect 4578 23364 4634 23420
rect 4634 23364 4638 23420
rect 4574 23360 4638 23364
rect 4654 23420 4718 23424
rect 4654 23364 4658 23420
rect 4658 23364 4714 23420
rect 4714 23364 4718 23420
rect 4654 23360 4718 23364
rect 4734 23420 4798 23424
rect 4734 23364 4738 23420
rect 4738 23364 4794 23420
rect 4794 23364 4798 23420
rect 4734 23360 4798 23364
rect 11578 23420 11642 23424
rect 11578 23364 11582 23420
rect 11582 23364 11638 23420
rect 11638 23364 11642 23420
rect 11578 23360 11642 23364
rect 11658 23420 11722 23424
rect 11658 23364 11662 23420
rect 11662 23364 11718 23420
rect 11718 23364 11722 23420
rect 11658 23360 11722 23364
rect 11738 23420 11802 23424
rect 11738 23364 11742 23420
rect 11742 23364 11798 23420
rect 11798 23364 11802 23420
rect 11738 23360 11802 23364
rect 11818 23420 11882 23424
rect 11818 23364 11822 23420
rect 11822 23364 11878 23420
rect 11878 23364 11882 23420
rect 11818 23360 11882 23364
rect 18662 23420 18726 23424
rect 18662 23364 18666 23420
rect 18666 23364 18722 23420
rect 18722 23364 18726 23420
rect 18662 23360 18726 23364
rect 18742 23420 18806 23424
rect 18742 23364 18746 23420
rect 18746 23364 18802 23420
rect 18802 23364 18806 23420
rect 18742 23360 18806 23364
rect 18822 23420 18886 23424
rect 18822 23364 18826 23420
rect 18826 23364 18882 23420
rect 18882 23364 18886 23420
rect 18822 23360 18886 23364
rect 18902 23420 18966 23424
rect 18902 23364 18906 23420
rect 18906 23364 18962 23420
rect 18962 23364 18966 23420
rect 18902 23360 18966 23364
rect 25746 23420 25810 23424
rect 25746 23364 25750 23420
rect 25750 23364 25806 23420
rect 25806 23364 25810 23420
rect 25746 23360 25810 23364
rect 25826 23420 25890 23424
rect 25826 23364 25830 23420
rect 25830 23364 25886 23420
rect 25886 23364 25890 23420
rect 25826 23360 25890 23364
rect 25906 23420 25970 23424
rect 25906 23364 25910 23420
rect 25910 23364 25966 23420
rect 25966 23364 25970 23420
rect 25906 23360 25970 23364
rect 25986 23420 26050 23424
rect 25986 23364 25990 23420
rect 25990 23364 26046 23420
rect 26046 23364 26050 23420
rect 25986 23360 26050 23364
rect 21036 22944 21100 22948
rect 21036 22888 21086 22944
rect 21086 22888 21100 22944
rect 21036 22884 21100 22888
rect 8036 22876 8100 22880
rect 8036 22820 8040 22876
rect 8040 22820 8096 22876
rect 8096 22820 8100 22876
rect 8036 22816 8100 22820
rect 8116 22876 8180 22880
rect 8116 22820 8120 22876
rect 8120 22820 8176 22876
rect 8176 22820 8180 22876
rect 8116 22816 8180 22820
rect 8196 22876 8260 22880
rect 8196 22820 8200 22876
rect 8200 22820 8256 22876
rect 8256 22820 8260 22876
rect 8196 22816 8260 22820
rect 8276 22876 8340 22880
rect 8276 22820 8280 22876
rect 8280 22820 8336 22876
rect 8336 22820 8340 22876
rect 8276 22816 8340 22820
rect 15120 22876 15184 22880
rect 15120 22820 15124 22876
rect 15124 22820 15180 22876
rect 15180 22820 15184 22876
rect 15120 22816 15184 22820
rect 15200 22876 15264 22880
rect 15200 22820 15204 22876
rect 15204 22820 15260 22876
rect 15260 22820 15264 22876
rect 15200 22816 15264 22820
rect 15280 22876 15344 22880
rect 15280 22820 15284 22876
rect 15284 22820 15340 22876
rect 15340 22820 15344 22876
rect 15280 22816 15344 22820
rect 15360 22876 15424 22880
rect 15360 22820 15364 22876
rect 15364 22820 15420 22876
rect 15420 22820 15424 22876
rect 15360 22816 15424 22820
rect 22204 22876 22268 22880
rect 22204 22820 22208 22876
rect 22208 22820 22264 22876
rect 22264 22820 22268 22876
rect 22204 22816 22268 22820
rect 22284 22876 22348 22880
rect 22284 22820 22288 22876
rect 22288 22820 22344 22876
rect 22344 22820 22348 22876
rect 22284 22816 22348 22820
rect 22364 22876 22428 22880
rect 22364 22820 22368 22876
rect 22368 22820 22424 22876
rect 22424 22820 22428 22876
rect 22364 22816 22428 22820
rect 22444 22876 22508 22880
rect 22444 22820 22448 22876
rect 22448 22820 22504 22876
rect 22504 22820 22508 22876
rect 22444 22816 22508 22820
rect 29288 22876 29352 22880
rect 29288 22820 29292 22876
rect 29292 22820 29348 22876
rect 29348 22820 29352 22876
rect 29288 22816 29352 22820
rect 29368 22876 29432 22880
rect 29368 22820 29372 22876
rect 29372 22820 29428 22876
rect 29428 22820 29432 22876
rect 29368 22816 29432 22820
rect 29448 22876 29512 22880
rect 29448 22820 29452 22876
rect 29452 22820 29508 22876
rect 29508 22820 29512 22876
rect 29448 22816 29512 22820
rect 29528 22876 29592 22880
rect 29528 22820 29532 22876
rect 29532 22820 29588 22876
rect 29588 22820 29592 22876
rect 29528 22816 29592 22820
rect 4494 22332 4558 22336
rect 4494 22276 4498 22332
rect 4498 22276 4554 22332
rect 4554 22276 4558 22332
rect 4494 22272 4558 22276
rect 4574 22332 4638 22336
rect 4574 22276 4578 22332
rect 4578 22276 4634 22332
rect 4634 22276 4638 22332
rect 4574 22272 4638 22276
rect 4654 22332 4718 22336
rect 4654 22276 4658 22332
rect 4658 22276 4714 22332
rect 4714 22276 4718 22332
rect 4654 22272 4718 22276
rect 4734 22332 4798 22336
rect 4734 22276 4738 22332
rect 4738 22276 4794 22332
rect 4794 22276 4798 22332
rect 4734 22272 4798 22276
rect 11578 22332 11642 22336
rect 11578 22276 11582 22332
rect 11582 22276 11638 22332
rect 11638 22276 11642 22332
rect 11578 22272 11642 22276
rect 11658 22332 11722 22336
rect 11658 22276 11662 22332
rect 11662 22276 11718 22332
rect 11718 22276 11722 22332
rect 11658 22272 11722 22276
rect 11738 22332 11802 22336
rect 11738 22276 11742 22332
rect 11742 22276 11798 22332
rect 11798 22276 11802 22332
rect 11738 22272 11802 22276
rect 11818 22332 11882 22336
rect 11818 22276 11822 22332
rect 11822 22276 11878 22332
rect 11878 22276 11882 22332
rect 11818 22272 11882 22276
rect 18662 22332 18726 22336
rect 18662 22276 18666 22332
rect 18666 22276 18722 22332
rect 18722 22276 18726 22332
rect 18662 22272 18726 22276
rect 18742 22332 18806 22336
rect 18742 22276 18746 22332
rect 18746 22276 18802 22332
rect 18802 22276 18806 22332
rect 18742 22272 18806 22276
rect 18822 22332 18886 22336
rect 18822 22276 18826 22332
rect 18826 22276 18882 22332
rect 18882 22276 18886 22332
rect 18822 22272 18886 22276
rect 18902 22332 18966 22336
rect 18902 22276 18906 22332
rect 18906 22276 18962 22332
rect 18962 22276 18966 22332
rect 18902 22272 18966 22276
rect 25746 22332 25810 22336
rect 25746 22276 25750 22332
rect 25750 22276 25806 22332
rect 25806 22276 25810 22332
rect 25746 22272 25810 22276
rect 25826 22332 25890 22336
rect 25826 22276 25830 22332
rect 25830 22276 25886 22332
rect 25886 22276 25890 22332
rect 25826 22272 25890 22276
rect 25906 22332 25970 22336
rect 25906 22276 25910 22332
rect 25910 22276 25966 22332
rect 25966 22276 25970 22332
rect 25906 22272 25970 22276
rect 25986 22332 26050 22336
rect 25986 22276 25990 22332
rect 25990 22276 26046 22332
rect 26046 22276 26050 22332
rect 25986 22272 26050 22276
rect 8036 21788 8100 21792
rect 8036 21732 8040 21788
rect 8040 21732 8096 21788
rect 8096 21732 8100 21788
rect 8036 21728 8100 21732
rect 8116 21788 8180 21792
rect 8116 21732 8120 21788
rect 8120 21732 8176 21788
rect 8176 21732 8180 21788
rect 8116 21728 8180 21732
rect 8196 21788 8260 21792
rect 8196 21732 8200 21788
rect 8200 21732 8256 21788
rect 8256 21732 8260 21788
rect 8196 21728 8260 21732
rect 8276 21788 8340 21792
rect 8276 21732 8280 21788
rect 8280 21732 8336 21788
rect 8336 21732 8340 21788
rect 8276 21728 8340 21732
rect 15120 21788 15184 21792
rect 15120 21732 15124 21788
rect 15124 21732 15180 21788
rect 15180 21732 15184 21788
rect 15120 21728 15184 21732
rect 15200 21788 15264 21792
rect 15200 21732 15204 21788
rect 15204 21732 15260 21788
rect 15260 21732 15264 21788
rect 15200 21728 15264 21732
rect 15280 21788 15344 21792
rect 15280 21732 15284 21788
rect 15284 21732 15340 21788
rect 15340 21732 15344 21788
rect 15280 21728 15344 21732
rect 15360 21788 15424 21792
rect 15360 21732 15364 21788
rect 15364 21732 15420 21788
rect 15420 21732 15424 21788
rect 15360 21728 15424 21732
rect 22204 21788 22268 21792
rect 22204 21732 22208 21788
rect 22208 21732 22264 21788
rect 22264 21732 22268 21788
rect 22204 21728 22268 21732
rect 22284 21788 22348 21792
rect 22284 21732 22288 21788
rect 22288 21732 22344 21788
rect 22344 21732 22348 21788
rect 22284 21728 22348 21732
rect 22364 21788 22428 21792
rect 22364 21732 22368 21788
rect 22368 21732 22424 21788
rect 22424 21732 22428 21788
rect 22364 21728 22428 21732
rect 22444 21788 22508 21792
rect 22444 21732 22448 21788
rect 22448 21732 22504 21788
rect 22504 21732 22508 21788
rect 22444 21728 22508 21732
rect 29288 21788 29352 21792
rect 29288 21732 29292 21788
rect 29292 21732 29348 21788
rect 29348 21732 29352 21788
rect 29288 21728 29352 21732
rect 29368 21788 29432 21792
rect 29368 21732 29372 21788
rect 29372 21732 29428 21788
rect 29428 21732 29432 21788
rect 29368 21728 29432 21732
rect 29448 21788 29512 21792
rect 29448 21732 29452 21788
rect 29452 21732 29508 21788
rect 29508 21732 29512 21788
rect 29448 21728 29512 21732
rect 29528 21788 29592 21792
rect 29528 21732 29532 21788
rect 29532 21732 29588 21788
rect 29588 21732 29592 21788
rect 29528 21728 29592 21732
rect 4494 21244 4558 21248
rect 4494 21188 4498 21244
rect 4498 21188 4554 21244
rect 4554 21188 4558 21244
rect 4494 21184 4558 21188
rect 4574 21244 4638 21248
rect 4574 21188 4578 21244
rect 4578 21188 4634 21244
rect 4634 21188 4638 21244
rect 4574 21184 4638 21188
rect 4654 21244 4718 21248
rect 4654 21188 4658 21244
rect 4658 21188 4714 21244
rect 4714 21188 4718 21244
rect 4654 21184 4718 21188
rect 4734 21244 4798 21248
rect 4734 21188 4738 21244
rect 4738 21188 4794 21244
rect 4794 21188 4798 21244
rect 4734 21184 4798 21188
rect 11578 21244 11642 21248
rect 11578 21188 11582 21244
rect 11582 21188 11638 21244
rect 11638 21188 11642 21244
rect 11578 21184 11642 21188
rect 11658 21244 11722 21248
rect 11658 21188 11662 21244
rect 11662 21188 11718 21244
rect 11718 21188 11722 21244
rect 11658 21184 11722 21188
rect 11738 21244 11802 21248
rect 11738 21188 11742 21244
rect 11742 21188 11798 21244
rect 11798 21188 11802 21244
rect 11738 21184 11802 21188
rect 11818 21244 11882 21248
rect 11818 21188 11822 21244
rect 11822 21188 11878 21244
rect 11878 21188 11882 21244
rect 11818 21184 11882 21188
rect 18662 21244 18726 21248
rect 18662 21188 18666 21244
rect 18666 21188 18722 21244
rect 18722 21188 18726 21244
rect 18662 21184 18726 21188
rect 18742 21244 18806 21248
rect 18742 21188 18746 21244
rect 18746 21188 18802 21244
rect 18802 21188 18806 21244
rect 18742 21184 18806 21188
rect 18822 21244 18886 21248
rect 18822 21188 18826 21244
rect 18826 21188 18882 21244
rect 18882 21188 18886 21244
rect 18822 21184 18886 21188
rect 18902 21244 18966 21248
rect 18902 21188 18906 21244
rect 18906 21188 18962 21244
rect 18962 21188 18966 21244
rect 18902 21184 18966 21188
rect 25746 21244 25810 21248
rect 25746 21188 25750 21244
rect 25750 21188 25806 21244
rect 25806 21188 25810 21244
rect 25746 21184 25810 21188
rect 25826 21244 25890 21248
rect 25826 21188 25830 21244
rect 25830 21188 25886 21244
rect 25886 21188 25890 21244
rect 25826 21184 25890 21188
rect 25906 21244 25970 21248
rect 25906 21188 25910 21244
rect 25910 21188 25966 21244
rect 25966 21188 25970 21244
rect 25906 21184 25970 21188
rect 25986 21244 26050 21248
rect 25986 21188 25990 21244
rect 25990 21188 26046 21244
rect 26046 21188 26050 21244
rect 25986 21184 26050 21188
rect 8036 20700 8100 20704
rect 8036 20644 8040 20700
rect 8040 20644 8096 20700
rect 8096 20644 8100 20700
rect 8036 20640 8100 20644
rect 8116 20700 8180 20704
rect 8116 20644 8120 20700
rect 8120 20644 8176 20700
rect 8176 20644 8180 20700
rect 8116 20640 8180 20644
rect 8196 20700 8260 20704
rect 8196 20644 8200 20700
rect 8200 20644 8256 20700
rect 8256 20644 8260 20700
rect 8196 20640 8260 20644
rect 8276 20700 8340 20704
rect 8276 20644 8280 20700
rect 8280 20644 8336 20700
rect 8336 20644 8340 20700
rect 8276 20640 8340 20644
rect 15120 20700 15184 20704
rect 15120 20644 15124 20700
rect 15124 20644 15180 20700
rect 15180 20644 15184 20700
rect 15120 20640 15184 20644
rect 15200 20700 15264 20704
rect 15200 20644 15204 20700
rect 15204 20644 15260 20700
rect 15260 20644 15264 20700
rect 15200 20640 15264 20644
rect 15280 20700 15344 20704
rect 15280 20644 15284 20700
rect 15284 20644 15340 20700
rect 15340 20644 15344 20700
rect 15280 20640 15344 20644
rect 15360 20700 15424 20704
rect 15360 20644 15364 20700
rect 15364 20644 15420 20700
rect 15420 20644 15424 20700
rect 15360 20640 15424 20644
rect 22204 20700 22268 20704
rect 22204 20644 22208 20700
rect 22208 20644 22264 20700
rect 22264 20644 22268 20700
rect 22204 20640 22268 20644
rect 22284 20700 22348 20704
rect 22284 20644 22288 20700
rect 22288 20644 22344 20700
rect 22344 20644 22348 20700
rect 22284 20640 22348 20644
rect 22364 20700 22428 20704
rect 22364 20644 22368 20700
rect 22368 20644 22424 20700
rect 22424 20644 22428 20700
rect 22364 20640 22428 20644
rect 22444 20700 22508 20704
rect 22444 20644 22448 20700
rect 22448 20644 22504 20700
rect 22504 20644 22508 20700
rect 22444 20640 22508 20644
rect 29288 20700 29352 20704
rect 29288 20644 29292 20700
rect 29292 20644 29348 20700
rect 29348 20644 29352 20700
rect 29288 20640 29352 20644
rect 29368 20700 29432 20704
rect 29368 20644 29372 20700
rect 29372 20644 29428 20700
rect 29428 20644 29432 20700
rect 29368 20640 29432 20644
rect 29448 20700 29512 20704
rect 29448 20644 29452 20700
rect 29452 20644 29508 20700
rect 29508 20644 29512 20700
rect 29448 20640 29512 20644
rect 29528 20700 29592 20704
rect 29528 20644 29532 20700
rect 29532 20644 29588 20700
rect 29588 20644 29592 20700
rect 29528 20640 29592 20644
rect 4494 20156 4558 20160
rect 4494 20100 4498 20156
rect 4498 20100 4554 20156
rect 4554 20100 4558 20156
rect 4494 20096 4558 20100
rect 4574 20156 4638 20160
rect 4574 20100 4578 20156
rect 4578 20100 4634 20156
rect 4634 20100 4638 20156
rect 4574 20096 4638 20100
rect 4654 20156 4718 20160
rect 4654 20100 4658 20156
rect 4658 20100 4714 20156
rect 4714 20100 4718 20156
rect 4654 20096 4718 20100
rect 4734 20156 4798 20160
rect 4734 20100 4738 20156
rect 4738 20100 4794 20156
rect 4794 20100 4798 20156
rect 4734 20096 4798 20100
rect 11578 20156 11642 20160
rect 11578 20100 11582 20156
rect 11582 20100 11638 20156
rect 11638 20100 11642 20156
rect 11578 20096 11642 20100
rect 11658 20156 11722 20160
rect 11658 20100 11662 20156
rect 11662 20100 11718 20156
rect 11718 20100 11722 20156
rect 11658 20096 11722 20100
rect 11738 20156 11802 20160
rect 11738 20100 11742 20156
rect 11742 20100 11798 20156
rect 11798 20100 11802 20156
rect 11738 20096 11802 20100
rect 11818 20156 11882 20160
rect 11818 20100 11822 20156
rect 11822 20100 11878 20156
rect 11878 20100 11882 20156
rect 11818 20096 11882 20100
rect 18662 20156 18726 20160
rect 18662 20100 18666 20156
rect 18666 20100 18722 20156
rect 18722 20100 18726 20156
rect 18662 20096 18726 20100
rect 18742 20156 18806 20160
rect 18742 20100 18746 20156
rect 18746 20100 18802 20156
rect 18802 20100 18806 20156
rect 18742 20096 18806 20100
rect 18822 20156 18886 20160
rect 18822 20100 18826 20156
rect 18826 20100 18882 20156
rect 18882 20100 18886 20156
rect 18822 20096 18886 20100
rect 18902 20156 18966 20160
rect 18902 20100 18906 20156
rect 18906 20100 18962 20156
rect 18962 20100 18966 20156
rect 18902 20096 18966 20100
rect 25746 20156 25810 20160
rect 25746 20100 25750 20156
rect 25750 20100 25806 20156
rect 25806 20100 25810 20156
rect 25746 20096 25810 20100
rect 25826 20156 25890 20160
rect 25826 20100 25830 20156
rect 25830 20100 25886 20156
rect 25886 20100 25890 20156
rect 25826 20096 25890 20100
rect 25906 20156 25970 20160
rect 25906 20100 25910 20156
rect 25910 20100 25966 20156
rect 25966 20100 25970 20156
rect 25906 20096 25970 20100
rect 25986 20156 26050 20160
rect 25986 20100 25990 20156
rect 25990 20100 26046 20156
rect 26046 20100 26050 20156
rect 25986 20096 26050 20100
rect 8036 19612 8100 19616
rect 8036 19556 8040 19612
rect 8040 19556 8096 19612
rect 8096 19556 8100 19612
rect 8036 19552 8100 19556
rect 8116 19612 8180 19616
rect 8116 19556 8120 19612
rect 8120 19556 8176 19612
rect 8176 19556 8180 19612
rect 8116 19552 8180 19556
rect 8196 19612 8260 19616
rect 8196 19556 8200 19612
rect 8200 19556 8256 19612
rect 8256 19556 8260 19612
rect 8196 19552 8260 19556
rect 8276 19612 8340 19616
rect 8276 19556 8280 19612
rect 8280 19556 8336 19612
rect 8336 19556 8340 19612
rect 8276 19552 8340 19556
rect 15120 19612 15184 19616
rect 15120 19556 15124 19612
rect 15124 19556 15180 19612
rect 15180 19556 15184 19612
rect 15120 19552 15184 19556
rect 15200 19612 15264 19616
rect 15200 19556 15204 19612
rect 15204 19556 15260 19612
rect 15260 19556 15264 19612
rect 15200 19552 15264 19556
rect 15280 19612 15344 19616
rect 15280 19556 15284 19612
rect 15284 19556 15340 19612
rect 15340 19556 15344 19612
rect 15280 19552 15344 19556
rect 15360 19612 15424 19616
rect 15360 19556 15364 19612
rect 15364 19556 15420 19612
rect 15420 19556 15424 19612
rect 15360 19552 15424 19556
rect 22204 19612 22268 19616
rect 22204 19556 22208 19612
rect 22208 19556 22264 19612
rect 22264 19556 22268 19612
rect 22204 19552 22268 19556
rect 22284 19612 22348 19616
rect 22284 19556 22288 19612
rect 22288 19556 22344 19612
rect 22344 19556 22348 19612
rect 22284 19552 22348 19556
rect 22364 19612 22428 19616
rect 22364 19556 22368 19612
rect 22368 19556 22424 19612
rect 22424 19556 22428 19612
rect 22364 19552 22428 19556
rect 22444 19612 22508 19616
rect 22444 19556 22448 19612
rect 22448 19556 22504 19612
rect 22504 19556 22508 19612
rect 22444 19552 22508 19556
rect 29288 19612 29352 19616
rect 29288 19556 29292 19612
rect 29292 19556 29348 19612
rect 29348 19556 29352 19612
rect 29288 19552 29352 19556
rect 29368 19612 29432 19616
rect 29368 19556 29372 19612
rect 29372 19556 29428 19612
rect 29428 19556 29432 19612
rect 29368 19552 29432 19556
rect 29448 19612 29512 19616
rect 29448 19556 29452 19612
rect 29452 19556 29508 19612
rect 29508 19556 29512 19612
rect 29448 19552 29512 19556
rect 29528 19612 29592 19616
rect 29528 19556 29532 19612
rect 29532 19556 29588 19612
rect 29588 19556 29592 19612
rect 29528 19552 29592 19556
rect 4494 19068 4558 19072
rect 4494 19012 4498 19068
rect 4498 19012 4554 19068
rect 4554 19012 4558 19068
rect 4494 19008 4558 19012
rect 4574 19068 4638 19072
rect 4574 19012 4578 19068
rect 4578 19012 4634 19068
rect 4634 19012 4638 19068
rect 4574 19008 4638 19012
rect 4654 19068 4718 19072
rect 4654 19012 4658 19068
rect 4658 19012 4714 19068
rect 4714 19012 4718 19068
rect 4654 19008 4718 19012
rect 4734 19068 4798 19072
rect 4734 19012 4738 19068
rect 4738 19012 4794 19068
rect 4794 19012 4798 19068
rect 4734 19008 4798 19012
rect 11578 19068 11642 19072
rect 11578 19012 11582 19068
rect 11582 19012 11638 19068
rect 11638 19012 11642 19068
rect 11578 19008 11642 19012
rect 11658 19068 11722 19072
rect 11658 19012 11662 19068
rect 11662 19012 11718 19068
rect 11718 19012 11722 19068
rect 11658 19008 11722 19012
rect 11738 19068 11802 19072
rect 11738 19012 11742 19068
rect 11742 19012 11798 19068
rect 11798 19012 11802 19068
rect 11738 19008 11802 19012
rect 11818 19068 11882 19072
rect 11818 19012 11822 19068
rect 11822 19012 11878 19068
rect 11878 19012 11882 19068
rect 11818 19008 11882 19012
rect 18662 19068 18726 19072
rect 18662 19012 18666 19068
rect 18666 19012 18722 19068
rect 18722 19012 18726 19068
rect 18662 19008 18726 19012
rect 18742 19068 18806 19072
rect 18742 19012 18746 19068
rect 18746 19012 18802 19068
rect 18802 19012 18806 19068
rect 18742 19008 18806 19012
rect 18822 19068 18886 19072
rect 18822 19012 18826 19068
rect 18826 19012 18882 19068
rect 18882 19012 18886 19068
rect 18822 19008 18886 19012
rect 18902 19068 18966 19072
rect 18902 19012 18906 19068
rect 18906 19012 18962 19068
rect 18962 19012 18966 19068
rect 18902 19008 18966 19012
rect 25746 19068 25810 19072
rect 25746 19012 25750 19068
rect 25750 19012 25806 19068
rect 25806 19012 25810 19068
rect 25746 19008 25810 19012
rect 25826 19068 25890 19072
rect 25826 19012 25830 19068
rect 25830 19012 25886 19068
rect 25886 19012 25890 19068
rect 25826 19008 25890 19012
rect 25906 19068 25970 19072
rect 25906 19012 25910 19068
rect 25910 19012 25966 19068
rect 25966 19012 25970 19068
rect 25906 19008 25970 19012
rect 25986 19068 26050 19072
rect 25986 19012 25990 19068
rect 25990 19012 26046 19068
rect 26046 19012 26050 19068
rect 25986 19008 26050 19012
rect 8036 18524 8100 18528
rect 8036 18468 8040 18524
rect 8040 18468 8096 18524
rect 8096 18468 8100 18524
rect 8036 18464 8100 18468
rect 8116 18524 8180 18528
rect 8116 18468 8120 18524
rect 8120 18468 8176 18524
rect 8176 18468 8180 18524
rect 8116 18464 8180 18468
rect 8196 18524 8260 18528
rect 8196 18468 8200 18524
rect 8200 18468 8256 18524
rect 8256 18468 8260 18524
rect 8196 18464 8260 18468
rect 8276 18524 8340 18528
rect 8276 18468 8280 18524
rect 8280 18468 8336 18524
rect 8336 18468 8340 18524
rect 8276 18464 8340 18468
rect 15120 18524 15184 18528
rect 15120 18468 15124 18524
rect 15124 18468 15180 18524
rect 15180 18468 15184 18524
rect 15120 18464 15184 18468
rect 15200 18524 15264 18528
rect 15200 18468 15204 18524
rect 15204 18468 15260 18524
rect 15260 18468 15264 18524
rect 15200 18464 15264 18468
rect 15280 18524 15344 18528
rect 15280 18468 15284 18524
rect 15284 18468 15340 18524
rect 15340 18468 15344 18524
rect 15280 18464 15344 18468
rect 15360 18524 15424 18528
rect 15360 18468 15364 18524
rect 15364 18468 15420 18524
rect 15420 18468 15424 18524
rect 15360 18464 15424 18468
rect 22204 18524 22268 18528
rect 22204 18468 22208 18524
rect 22208 18468 22264 18524
rect 22264 18468 22268 18524
rect 22204 18464 22268 18468
rect 22284 18524 22348 18528
rect 22284 18468 22288 18524
rect 22288 18468 22344 18524
rect 22344 18468 22348 18524
rect 22284 18464 22348 18468
rect 22364 18524 22428 18528
rect 22364 18468 22368 18524
rect 22368 18468 22424 18524
rect 22424 18468 22428 18524
rect 22364 18464 22428 18468
rect 22444 18524 22508 18528
rect 22444 18468 22448 18524
rect 22448 18468 22504 18524
rect 22504 18468 22508 18524
rect 22444 18464 22508 18468
rect 29288 18524 29352 18528
rect 29288 18468 29292 18524
rect 29292 18468 29348 18524
rect 29348 18468 29352 18524
rect 29288 18464 29352 18468
rect 29368 18524 29432 18528
rect 29368 18468 29372 18524
rect 29372 18468 29428 18524
rect 29428 18468 29432 18524
rect 29368 18464 29432 18468
rect 29448 18524 29512 18528
rect 29448 18468 29452 18524
rect 29452 18468 29508 18524
rect 29508 18468 29512 18524
rect 29448 18464 29512 18468
rect 29528 18524 29592 18528
rect 29528 18468 29532 18524
rect 29532 18468 29588 18524
rect 29588 18468 29592 18524
rect 29528 18464 29592 18468
rect 4494 17980 4558 17984
rect 4494 17924 4498 17980
rect 4498 17924 4554 17980
rect 4554 17924 4558 17980
rect 4494 17920 4558 17924
rect 4574 17980 4638 17984
rect 4574 17924 4578 17980
rect 4578 17924 4634 17980
rect 4634 17924 4638 17980
rect 4574 17920 4638 17924
rect 4654 17980 4718 17984
rect 4654 17924 4658 17980
rect 4658 17924 4714 17980
rect 4714 17924 4718 17980
rect 4654 17920 4718 17924
rect 4734 17980 4798 17984
rect 4734 17924 4738 17980
rect 4738 17924 4794 17980
rect 4794 17924 4798 17980
rect 4734 17920 4798 17924
rect 11578 17980 11642 17984
rect 11578 17924 11582 17980
rect 11582 17924 11638 17980
rect 11638 17924 11642 17980
rect 11578 17920 11642 17924
rect 11658 17980 11722 17984
rect 11658 17924 11662 17980
rect 11662 17924 11718 17980
rect 11718 17924 11722 17980
rect 11658 17920 11722 17924
rect 11738 17980 11802 17984
rect 11738 17924 11742 17980
rect 11742 17924 11798 17980
rect 11798 17924 11802 17980
rect 11738 17920 11802 17924
rect 11818 17980 11882 17984
rect 11818 17924 11822 17980
rect 11822 17924 11878 17980
rect 11878 17924 11882 17980
rect 11818 17920 11882 17924
rect 18662 17980 18726 17984
rect 18662 17924 18666 17980
rect 18666 17924 18722 17980
rect 18722 17924 18726 17980
rect 18662 17920 18726 17924
rect 18742 17980 18806 17984
rect 18742 17924 18746 17980
rect 18746 17924 18802 17980
rect 18802 17924 18806 17980
rect 18742 17920 18806 17924
rect 18822 17980 18886 17984
rect 18822 17924 18826 17980
rect 18826 17924 18882 17980
rect 18882 17924 18886 17980
rect 18822 17920 18886 17924
rect 18902 17980 18966 17984
rect 18902 17924 18906 17980
rect 18906 17924 18962 17980
rect 18962 17924 18966 17980
rect 18902 17920 18966 17924
rect 25746 17980 25810 17984
rect 25746 17924 25750 17980
rect 25750 17924 25806 17980
rect 25806 17924 25810 17980
rect 25746 17920 25810 17924
rect 25826 17980 25890 17984
rect 25826 17924 25830 17980
rect 25830 17924 25886 17980
rect 25886 17924 25890 17980
rect 25826 17920 25890 17924
rect 25906 17980 25970 17984
rect 25906 17924 25910 17980
rect 25910 17924 25966 17980
rect 25966 17924 25970 17980
rect 25906 17920 25970 17924
rect 25986 17980 26050 17984
rect 25986 17924 25990 17980
rect 25990 17924 26046 17980
rect 26046 17924 26050 17980
rect 25986 17920 26050 17924
rect 8036 17436 8100 17440
rect 8036 17380 8040 17436
rect 8040 17380 8096 17436
rect 8096 17380 8100 17436
rect 8036 17376 8100 17380
rect 8116 17436 8180 17440
rect 8116 17380 8120 17436
rect 8120 17380 8176 17436
rect 8176 17380 8180 17436
rect 8116 17376 8180 17380
rect 8196 17436 8260 17440
rect 8196 17380 8200 17436
rect 8200 17380 8256 17436
rect 8256 17380 8260 17436
rect 8196 17376 8260 17380
rect 8276 17436 8340 17440
rect 8276 17380 8280 17436
rect 8280 17380 8336 17436
rect 8336 17380 8340 17436
rect 8276 17376 8340 17380
rect 15120 17436 15184 17440
rect 15120 17380 15124 17436
rect 15124 17380 15180 17436
rect 15180 17380 15184 17436
rect 15120 17376 15184 17380
rect 15200 17436 15264 17440
rect 15200 17380 15204 17436
rect 15204 17380 15260 17436
rect 15260 17380 15264 17436
rect 15200 17376 15264 17380
rect 15280 17436 15344 17440
rect 15280 17380 15284 17436
rect 15284 17380 15340 17436
rect 15340 17380 15344 17436
rect 15280 17376 15344 17380
rect 15360 17436 15424 17440
rect 15360 17380 15364 17436
rect 15364 17380 15420 17436
rect 15420 17380 15424 17436
rect 15360 17376 15424 17380
rect 22204 17436 22268 17440
rect 22204 17380 22208 17436
rect 22208 17380 22264 17436
rect 22264 17380 22268 17436
rect 22204 17376 22268 17380
rect 22284 17436 22348 17440
rect 22284 17380 22288 17436
rect 22288 17380 22344 17436
rect 22344 17380 22348 17436
rect 22284 17376 22348 17380
rect 22364 17436 22428 17440
rect 22364 17380 22368 17436
rect 22368 17380 22424 17436
rect 22424 17380 22428 17436
rect 22364 17376 22428 17380
rect 22444 17436 22508 17440
rect 22444 17380 22448 17436
rect 22448 17380 22504 17436
rect 22504 17380 22508 17436
rect 22444 17376 22508 17380
rect 29288 17436 29352 17440
rect 29288 17380 29292 17436
rect 29292 17380 29348 17436
rect 29348 17380 29352 17436
rect 29288 17376 29352 17380
rect 29368 17436 29432 17440
rect 29368 17380 29372 17436
rect 29372 17380 29428 17436
rect 29428 17380 29432 17436
rect 29368 17376 29432 17380
rect 29448 17436 29512 17440
rect 29448 17380 29452 17436
rect 29452 17380 29508 17436
rect 29508 17380 29512 17436
rect 29448 17376 29512 17380
rect 29528 17436 29592 17440
rect 29528 17380 29532 17436
rect 29532 17380 29588 17436
rect 29588 17380 29592 17436
rect 29528 17376 29592 17380
rect 4494 16892 4558 16896
rect 4494 16836 4498 16892
rect 4498 16836 4554 16892
rect 4554 16836 4558 16892
rect 4494 16832 4558 16836
rect 4574 16892 4638 16896
rect 4574 16836 4578 16892
rect 4578 16836 4634 16892
rect 4634 16836 4638 16892
rect 4574 16832 4638 16836
rect 4654 16892 4718 16896
rect 4654 16836 4658 16892
rect 4658 16836 4714 16892
rect 4714 16836 4718 16892
rect 4654 16832 4718 16836
rect 4734 16892 4798 16896
rect 4734 16836 4738 16892
rect 4738 16836 4794 16892
rect 4794 16836 4798 16892
rect 4734 16832 4798 16836
rect 11578 16892 11642 16896
rect 11578 16836 11582 16892
rect 11582 16836 11638 16892
rect 11638 16836 11642 16892
rect 11578 16832 11642 16836
rect 11658 16892 11722 16896
rect 11658 16836 11662 16892
rect 11662 16836 11718 16892
rect 11718 16836 11722 16892
rect 11658 16832 11722 16836
rect 11738 16892 11802 16896
rect 11738 16836 11742 16892
rect 11742 16836 11798 16892
rect 11798 16836 11802 16892
rect 11738 16832 11802 16836
rect 11818 16892 11882 16896
rect 11818 16836 11822 16892
rect 11822 16836 11878 16892
rect 11878 16836 11882 16892
rect 11818 16832 11882 16836
rect 18662 16892 18726 16896
rect 18662 16836 18666 16892
rect 18666 16836 18722 16892
rect 18722 16836 18726 16892
rect 18662 16832 18726 16836
rect 18742 16892 18806 16896
rect 18742 16836 18746 16892
rect 18746 16836 18802 16892
rect 18802 16836 18806 16892
rect 18742 16832 18806 16836
rect 18822 16892 18886 16896
rect 18822 16836 18826 16892
rect 18826 16836 18882 16892
rect 18882 16836 18886 16892
rect 18822 16832 18886 16836
rect 18902 16892 18966 16896
rect 18902 16836 18906 16892
rect 18906 16836 18962 16892
rect 18962 16836 18966 16892
rect 18902 16832 18966 16836
rect 25746 16892 25810 16896
rect 25746 16836 25750 16892
rect 25750 16836 25806 16892
rect 25806 16836 25810 16892
rect 25746 16832 25810 16836
rect 25826 16892 25890 16896
rect 25826 16836 25830 16892
rect 25830 16836 25886 16892
rect 25886 16836 25890 16892
rect 25826 16832 25890 16836
rect 25906 16892 25970 16896
rect 25906 16836 25910 16892
rect 25910 16836 25966 16892
rect 25966 16836 25970 16892
rect 25906 16832 25970 16836
rect 25986 16892 26050 16896
rect 25986 16836 25990 16892
rect 25990 16836 26046 16892
rect 26046 16836 26050 16892
rect 25986 16832 26050 16836
rect 20668 16688 20732 16692
rect 20668 16632 20682 16688
rect 20682 16632 20732 16688
rect 20668 16628 20732 16632
rect 8036 16348 8100 16352
rect 8036 16292 8040 16348
rect 8040 16292 8096 16348
rect 8096 16292 8100 16348
rect 8036 16288 8100 16292
rect 8116 16348 8180 16352
rect 8116 16292 8120 16348
rect 8120 16292 8176 16348
rect 8176 16292 8180 16348
rect 8116 16288 8180 16292
rect 8196 16348 8260 16352
rect 8196 16292 8200 16348
rect 8200 16292 8256 16348
rect 8256 16292 8260 16348
rect 8196 16288 8260 16292
rect 8276 16348 8340 16352
rect 8276 16292 8280 16348
rect 8280 16292 8336 16348
rect 8336 16292 8340 16348
rect 8276 16288 8340 16292
rect 15120 16348 15184 16352
rect 15120 16292 15124 16348
rect 15124 16292 15180 16348
rect 15180 16292 15184 16348
rect 15120 16288 15184 16292
rect 15200 16348 15264 16352
rect 15200 16292 15204 16348
rect 15204 16292 15260 16348
rect 15260 16292 15264 16348
rect 15200 16288 15264 16292
rect 15280 16348 15344 16352
rect 15280 16292 15284 16348
rect 15284 16292 15340 16348
rect 15340 16292 15344 16348
rect 15280 16288 15344 16292
rect 15360 16348 15424 16352
rect 15360 16292 15364 16348
rect 15364 16292 15420 16348
rect 15420 16292 15424 16348
rect 15360 16288 15424 16292
rect 22204 16348 22268 16352
rect 22204 16292 22208 16348
rect 22208 16292 22264 16348
rect 22264 16292 22268 16348
rect 22204 16288 22268 16292
rect 22284 16348 22348 16352
rect 22284 16292 22288 16348
rect 22288 16292 22344 16348
rect 22344 16292 22348 16348
rect 22284 16288 22348 16292
rect 22364 16348 22428 16352
rect 22364 16292 22368 16348
rect 22368 16292 22424 16348
rect 22424 16292 22428 16348
rect 22364 16288 22428 16292
rect 22444 16348 22508 16352
rect 22444 16292 22448 16348
rect 22448 16292 22504 16348
rect 22504 16292 22508 16348
rect 22444 16288 22508 16292
rect 29288 16348 29352 16352
rect 29288 16292 29292 16348
rect 29292 16292 29348 16348
rect 29348 16292 29352 16348
rect 29288 16288 29352 16292
rect 29368 16348 29432 16352
rect 29368 16292 29372 16348
rect 29372 16292 29428 16348
rect 29428 16292 29432 16348
rect 29368 16288 29432 16292
rect 29448 16348 29512 16352
rect 29448 16292 29452 16348
rect 29452 16292 29508 16348
rect 29508 16292 29512 16348
rect 29448 16288 29512 16292
rect 29528 16348 29592 16352
rect 29528 16292 29532 16348
rect 29532 16292 29588 16348
rect 29588 16292 29592 16348
rect 29528 16288 29592 16292
rect 4494 15804 4558 15808
rect 4494 15748 4498 15804
rect 4498 15748 4554 15804
rect 4554 15748 4558 15804
rect 4494 15744 4558 15748
rect 4574 15804 4638 15808
rect 4574 15748 4578 15804
rect 4578 15748 4634 15804
rect 4634 15748 4638 15804
rect 4574 15744 4638 15748
rect 4654 15804 4718 15808
rect 4654 15748 4658 15804
rect 4658 15748 4714 15804
rect 4714 15748 4718 15804
rect 4654 15744 4718 15748
rect 4734 15804 4798 15808
rect 4734 15748 4738 15804
rect 4738 15748 4794 15804
rect 4794 15748 4798 15804
rect 4734 15744 4798 15748
rect 11578 15804 11642 15808
rect 11578 15748 11582 15804
rect 11582 15748 11638 15804
rect 11638 15748 11642 15804
rect 11578 15744 11642 15748
rect 11658 15804 11722 15808
rect 11658 15748 11662 15804
rect 11662 15748 11718 15804
rect 11718 15748 11722 15804
rect 11658 15744 11722 15748
rect 11738 15804 11802 15808
rect 11738 15748 11742 15804
rect 11742 15748 11798 15804
rect 11798 15748 11802 15804
rect 11738 15744 11802 15748
rect 11818 15804 11882 15808
rect 11818 15748 11822 15804
rect 11822 15748 11878 15804
rect 11878 15748 11882 15804
rect 11818 15744 11882 15748
rect 18662 15804 18726 15808
rect 18662 15748 18666 15804
rect 18666 15748 18722 15804
rect 18722 15748 18726 15804
rect 18662 15744 18726 15748
rect 18742 15804 18806 15808
rect 18742 15748 18746 15804
rect 18746 15748 18802 15804
rect 18802 15748 18806 15804
rect 18742 15744 18806 15748
rect 18822 15804 18886 15808
rect 18822 15748 18826 15804
rect 18826 15748 18882 15804
rect 18882 15748 18886 15804
rect 18822 15744 18886 15748
rect 18902 15804 18966 15808
rect 18902 15748 18906 15804
rect 18906 15748 18962 15804
rect 18962 15748 18966 15804
rect 18902 15744 18966 15748
rect 25746 15804 25810 15808
rect 25746 15748 25750 15804
rect 25750 15748 25806 15804
rect 25806 15748 25810 15804
rect 25746 15744 25810 15748
rect 25826 15804 25890 15808
rect 25826 15748 25830 15804
rect 25830 15748 25886 15804
rect 25886 15748 25890 15804
rect 25826 15744 25890 15748
rect 25906 15804 25970 15808
rect 25906 15748 25910 15804
rect 25910 15748 25966 15804
rect 25966 15748 25970 15804
rect 25906 15744 25970 15748
rect 25986 15804 26050 15808
rect 25986 15748 25990 15804
rect 25990 15748 26046 15804
rect 26046 15748 26050 15804
rect 25986 15744 26050 15748
rect 8036 15260 8100 15264
rect 8036 15204 8040 15260
rect 8040 15204 8096 15260
rect 8096 15204 8100 15260
rect 8036 15200 8100 15204
rect 8116 15260 8180 15264
rect 8116 15204 8120 15260
rect 8120 15204 8176 15260
rect 8176 15204 8180 15260
rect 8116 15200 8180 15204
rect 8196 15260 8260 15264
rect 8196 15204 8200 15260
rect 8200 15204 8256 15260
rect 8256 15204 8260 15260
rect 8196 15200 8260 15204
rect 8276 15260 8340 15264
rect 8276 15204 8280 15260
rect 8280 15204 8336 15260
rect 8336 15204 8340 15260
rect 8276 15200 8340 15204
rect 15120 15260 15184 15264
rect 15120 15204 15124 15260
rect 15124 15204 15180 15260
rect 15180 15204 15184 15260
rect 15120 15200 15184 15204
rect 15200 15260 15264 15264
rect 15200 15204 15204 15260
rect 15204 15204 15260 15260
rect 15260 15204 15264 15260
rect 15200 15200 15264 15204
rect 15280 15260 15344 15264
rect 15280 15204 15284 15260
rect 15284 15204 15340 15260
rect 15340 15204 15344 15260
rect 15280 15200 15344 15204
rect 15360 15260 15424 15264
rect 15360 15204 15364 15260
rect 15364 15204 15420 15260
rect 15420 15204 15424 15260
rect 15360 15200 15424 15204
rect 22204 15260 22268 15264
rect 22204 15204 22208 15260
rect 22208 15204 22264 15260
rect 22264 15204 22268 15260
rect 22204 15200 22268 15204
rect 22284 15260 22348 15264
rect 22284 15204 22288 15260
rect 22288 15204 22344 15260
rect 22344 15204 22348 15260
rect 22284 15200 22348 15204
rect 22364 15260 22428 15264
rect 22364 15204 22368 15260
rect 22368 15204 22424 15260
rect 22424 15204 22428 15260
rect 22364 15200 22428 15204
rect 22444 15260 22508 15264
rect 22444 15204 22448 15260
rect 22448 15204 22504 15260
rect 22504 15204 22508 15260
rect 22444 15200 22508 15204
rect 29288 15260 29352 15264
rect 29288 15204 29292 15260
rect 29292 15204 29348 15260
rect 29348 15204 29352 15260
rect 29288 15200 29352 15204
rect 29368 15260 29432 15264
rect 29368 15204 29372 15260
rect 29372 15204 29428 15260
rect 29428 15204 29432 15260
rect 29368 15200 29432 15204
rect 29448 15260 29512 15264
rect 29448 15204 29452 15260
rect 29452 15204 29508 15260
rect 29508 15204 29512 15260
rect 29448 15200 29512 15204
rect 29528 15260 29592 15264
rect 29528 15204 29532 15260
rect 29532 15204 29588 15260
rect 29588 15204 29592 15260
rect 29528 15200 29592 15204
rect 4494 14716 4558 14720
rect 4494 14660 4498 14716
rect 4498 14660 4554 14716
rect 4554 14660 4558 14716
rect 4494 14656 4558 14660
rect 4574 14716 4638 14720
rect 4574 14660 4578 14716
rect 4578 14660 4634 14716
rect 4634 14660 4638 14716
rect 4574 14656 4638 14660
rect 4654 14716 4718 14720
rect 4654 14660 4658 14716
rect 4658 14660 4714 14716
rect 4714 14660 4718 14716
rect 4654 14656 4718 14660
rect 4734 14716 4798 14720
rect 4734 14660 4738 14716
rect 4738 14660 4794 14716
rect 4794 14660 4798 14716
rect 4734 14656 4798 14660
rect 11578 14716 11642 14720
rect 11578 14660 11582 14716
rect 11582 14660 11638 14716
rect 11638 14660 11642 14716
rect 11578 14656 11642 14660
rect 11658 14716 11722 14720
rect 11658 14660 11662 14716
rect 11662 14660 11718 14716
rect 11718 14660 11722 14716
rect 11658 14656 11722 14660
rect 11738 14716 11802 14720
rect 11738 14660 11742 14716
rect 11742 14660 11798 14716
rect 11798 14660 11802 14716
rect 11738 14656 11802 14660
rect 11818 14716 11882 14720
rect 11818 14660 11822 14716
rect 11822 14660 11878 14716
rect 11878 14660 11882 14716
rect 11818 14656 11882 14660
rect 18662 14716 18726 14720
rect 18662 14660 18666 14716
rect 18666 14660 18722 14716
rect 18722 14660 18726 14716
rect 18662 14656 18726 14660
rect 18742 14716 18806 14720
rect 18742 14660 18746 14716
rect 18746 14660 18802 14716
rect 18802 14660 18806 14716
rect 18742 14656 18806 14660
rect 18822 14716 18886 14720
rect 18822 14660 18826 14716
rect 18826 14660 18882 14716
rect 18882 14660 18886 14716
rect 18822 14656 18886 14660
rect 18902 14716 18966 14720
rect 18902 14660 18906 14716
rect 18906 14660 18962 14716
rect 18962 14660 18966 14716
rect 18902 14656 18966 14660
rect 25746 14716 25810 14720
rect 25746 14660 25750 14716
rect 25750 14660 25806 14716
rect 25806 14660 25810 14716
rect 25746 14656 25810 14660
rect 25826 14716 25890 14720
rect 25826 14660 25830 14716
rect 25830 14660 25886 14716
rect 25886 14660 25890 14716
rect 25826 14656 25890 14660
rect 25906 14716 25970 14720
rect 25906 14660 25910 14716
rect 25910 14660 25966 14716
rect 25966 14660 25970 14716
rect 25906 14656 25970 14660
rect 25986 14716 26050 14720
rect 25986 14660 25990 14716
rect 25990 14660 26046 14716
rect 26046 14660 26050 14716
rect 25986 14656 26050 14660
rect 8036 14172 8100 14176
rect 8036 14116 8040 14172
rect 8040 14116 8096 14172
rect 8096 14116 8100 14172
rect 8036 14112 8100 14116
rect 8116 14172 8180 14176
rect 8116 14116 8120 14172
rect 8120 14116 8176 14172
rect 8176 14116 8180 14172
rect 8116 14112 8180 14116
rect 8196 14172 8260 14176
rect 8196 14116 8200 14172
rect 8200 14116 8256 14172
rect 8256 14116 8260 14172
rect 8196 14112 8260 14116
rect 8276 14172 8340 14176
rect 8276 14116 8280 14172
rect 8280 14116 8336 14172
rect 8336 14116 8340 14172
rect 8276 14112 8340 14116
rect 15120 14172 15184 14176
rect 15120 14116 15124 14172
rect 15124 14116 15180 14172
rect 15180 14116 15184 14172
rect 15120 14112 15184 14116
rect 15200 14172 15264 14176
rect 15200 14116 15204 14172
rect 15204 14116 15260 14172
rect 15260 14116 15264 14172
rect 15200 14112 15264 14116
rect 15280 14172 15344 14176
rect 15280 14116 15284 14172
rect 15284 14116 15340 14172
rect 15340 14116 15344 14172
rect 15280 14112 15344 14116
rect 15360 14172 15424 14176
rect 15360 14116 15364 14172
rect 15364 14116 15420 14172
rect 15420 14116 15424 14172
rect 15360 14112 15424 14116
rect 22204 14172 22268 14176
rect 22204 14116 22208 14172
rect 22208 14116 22264 14172
rect 22264 14116 22268 14172
rect 22204 14112 22268 14116
rect 22284 14172 22348 14176
rect 22284 14116 22288 14172
rect 22288 14116 22344 14172
rect 22344 14116 22348 14172
rect 22284 14112 22348 14116
rect 22364 14172 22428 14176
rect 22364 14116 22368 14172
rect 22368 14116 22424 14172
rect 22424 14116 22428 14172
rect 22364 14112 22428 14116
rect 22444 14172 22508 14176
rect 22444 14116 22448 14172
rect 22448 14116 22504 14172
rect 22504 14116 22508 14172
rect 22444 14112 22508 14116
rect 29288 14172 29352 14176
rect 29288 14116 29292 14172
rect 29292 14116 29348 14172
rect 29348 14116 29352 14172
rect 29288 14112 29352 14116
rect 29368 14172 29432 14176
rect 29368 14116 29372 14172
rect 29372 14116 29428 14172
rect 29428 14116 29432 14172
rect 29368 14112 29432 14116
rect 29448 14172 29512 14176
rect 29448 14116 29452 14172
rect 29452 14116 29508 14172
rect 29508 14116 29512 14172
rect 29448 14112 29512 14116
rect 29528 14172 29592 14176
rect 29528 14116 29532 14172
rect 29532 14116 29588 14172
rect 29588 14116 29592 14172
rect 29528 14112 29592 14116
rect 4494 13628 4558 13632
rect 4494 13572 4498 13628
rect 4498 13572 4554 13628
rect 4554 13572 4558 13628
rect 4494 13568 4558 13572
rect 4574 13628 4638 13632
rect 4574 13572 4578 13628
rect 4578 13572 4634 13628
rect 4634 13572 4638 13628
rect 4574 13568 4638 13572
rect 4654 13628 4718 13632
rect 4654 13572 4658 13628
rect 4658 13572 4714 13628
rect 4714 13572 4718 13628
rect 4654 13568 4718 13572
rect 4734 13628 4798 13632
rect 4734 13572 4738 13628
rect 4738 13572 4794 13628
rect 4794 13572 4798 13628
rect 4734 13568 4798 13572
rect 11578 13628 11642 13632
rect 11578 13572 11582 13628
rect 11582 13572 11638 13628
rect 11638 13572 11642 13628
rect 11578 13568 11642 13572
rect 11658 13628 11722 13632
rect 11658 13572 11662 13628
rect 11662 13572 11718 13628
rect 11718 13572 11722 13628
rect 11658 13568 11722 13572
rect 11738 13628 11802 13632
rect 11738 13572 11742 13628
rect 11742 13572 11798 13628
rect 11798 13572 11802 13628
rect 11738 13568 11802 13572
rect 11818 13628 11882 13632
rect 11818 13572 11822 13628
rect 11822 13572 11878 13628
rect 11878 13572 11882 13628
rect 11818 13568 11882 13572
rect 18662 13628 18726 13632
rect 18662 13572 18666 13628
rect 18666 13572 18722 13628
rect 18722 13572 18726 13628
rect 18662 13568 18726 13572
rect 18742 13628 18806 13632
rect 18742 13572 18746 13628
rect 18746 13572 18802 13628
rect 18802 13572 18806 13628
rect 18742 13568 18806 13572
rect 18822 13628 18886 13632
rect 18822 13572 18826 13628
rect 18826 13572 18882 13628
rect 18882 13572 18886 13628
rect 18822 13568 18886 13572
rect 18902 13628 18966 13632
rect 18902 13572 18906 13628
rect 18906 13572 18962 13628
rect 18962 13572 18966 13628
rect 18902 13568 18966 13572
rect 25746 13628 25810 13632
rect 25746 13572 25750 13628
rect 25750 13572 25806 13628
rect 25806 13572 25810 13628
rect 25746 13568 25810 13572
rect 25826 13628 25890 13632
rect 25826 13572 25830 13628
rect 25830 13572 25886 13628
rect 25886 13572 25890 13628
rect 25826 13568 25890 13572
rect 25906 13628 25970 13632
rect 25906 13572 25910 13628
rect 25910 13572 25966 13628
rect 25966 13572 25970 13628
rect 25906 13568 25970 13572
rect 25986 13628 26050 13632
rect 25986 13572 25990 13628
rect 25990 13572 26046 13628
rect 26046 13572 26050 13628
rect 25986 13568 26050 13572
rect 8036 13084 8100 13088
rect 8036 13028 8040 13084
rect 8040 13028 8096 13084
rect 8096 13028 8100 13084
rect 8036 13024 8100 13028
rect 8116 13084 8180 13088
rect 8116 13028 8120 13084
rect 8120 13028 8176 13084
rect 8176 13028 8180 13084
rect 8116 13024 8180 13028
rect 8196 13084 8260 13088
rect 8196 13028 8200 13084
rect 8200 13028 8256 13084
rect 8256 13028 8260 13084
rect 8196 13024 8260 13028
rect 8276 13084 8340 13088
rect 8276 13028 8280 13084
rect 8280 13028 8336 13084
rect 8336 13028 8340 13084
rect 8276 13024 8340 13028
rect 15120 13084 15184 13088
rect 15120 13028 15124 13084
rect 15124 13028 15180 13084
rect 15180 13028 15184 13084
rect 15120 13024 15184 13028
rect 15200 13084 15264 13088
rect 15200 13028 15204 13084
rect 15204 13028 15260 13084
rect 15260 13028 15264 13084
rect 15200 13024 15264 13028
rect 15280 13084 15344 13088
rect 15280 13028 15284 13084
rect 15284 13028 15340 13084
rect 15340 13028 15344 13084
rect 15280 13024 15344 13028
rect 15360 13084 15424 13088
rect 15360 13028 15364 13084
rect 15364 13028 15420 13084
rect 15420 13028 15424 13084
rect 15360 13024 15424 13028
rect 22204 13084 22268 13088
rect 22204 13028 22208 13084
rect 22208 13028 22264 13084
rect 22264 13028 22268 13084
rect 22204 13024 22268 13028
rect 22284 13084 22348 13088
rect 22284 13028 22288 13084
rect 22288 13028 22344 13084
rect 22344 13028 22348 13084
rect 22284 13024 22348 13028
rect 22364 13084 22428 13088
rect 22364 13028 22368 13084
rect 22368 13028 22424 13084
rect 22424 13028 22428 13084
rect 22364 13024 22428 13028
rect 22444 13084 22508 13088
rect 22444 13028 22448 13084
rect 22448 13028 22504 13084
rect 22504 13028 22508 13084
rect 22444 13024 22508 13028
rect 29288 13084 29352 13088
rect 29288 13028 29292 13084
rect 29292 13028 29348 13084
rect 29348 13028 29352 13084
rect 29288 13024 29352 13028
rect 29368 13084 29432 13088
rect 29368 13028 29372 13084
rect 29372 13028 29428 13084
rect 29428 13028 29432 13084
rect 29368 13024 29432 13028
rect 29448 13084 29512 13088
rect 29448 13028 29452 13084
rect 29452 13028 29508 13084
rect 29508 13028 29512 13084
rect 29448 13024 29512 13028
rect 29528 13084 29592 13088
rect 29528 13028 29532 13084
rect 29532 13028 29588 13084
rect 29588 13028 29592 13084
rect 29528 13024 29592 13028
rect 21036 12956 21100 13020
rect 4494 12540 4558 12544
rect 4494 12484 4498 12540
rect 4498 12484 4554 12540
rect 4554 12484 4558 12540
rect 4494 12480 4558 12484
rect 4574 12540 4638 12544
rect 4574 12484 4578 12540
rect 4578 12484 4634 12540
rect 4634 12484 4638 12540
rect 4574 12480 4638 12484
rect 4654 12540 4718 12544
rect 4654 12484 4658 12540
rect 4658 12484 4714 12540
rect 4714 12484 4718 12540
rect 4654 12480 4718 12484
rect 4734 12540 4798 12544
rect 4734 12484 4738 12540
rect 4738 12484 4794 12540
rect 4794 12484 4798 12540
rect 4734 12480 4798 12484
rect 11578 12540 11642 12544
rect 11578 12484 11582 12540
rect 11582 12484 11638 12540
rect 11638 12484 11642 12540
rect 11578 12480 11642 12484
rect 11658 12540 11722 12544
rect 11658 12484 11662 12540
rect 11662 12484 11718 12540
rect 11718 12484 11722 12540
rect 11658 12480 11722 12484
rect 11738 12540 11802 12544
rect 11738 12484 11742 12540
rect 11742 12484 11798 12540
rect 11798 12484 11802 12540
rect 11738 12480 11802 12484
rect 11818 12540 11882 12544
rect 11818 12484 11822 12540
rect 11822 12484 11878 12540
rect 11878 12484 11882 12540
rect 11818 12480 11882 12484
rect 18662 12540 18726 12544
rect 18662 12484 18666 12540
rect 18666 12484 18722 12540
rect 18722 12484 18726 12540
rect 18662 12480 18726 12484
rect 18742 12540 18806 12544
rect 18742 12484 18746 12540
rect 18746 12484 18802 12540
rect 18802 12484 18806 12540
rect 18742 12480 18806 12484
rect 18822 12540 18886 12544
rect 18822 12484 18826 12540
rect 18826 12484 18882 12540
rect 18882 12484 18886 12540
rect 18822 12480 18886 12484
rect 18902 12540 18966 12544
rect 18902 12484 18906 12540
rect 18906 12484 18962 12540
rect 18962 12484 18966 12540
rect 18902 12480 18966 12484
rect 25746 12540 25810 12544
rect 25746 12484 25750 12540
rect 25750 12484 25806 12540
rect 25806 12484 25810 12540
rect 25746 12480 25810 12484
rect 25826 12540 25890 12544
rect 25826 12484 25830 12540
rect 25830 12484 25886 12540
rect 25886 12484 25890 12540
rect 25826 12480 25890 12484
rect 25906 12540 25970 12544
rect 25906 12484 25910 12540
rect 25910 12484 25966 12540
rect 25966 12484 25970 12540
rect 25906 12480 25970 12484
rect 25986 12540 26050 12544
rect 25986 12484 25990 12540
rect 25990 12484 26046 12540
rect 26046 12484 26050 12540
rect 25986 12480 26050 12484
rect 20668 12140 20732 12204
rect 8036 11996 8100 12000
rect 8036 11940 8040 11996
rect 8040 11940 8096 11996
rect 8096 11940 8100 11996
rect 8036 11936 8100 11940
rect 8116 11996 8180 12000
rect 8116 11940 8120 11996
rect 8120 11940 8176 11996
rect 8176 11940 8180 11996
rect 8116 11936 8180 11940
rect 8196 11996 8260 12000
rect 8196 11940 8200 11996
rect 8200 11940 8256 11996
rect 8256 11940 8260 11996
rect 8196 11936 8260 11940
rect 8276 11996 8340 12000
rect 8276 11940 8280 11996
rect 8280 11940 8336 11996
rect 8336 11940 8340 11996
rect 8276 11936 8340 11940
rect 15120 11996 15184 12000
rect 15120 11940 15124 11996
rect 15124 11940 15180 11996
rect 15180 11940 15184 11996
rect 15120 11936 15184 11940
rect 15200 11996 15264 12000
rect 15200 11940 15204 11996
rect 15204 11940 15260 11996
rect 15260 11940 15264 11996
rect 15200 11936 15264 11940
rect 15280 11996 15344 12000
rect 15280 11940 15284 11996
rect 15284 11940 15340 11996
rect 15340 11940 15344 11996
rect 15280 11936 15344 11940
rect 15360 11996 15424 12000
rect 15360 11940 15364 11996
rect 15364 11940 15420 11996
rect 15420 11940 15424 11996
rect 15360 11936 15424 11940
rect 22204 11996 22268 12000
rect 22204 11940 22208 11996
rect 22208 11940 22264 11996
rect 22264 11940 22268 11996
rect 22204 11936 22268 11940
rect 22284 11996 22348 12000
rect 22284 11940 22288 11996
rect 22288 11940 22344 11996
rect 22344 11940 22348 11996
rect 22284 11936 22348 11940
rect 22364 11996 22428 12000
rect 22364 11940 22368 11996
rect 22368 11940 22424 11996
rect 22424 11940 22428 11996
rect 22364 11936 22428 11940
rect 22444 11996 22508 12000
rect 22444 11940 22448 11996
rect 22448 11940 22504 11996
rect 22504 11940 22508 11996
rect 22444 11936 22508 11940
rect 29288 11996 29352 12000
rect 29288 11940 29292 11996
rect 29292 11940 29348 11996
rect 29348 11940 29352 11996
rect 29288 11936 29352 11940
rect 29368 11996 29432 12000
rect 29368 11940 29372 11996
rect 29372 11940 29428 11996
rect 29428 11940 29432 11996
rect 29368 11936 29432 11940
rect 29448 11996 29512 12000
rect 29448 11940 29452 11996
rect 29452 11940 29508 11996
rect 29508 11940 29512 11996
rect 29448 11936 29512 11940
rect 29528 11996 29592 12000
rect 29528 11940 29532 11996
rect 29532 11940 29588 11996
rect 29588 11940 29592 11996
rect 29528 11936 29592 11940
rect 4494 11452 4558 11456
rect 4494 11396 4498 11452
rect 4498 11396 4554 11452
rect 4554 11396 4558 11452
rect 4494 11392 4558 11396
rect 4574 11452 4638 11456
rect 4574 11396 4578 11452
rect 4578 11396 4634 11452
rect 4634 11396 4638 11452
rect 4574 11392 4638 11396
rect 4654 11452 4718 11456
rect 4654 11396 4658 11452
rect 4658 11396 4714 11452
rect 4714 11396 4718 11452
rect 4654 11392 4718 11396
rect 4734 11452 4798 11456
rect 4734 11396 4738 11452
rect 4738 11396 4794 11452
rect 4794 11396 4798 11452
rect 4734 11392 4798 11396
rect 11578 11452 11642 11456
rect 11578 11396 11582 11452
rect 11582 11396 11638 11452
rect 11638 11396 11642 11452
rect 11578 11392 11642 11396
rect 11658 11452 11722 11456
rect 11658 11396 11662 11452
rect 11662 11396 11718 11452
rect 11718 11396 11722 11452
rect 11658 11392 11722 11396
rect 11738 11452 11802 11456
rect 11738 11396 11742 11452
rect 11742 11396 11798 11452
rect 11798 11396 11802 11452
rect 11738 11392 11802 11396
rect 11818 11452 11882 11456
rect 11818 11396 11822 11452
rect 11822 11396 11878 11452
rect 11878 11396 11882 11452
rect 11818 11392 11882 11396
rect 18662 11452 18726 11456
rect 18662 11396 18666 11452
rect 18666 11396 18722 11452
rect 18722 11396 18726 11452
rect 18662 11392 18726 11396
rect 18742 11452 18806 11456
rect 18742 11396 18746 11452
rect 18746 11396 18802 11452
rect 18802 11396 18806 11452
rect 18742 11392 18806 11396
rect 18822 11452 18886 11456
rect 18822 11396 18826 11452
rect 18826 11396 18882 11452
rect 18882 11396 18886 11452
rect 18822 11392 18886 11396
rect 18902 11452 18966 11456
rect 18902 11396 18906 11452
rect 18906 11396 18962 11452
rect 18962 11396 18966 11452
rect 18902 11392 18966 11396
rect 25746 11452 25810 11456
rect 25746 11396 25750 11452
rect 25750 11396 25806 11452
rect 25806 11396 25810 11452
rect 25746 11392 25810 11396
rect 25826 11452 25890 11456
rect 25826 11396 25830 11452
rect 25830 11396 25886 11452
rect 25886 11396 25890 11452
rect 25826 11392 25890 11396
rect 25906 11452 25970 11456
rect 25906 11396 25910 11452
rect 25910 11396 25966 11452
rect 25966 11396 25970 11452
rect 25906 11392 25970 11396
rect 25986 11452 26050 11456
rect 25986 11396 25990 11452
rect 25990 11396 26046 11452
rect 26046 11396 26050 11452
rect 25986 11392 26050 11396
rect 8036 10908 8100 10912
rect 8036 10852 8040 10908
rect 8040 10852 8096 10908
rect 8096 10852 8100 10908
rect 8036 10848 8100 10852
rect 8116 10908 8180 10912
rect 8116 10852 8120 10908
rect 8120 10852 8176 10908
rect 8176 10852 8180 10908
rect 8116 10848 8180 10852
rect 8196 10908 8260 10912
rect 8196 10852 8200 10908
rect 8200 10852 8256 10908
rect 8256 10852 8260 10908
rect 8196 10848 8260 10852
rect 8276 10908 8340 10912
rect 8276 10852 8280 10908
rect 8280 10852 8336 10908
rect 8336 10852 8340 10908
rect 8276 10848 8340 10852
rect 15120 10908 15184 10912
rect 15120 10852 15124 10908
rect 15124 10852 15180 10908
rect 15180 10852 15184 10908
rect 15120 10848 15184 10852
rect 15200 10908 15264 10912
rect 15200 10852 15204 10908
rect 15204 10852 15260 10908
rect 15260 10852 15264 10908
rect 15200 10848 15264 10852
rect 15280 10908 15344 10912
rect 15280 10852 15284 10908
rect 15284 10852 15340 10908
rect 15340 10852 15344 10908
rect 15280 10848 15344 10852
rect 15360 10908 15424 10912
rect 15360 10852 15364 10908
rect 15364 10852 15420 10908
rect 15420 10852 15424 10908
rect 15360 10848 15424 10852
rect 22204 10908 22268 10912
rect 22204 10852 22208 10908
rect 22208 10852 22264 10908
rect 22264 10852 22268 10908
rect 22204 10848 22268 10852
rect 22284 10908 22348 10912
rect 22284 10852 22288 10908
rect 22288 10852 22344 10908
rect 22344 10852 22348 10908
rect 22284 10848 22348 10852
rect 22364 10908 22428 10912
rect 22364 10852 22368 10908
rect 22368 10852 22424 10908
rect 22424 10852 22428 10908
rect 22364 10848 22428 10852
rect 22444 10908 22508 10912
rect 22444 10852 22448 10908
rect 22448 10852 22504 10908
rect 22504 10852 22508 10908
rect 22444 10848 22508 10852
rect 29288 10908 29352 10912
rect 29288 10852 29292 10908
rect 29292 10852 29348 10908
rect 29348 10852 29352 10908
rect 29288 10848 29352 10852
rect 29368 10908 29432 10912
rect 29368 10852 29372 10908
rect 29372 10852 29428 10908
rect 29428 10852 29432 10908
rect 29368 10848 29432 10852
rect 29448 10908 29512 10912
rect 29448 10852 29452 10908
rect 29452 10852 29508 10908
rect 29508 10852 29512 10908
rect 29448 10848 29512 10852
rect 29528 10908 29592 10912
rect 29528 10852 29532 10908
rect 29532 10852 29588 10908
rect 29588 10852 29592 10908
rect 29528 10848 29592 10852
rect 4494 10364 4558 10368
rect 4494 10308 4498 10364
rect 4498 10308 4554 10364
rect 4554 10308 4558 10364
rect 4494 10304 4558 10308
rect 4574 10364 4638 10368
rect 4574 10308 4578 10364
rect 4578 10308 4634 10364
rect 4634 10308 4638 10364
rect 4574 10304 4638 10308
rect 4654 10364 4718 10368
rect 4654 10308 4658 10364
rect 4658 10308 4714 10364
rect 4714 10308 4718 10364
rect 4654 10304 4718 10308
rect 4734 10364 4798 10368
rect 4734 10308 4738 10364
rect 4738 10308 4794 10364
rect 4794 10308 4798 10364
rect 4734 10304 4798 10308
rect 11578 10364 11642 10368
rect 11578 10308 11582 10364
rect 11582 10308 11638 10364
rect 11638 10308 11642 10364
rect 11578 10304 11642 10308
rect 11658 10364 11722 10368
rect 11658 10308 11662 10364
rect 11662 10308 11718 10364
rect 11718 10308 11722 10364
rect 11658 10304 11722 10308
rect 11738 10364 11802 10368
rect 11738 10308 11742 10364
rect 11742 10308 11798 10364
rect 11798 10308 11802 10364
rect 11738 10304 11802 10308
rect 11818 10364 11882 10368
rect 11818 10308 11822 10364
rect 11822 10308 11878 10364
rect 11878 10308 11882 10364
rect 11818 10304 11882 10308
rect 18662 10364 18726 10368
rect 18662 10308 18666 10364
rect 18666 10308 18722 10364
rect 18722 10308 18726 10364
rect 18662 10304 18726 10308
rect 18742 10364 18806 10368
rect 18742 10308 18746 10364
rect 18746 10308 18802 10364
rect 18802 10308 18806 10364
rect 18742 10304 18806 10308
rect 18822 10364 18886 10368
rect 18822 10308 18826 10364
rect 18826 10308 18882 10364
rect 18882 10308 18886 10364
rect 18822 10304 18886 10308
rect 18902 10364 18966 10368
rect 18902 10308 18906 10364
rect 18906 10308 18962 10364
rect 18962 10308 18966 10364
rect 18902 10304 18966 10308
rect 25746 10364 25810 10368
rect 25746 10308 25750 10364
rect 25750 10308 25806 10364
rect 25806 10308 25810 10364
rect 25746 10304 25810 10308
rect 25826 10364 25890 10368
rect 25826 10308 25830 10364
rect 25830 10308 25886 10364
rect 25886 10308 25890 10364
rect 25826 10304 25890 10308
rect 25906 10364 25970 10368
rect 25906 10308 25910 10364
rect 25910 10308 25966 10364
rect 25966 10308 25970 10364
rect 25906 10304 25970 10308
rect 25986 10364 26050 10368
rect 25986 10308 25990 10364
rect 25990 10308 26046 10364
rect 26046 10308 26050 10364
rect 25986 10304 26050 10308
rect 8036 9820 8100 9824
rect 8036 9764 8040 9820
rect 8040 9764 8096 9820
rect 8096 9764 8100 9820
rect 8036 9760 8100 9764
rect 8116 9820 8180 9824
rect 8116 9764 8120 9820
rect 8120 9764 8176 9820
rect 8176 9764 8180 9820
rect 8116 9760 8180 9764
rect 8196 9820 8260 9824
rect 8196 9764 8200 9820
rect 8200 9764 8256 9820
rect 8256 9764 8260 9820
rect 8196 9760 8260 9764
rect 8276 9820 8340 9824
rect 8276 9764 8280 9820
rect 8280 9764 8336 9820
rect 8336 9764 8340 9820
rect 8276 9760 8340 9764
rect 15120 9820 15184 9824
rect 15120 9764 15124 9820
rect 15124 9764 15180 9820
rect 15180 9764 15184 9820
rect 15120 9760 15184 9764
rect 15200 9820 15264 9824
rect 15200 9764 15204 9820
rect 15204 9764 15260 9820
rect 15260 9764 15264 9820
rect 15200 9760 15264 9764
rect 15280 9820 15344 9824
rect 15280 9764 15284 9820
rect 15284 9764 15340 9820
rect 15340 9764 15344 9820
rect 15280 9760 15344 9764
rect 15360 9820 15424 9824
rect 15360 9764 15364 9820
rect 15364 9764 15420 9820
rect 15420 9764 15424 9820
rect 15360 9760 15424 9764
rect 22204 9820 22268 9824
rect 22204 9764 22208 9820
rect 22208 9764 22264 9820
rect 22264 9764 22268 9820
rect 22204 9760 22268 9764
rect 22284 9820 22348 9824
rect 22284 9764 22288 9820
rect 22288 9764 22344 9820
rect 22344 9764 22348 9820
rect 22284 9760 22348 9764
rect 22364 9820 22428 9824
rect 22364 9764 22368 9820
rect 22368 9764 22424 9820
rect 22424 9764 22428 9820
rect 22364 9760 22428 9764
rect 22444 9820 22508 9824
rect 22444 9764 22448 9820
rect 22448 9764 22504 9820
rect 22504 9764 22508 9820
rect 22444 9760 22508 9764
rect 29288 9820 29352 9824
rect 29288 9764 29292 9820
rect 29292 9764 29348 9820
rect 29348 9764 29352 9820
rect 29288 9760 29352 9764
rect 29368 9820 29432 9824
rect 29368 9764 29372 9820
rect 29372 9764 29428 9820
rect 29428 9764 29432 9820
rect 29368 9760 29432 9764
rect 29448 9820 29512 9824
rect 29448 9764 29452 9820
rect 29452 9764 29508 9820
rect 29508 9764 29512 9820
rect 29448 9760 29512 9764
rect 29528 9820 29592 9824
rect 29528 9764 29532 9820
rect 29532 9764 29588 9820
rect 29588 9764 29592 9820
rect 29528 9760 29592 9764
rect 4494 9276 4558 9280
rect 4494 9220 4498 9276
rect 4498 9220 4554 9276
rect 4554 9220 4558 9276
rect 4494 9216 4558 9220
rect 4574 9276 4638 9280
rect 4574 9220 4578 9276
rect 4578 9220 4634 9276
rect 4634 9220 4638 9276
rect 4574 9216 4638 9220
rect 4654 9276 4718 9280
rect 4654 9220 4658 9276
rect 4658 9220 4714 9276
rect 4714 9220 4718 9276
rect 4654 9216 4718 9220
rect 4734 9276 4798 9280
rect 4734 9220 4738 9276
rect 4738 9220 4794 9276
rect 4794 9220 4798 9276
rect 4734 9216 4798 9220
rect 11578 9276 11642 9280
rect 11578 9220 11582 9276
rect 11582 9220 11638 9276
rect 11638 9220 11642 9276
rect 11578 9216 11642 9220
rect 11658 9276 11722 9280
rect 11658 9220 11662 9276
rect 11662 9220 11718 9276
rect 11718 9220 11722 9276
rect 11658 9216 11722 9220
rect 11738 9276 11802 9280
rect 11738 9220 11742 9276
rect 11742 9220 11798 9276
rect 11798 9220 11802 9276
rect 11738 9216 11802 9220
rect 11818 9276 11882 9280
rect 11818 9220 11822 9276
rect 11822 9220 11878 9276
rect 11878 9220 11882 9276
rect 11818 9216 11882 9220
rect 18662 9276 18726 9280
rect 18662 9220 18666 9276
rect 18666 9220 18722 9276
rect 18722 9220 18726 9276
rect 18662 9216 18726 9220
rect 18742 9276 18806 9280
rect 18742 9220 18746 9276
rect 18746 9220 18802 9276
rect 18802 9220 18806 9276
rect 18742 9216 18806 9220
rect 18822 9276 18886 9280
rect 18822 9220 18826 9276
rect 18826 9220 18882 9276
rect 18882 9220 18886 9276
rect 18822 9216 18886 9220
rect 18902 9276 18966 9280
rect 18902 9220 18906 9276
rect 18906 9220 18962 9276
rect 18962 9220 18966 9276
rect 18902 9216 18966 9220
rect 25746 9276 25810 9280
rect 25746 9220 25750 9276
rect 25750 9220 25806 9276
rect 25806 9220 25810 9276
rect 25746 9216 25810 9220
rect 25826 9276 25890 9280
rect 25826 9220 25830 9276
rect 25830 9220 25886 9276
rect 25886 9220 25890 9276
rect 25826 9216 25890 9220
rect 25906 9276 25970 9280
rect 25906 9220 25910 9276
rect 25910 9220 25966 9276
rect 25966 9220 25970 9276
rect 25906 9216 25970 9220
rect 25986 9276 26050 9280
rect 25986 9220 25990 9276
rect 25990 9220 26046 9276
rect 26046 9220 26050 9276
rect 25986 9216 26050 9220
rect 8036 8732 8100 8736
rect 8036 8676 8040 8732
rect 8040 8676 8096 8732
rect 8096 8676 8100 8732
rect 8036 8672 8100 8676
rect 8116 8732 8180 8736
rect 8116 8676 8120 8732
rect 8120 8676 8176 8732
rect 8176 8676 8180 8732
rect 8116 8672 8180 8676
rect 8196 8732 8260 8736
rect 8196 8676 8200 8732
rect 8200 8676 8256 8732
rect 8256 8676 8260 8732
rect 8196 8672 8260 8676
rect 8276 8732 8340 8736
rect 8276 8676 8280 8732
rect 8280 8676 8336 8732
rect 8336 8676 8340 8732
rect 8276 8672 8340 8676
rect 15120 8732 15184 8736
rect 15120 8676 15124 8732
rect 15124 8676 15180 8732
rect 15180 8676 15184 8732
rect 15120 8672 15184 8676
rect 15200 8732 15264 8736
rect 15200 8676 15204 8732
rect 15204 8676 15260 8732
rect 15260 8676 15264 8732
rect 15200 8672 15264 8676
rect 15280 8732 15344 8736
rect 15280 8676 15284 8732
rect 15284 8676 15340 8732
rect 15340 8676 15344 8732
rect 15280 8672 15344 8676
rect 15360 8732 15424 8736
rect 15360 8676 15364 8732
rect 15364 8676 15420 8732
rect 15420 8676 15424 8732
rect 15360 8672 15424 8676
rect 22204 8732 22268 8736
rect 22204 8676 22208 8732
rect 22208 8676 22264 8732
rect 22264 8676 22268 8732
rect 22204 8672 22268 8676
rect 22284 8732 22348 8736
rect 22284 8676 22288 8732
rect 22288 8676 22344 8732
rect 22344 8676 22348 8732
rect 22284 8672 22348 8676
rect 22364 8732 22428 8736
rect 22364 8676 22368 8732
rect 22368 8676 22424 8732
rect 22424 8676 22428 8732
rect 22364 8672 22428 8676
rect 22444 8732 22508 8736
rect 22444 8676 22448 8732
rect 22448 8676 22504 8732
rect 22504 8676 22508 8732
rect 22444 8672 22508 8676
rect 29288 8732 29352 8736
rect 29288 8676 29292 8732
rect 29292 8676 29348 8732
rect 29348 8676 29352 8732
rect 29288 8672 29352 8676
rect 29368 8732 29432 8736
rect 29368 8676 29372 8732
rect 29372 8676 29428 8732
rect 29428 8676 29432 8732
rect 29368 8672 29432 8676
rect 29448 8732 29512 8736
rect 29448 8676 29452 8732
rect 29452 8676 29508 8732
rect 29508 8676 29512 8732
rect 29448 8672 29512 8676
rect 29528 8732 29592 8736
rect 29528 8676 29532 8732
rect 29532 8676 29588 8732
rect 29588 8676 29592 8732
rect 29528 8672 29592 8676
rect 4494 8188 4558 8192
rect 4494 8132 4498 8188
rect 4498 8132 4554 8188
rect 4554 8132 4558 8188
rect 4494 8128 4558 8132
rect 4574 8188 4638 8192
rect 4574 8132 4578 8188
rect 4578 8132 4634 8188
rect 4634 8132 4638 8188
rect 4574 8128 4638 8132
rect 4654 8188 4718 8192
rect 4654 8132 4658 8188
rect 4658 8132 4714 8188
rect 4714 8132 4718 8188
rect 4654 8128 4718 8132
rect 4734 8188 4798 8192
rect 4734 8132 4738 8188
rect 4738 8132 4794 8188
rect 4794 8132 4798 8188
rect 4734 8128 4798 8132
rect 11578 8188 11642 8192
rect 11578 8132 11582 8188
rect 11582 8132 11638 8188
rect 11638 8132 11642 8188
rect 11578 8128 11642 8132
rect 11658 8188 11722 8192
rect 11658 8132 11662 8188
rect 11662 8132 11718 8188
rect 11718 8132 11722 8188
rect 11658 8128 11722 8132
rect 11738 8188 11802 8192
rect 11738 8132 11742 8188
rect 11742 8132 11798 8188
rect 11798 8132 11802 8188
rect 11738 8128 11802 8132
rect 11818 8188 11882 8192
rect 11818 8132 11822 8188
rect 11822 8132 11878 8188
rect 11878 8132 11882 8188
rect 11818 8128 11882 8132
rect 18662 8188 18726 8192
rect 18662 8132 18666 8188
rect 18666 8132 18722 8188
rect 18722 8132 18726 8188
rect 18662 8128 18726 8132
rect 18742 8188 18806 8192
rect 18742 8132 18746 8188
rect 18746 8132 18802 8188
rect 18802 8132 18806 8188
rect 18742 8128 18806 8132
rect 18822 8188 18886 8192
rect 18822 8132 18826 8188
rect 18826 8132 18882 8188
rect 18882 8132 18886 8188
rect 18822 8128 18886 8132
rect 18902 8188 18966 8192
rect 18902 8132 18906 8188
rect 18906 8132 18962 8188
rect 18962 8132 18966 8188
rect 18902 8128 18966 8132
rect 25746 8188 25810 8192
rect 25746 8132 25750 8188
rect 25750 8132 25806 8188
rect 25806 8132 25810 8188
rect 25746 8128 25810 8132
rect 25826 8188 25890 8192
rect 25826 8132 25830 8188
rect 25830 8132 25886 8188
rect 25886 8132 25890 8188
rect 25826 8128 25890 8132
rect 25906 8188 25970 8192
rect 25906 8132 25910 8188
rect 25910 8132 25966 8188
rect 25966 8132 25970 8188
rect 25906 8128 25970 8132
rect 25986 8188 26050 8192
rect 25986 8132 25990 8188
rect 25990 8132 26046 8188
rect 26046 8132 26050 8188
rect 25986 8128 26050 8132
rect 22692 7788 22756 7852
rect 8036 7644 8100 7648
rect 8036 7588 8040 7644
rect 8040 7588 8096 7644
rect 8096 7588 8100 7644
rect 8036 7584 8100 7588
rect 8116 7644 8180 7648
rect 8116 7588 8120 7644
rect 8120 7588 8176 7644
rect 8176 7588 8180 7644
rect 8116 7584 8180 7588
rect 8196 7644 8260 7648
rect 8196 7588 8200 7644
rect 8200 7588 8256 7644
rect 8256 7588 8260 7644
rect 8196 7584 8260 7588
rect 8276 7644 8340 7648
rect 8276 7588 8280 7644
rect 8280 7588 8336 7644
rect 8336 7588 8340 7644
rect 8276 7584 8340 7588
rect 15120 7644 15184 7648
rect 15120 7588 15124 7644
rect 15124 7588 15180 7644
rect 15180 7588 15184 7644
rect 15120 7584 15184 7588
rect 15200 7644 15264 7648
rect 15200 7588 15204 7644
rect 15204 7588 15260 7644
rect 15260 7588 15264 7644
rect 15200 7584 15264 7588
rect 15280 7644 15344 7648
rect 15280 7588 15284 7644
rect 15284 7588 15340 7644
rect 15340 7588 15344 7644
rect 15280 7584 15344 7588
rect 15360 7644 15424 7648
rect 15360 7588 15364 7644
rect 15364 7588 15420 7644
rect 15420 7588 15424 7644
rect 15360 7584 15424 7588
rect 22204 7644 22268 7648
rect 22204 7588 22208 7644
rect 22208 7588 22264 7644
rect 22264 7588 22268 7644
rect 22204 7584 22268 7588
rect 22284 7644 22348 7648
rect 22284 7588 22288 7644
rect 22288 7588 22344 7644
rect 22344 7588 22348 7644
rect 22284 7584 22348 7588
rect 22364 7644 22428 7648
rect 22364 7588 22368 7644
rect 22368 7588 22424 7644
rect 22424 7588 22428 7644
rect 22364 7584 22428 7588
rect 22444 7644 22508 7648
rect 22444 7588 22448 7644
rect 22448 7588 22504 7644
rect 22504 7588 22508 7644
rect 22444 7584 22508 7588
rect 29288 7644 29352 7648
rect 29288 7588 29292 7644
rect 29292 7588 29348 7644
rect 29348 7588 29352 7644
rect 29288 7584 29352 7588
rect 29368 7644 29432 7648
rect 29368 7588 29372 7644
rect 29372 7588 29428 7644
rect 29428 7588 29432 7644
rect 29368 7584 29432 7588
rect 29448 7644 29512 7648
rect 29448 7588 29452 7644
rect 29452 7588 29508 7644
rect 29508 7588 29512 7644
rect 29448 7584 29512 7588
rect 29528 7644 29592 7648
rect 29528 7588 29532 7644
rect 29532 7588 29588 7644
rect 29588 7588 29592 7644
rect 29528 7584 29592 7588
rect 4494 7100 4558 7104
rect 4494 7044 4498 7100
rect 4498 7044 4554 7100
rect 4554 7044 4558 7100
rect 4494 7040 4558 7044
rect 4574 7100 4638 7104
rect 4574 7044 4578 7100
rect 4578 7044 4634 7100
rect 4634 7044 4638 7100
rect 4574 7040 4638 7044
rect 4654 7100 4718 7104
rect 4654 7044 4658 7100
rect 4658 7044 4714 7100
rect 4714 7044 4718 7100
rect 4654 7040 4718 7044
rect 4734 7100 4798 7104
rect 4734 7044 4738 7100
rect 4738 7044 4794 7100
rect 4794 7044 4798 7100
rect 4734 7040 4798 7044
rect 11578 7100 11642 7104
rect 11578 7044 11582 7100
rect 11582 7044 11638 7100
rect 11638 7044 11642 7100
rect 11578 7040 11642 7044
rect 11658 7100 11722 7104
rect 11658 7044 11662 7100
rect 11662 7044 11718 7100
rect 11718 7044 11722 7100
rect 11658 7040 11722 7044
rect 11738 7100 11802 7104
rect 11738 7044 11742 7100
rect 11742 7044 11798 7100
rect 11798 7044 11802 7100
rect 11738 7040 11802 7044
rect 11818 7100 11882 7104
rect 11818 7044 11822 7100
rect 11822 7044 11878 7100
rect 11878 7044 11882 7100
rect 11818 7040 11882 7044
rect 18662 7100 18726 7104
rect 18662 7044 18666 7100
rect 18666 7044 18722 7100
rect 18722 7044 18726 7100
rect 18662 7040 18726 7044
rect 18742 7100 18806 7104
rect 18742 7044 18746 7100
rect 18746 7044 18802 7100
rect 18802 7044 18806 7100
rect 18742 7040 18806 7044
rect 18822 7100 18886 7104
rect 18822 7044 18826 7100
rect 18826 7044 18882 7100
rect 18882 7044 18886 7100
rect 18822 7040 18886 7044
rect 18902 7100 18966 7104
rect 18902 7044 18906 7100
rect 18906 7044 18962 7100
rect 18962 7044 18966 7100
rect 18902 7040 18966 7044
rect 25746 7100 25810 7104
rect 25746 7044 25750 7100
rect 25750 7044 25806 7100
rect 25806 7044 25810 7100
rect 25746 7040 25810 7044
rect 25826 7100 25890 7104
rect 25826 7044 25830 7100
rect 25830 7044 25886 7100
rect 25886 7044 25890 7100
rect 25826 7040 25890 7044
rect 25906 7100 25970 7104
rect 25906 7044 25910 7100
rect 25910 7044 25966 7100
rect 25966 7044 25970 7100
rect 25906 7040 25970 7044
rect 25986 7100 26050 7104
rect 25986 7044 25990 7100
rect 25990 7044 26046 7100
rect 26046 7044 26050 7100
rect 25986 7040 26050 7044
rect 8036 6556 8100 6560
rect 8036 6500 8040 6556
rect 8040 6500 8096 6556
rect 8096 6500 8100 6556
rect 8036 6496 8100 6500
rect 8116 6556 8180 6560
rect 8116 6500 8120 6556
rect 8120 6500 8176 6556
rect 8176 6500 8180 6556
rect 8116 6496 8180 6500
rect 8196 6556 8260 6560
rect 8196 6500 8200 6556
rect 8200 6500 8256 6556
rect 8256 6500 8260 6556
rect 8196 6496 8260 6500
rect 8276 6556 8340 6560
rect 8276 6500 8280 6556
rect 8280 6500 8336 6556
rect 8336 6500 8340 6556
rect 8276 6496 8340 6500
rect 15120 6556 15184 6560
rect 15120 6500 15124 6556
rect 15124 6500 15180 6556
rect 15180 6500 15184 6556
rect 15120 6496 15184 6500
rect 15200 6556 15264 6560
rect 15200 6500 15204 6556
rect 15204 6500 15260 6556
rect 15260 6500 15264 6556
rect 15200 6496 15264 6500
rect 15280 6556 15344 6560
rect 15280 6500 15284 6556
rect 15284 6500 15340 6556
rect 15340 6500 15344 6556
rect 15280 6496 15344 6500
rect 15360 6556 15424 6560
rect 15360 6500 15364 6556
rect 15364 6500 15420 6556
rect 15420 6500 15424 6556
rect 15360 6496 15424 6500
rect 22204 6556 22268 6560
rect 22204 6500 22208 6556
rect 22208 6500 22264 6556
rect 22264 6500 22268 6556
rect 22204 6496 22268 6500
rect 22284 6556 22348 6560
rect 22284 6500 22288 6556
rect 22288 6500 22344 6556
rect 22344 6500 22348 6556
rect 22284 6496 22348 6500
rect 22364 6556 22428 6560
rect 22364 6500 22368 6556
rect 22368 6500 22424 6556
rect 22424 6500 22428 6556
rect 22364 6496 22428 6500
rect 22444 6556 22508 6560
rect 22444 6500 22448 6556
rect 22448 6500 22504 6556
rect 22504 6500 22508 6556
rect 22444 6496 22508 6500
rect 29288 6556 29352 6560
rect 29288 6500 29292 6556
rect 29292 6500 29348 6556
rect 29348 6500 29352 6556
rect 29288 6496 29352 6500
rect 29368 6556 29432 6560
rect 29368 6500 29372 6556
rect 29372 6500 29428 6556
rect 29428 6500 29432 6556
rect 29368 6496 29432 6500
rect 29448 6556 29512 6560
rect 29448 6500 29452 6556
rect 29452 6500 29508 6556
rect 29508 6500 29512 6556
rect 29448 6496 29512 6500
rect 29528 6556 29592 6560
rect 29528 6500 29532 6556
rect 29532 6500 29588 6556
rect 29588 6500 29592 6556
rect 29528 6496 29592 6500
rect 4494 6012 4558 6016
rect 4494 5956 4498 6012
rect 4498 5956 4554 6012
rect 4554 5956 4558 6012
rect 4494 5952 4558 5956
rect 4574 6012 4638 6016
rect 4574 5956 4578 6012
rect 4578 5956 4634 6012
rect 4634 5956 4638 6012
rect 4574 5952 4638 5956
rect 4654 6012 4718 6016
rect 4654 5956 4658 6012
rect 4658 5956 4714 6012
rect 4714 5956 4718 6012
rect 4654 5952 4718 5956
rect 4734 6012 4798 6016
rect 4734 5956 4738 6012
rect 4738 5956 4794 6012
rect 4794 5956 4798 6012
rect 4734 5952 4798 5956
rect 11578 6012 11642 6016
rect 11578 5956 11582 6012
rect 11582 5956 11638 6012
rect 11638 5956 11642 6012
rect 11578 5952 11642 5956
rect 11658 6012 11722 6016
rect 11658 5956 11662 6012
rect 11662 5956 11718 6012
rect 11718 5956 11722 6012
rect 11658 5952 11722 5956
rect 11738 6012 11802 6016
rect 11738 5956 11742 6012
rect 11742 5956 11798 6012
rect 11798 5956 11802 6012
rect 11738 5952 11802 5956
rect 11818 6012 11882 6016
rect 11818 5956 11822 6012
rect 11822 5956 11878 6012
rect 11878 5956 11882 6012
rect 11818 5952 11882 5956
rect 18662 6012 18726 6016
rect 18662 5956 18666 6012
rect 18666 5956 18722 6012
rect 18722 5956 18726 6012
rect 18662 5952 18726 5956
rect 18742 6012 18806 6016
rect 18742 5956 18746 6012
rect 18746 5956 18802 6012
rect 18802 5956 18806 6012
rect 18742 5952 18806 5956
rect 18822 6012 18886 6016
rect 18822 5956 18826 6012
rect 18826 5956 18882 6012
rect 18882 5956 18886 6012
rect 18822 5952 18886 5956
rect 18902 6012 18966 6016
rect 18902 5956 18906 6012
rect 18906 5956 18962 6012
rect 18962 5956 18966 6012
rect 18902 5952 18966 5956
rect 25746 6012 25810 6016
rect 25746 5956 25750 6012
rect 25750 5956 25806 6012
rect 25806 5956 25810 6012
rect 25746 5952 25810 5956
rect 25826 6012 25890 6016
rect 25826 5956 25830 6012
rect 25830 5956 25886 6012
rect 25886 5956 25890 6012
rect 25826 5952 25890 5956
rect 25906 6012 25970 6016
rect 25906 5956 25910 6012
rect 25910 5956 25966 6012
rect 25966 5956 25970 6012
rect 25906 5952 25970 5956
rect 25986 6012 26050 6016
rect 25986 5956 25990 6012
rect 25990 5956 26046 6012
rect 26046 5956 26050 6012
rect 25986 5952 26050 5956
rect 8036 5468 8100 5472
rect 8036 5412 8040 5468
rect 8040 5412 8096 5468
rect 8096 5412 8100 5468
rect 8036 5408 8100 5412
rect 8116 5468 8180 5472
rect 8116 5412 8120 5468
rect 8120 5412 8176 5468
rect 8176 5412 8180 5468
rect 8116 5408 8180 5412
rect 8196 5468 8260 5472
rect 8196 5412 8200 5468
rect 8200 5412 8256 5468
rect 8256 5412 8260 5468
rect 8196 5408 8260 5412
rect 8276 5468 8340 5472
rect 8276 5412 8280 5468
rect 8280 5412 8336 5468
rect 8336 5412 8340 5468
rect 8276 5408 8340 5412
rect 15120 5468 15184 5472
rect 15120 5412 15124 5468
rect 15124 5412 15180 5468
rect 15180 5412 15184 5468
rect 15120 5408 15184 5412
rect 15200 5468 15264 5472
rect 15200 5412 15204 5468
rect 15204 5412 15260 5468
rect 15260 5412 15264 5468
rect 15200 5408 15264 5412
rect 15280 5468 15344 5472
rect 15280 5412 15284 5468
rect 15284 5412 15340 5468
rect 15340 5412 15344 5468
rect 15280 5408 15344 5412
rect 15360 5468 15424 5472
rect 15360 5412 15364 5468
rect 15364 5412 15420 5468
rect 15420 5412 15424 5468
rect 15360 5408 15424 5412
rect 22204 5468 22268 5472
rect 22204 5412 22208 5468
rect 22208 5412 22264 5468
rect 22264 5412 22268 5468
rect 22204 5408 22268 5412
rect 22284 5468 22348 5472
rect 22284 5412 22288 5468
rect 22288 5412 22344 5468
rect 22344 5412 22348 5468
rect 22284 5408 22348 5412
rect 22364 5468 22428 5472
rect 22364 5412 22368 5468
rect 22368 5412 22424 5468
rect 22424 5412 22428 5468
rect 22364 5408 22428 5412
rect 22444 5468 22508 5472
rect 22444 5412 22448 5468
rect 22448 5412 22504 5468
rect 22504 5412 22508 5468
rect 22444 5408 22508 5412
rect 29288 5468 29352 5472
rect 29288 5412 29292 5468
rect 29292 5412 29348 5468
rect 29348 5412 29352 5468
rect 29288 5408 29352 5412
rect 29368 5468 29432 5472
rect 29368 5412 29372 5468
rect 29372 5412 29428 5468
rect 29428 5412 29432 5468
rect 29368 5408 29432 5412
rect 29448 5468 29512 5472
rect 29448 5412 29452 5468
rect 29452 5412 29508 5468
rect 29508 5412 29512 5468
rect 29448 5408 29512 5412
rect 29528 5468 29592 5472
rect 29528 5412 29532 5468
rect 29532 5412 29588 5468
rect 29588 5412 29592 5468
rect 29528 5408 29592 5412
rect 27844 5068 27908 5132
rect 4494 4924 4558 4928
rect 4494 4868 4498 4924
rect 4498 4868 4554 4924
rect 4554 4868 4558 4924
rect 4494 4864 4558 4868
rect 4574 4924 4638 4928
rect 4574 4868 4578 4924
rect 4578 4868 4634 4924
rect 4634 4868 4638 4924
rect 4574 4864 4638 4868
rect 4654 4924 4718 4928
rect 4654 4868 4658 4924
rect 4658 4868 4714 4924
rect 4714 4868 4718 4924
rect 4654 4864 4718 4868
rect 4734 4924 4798 4928
rect 4734 4868 4738 4924
rect 4738 4868 4794 4924
rect 4794 4868 4798 4924
rect 4734 4864 4798 4868
rect 11578 4924 11642 4928
rect 11578 4868 11582 4924
rect 11582 4868 11638 4924
rect 11638 4868 11642 4924
rect 11578 4864 11642 4868
rect 11658 4924 11722 4928
rect 11658 4868 11662 4924
rect 11662 4868 11718 4924
rect 11718 4868 11722 4924
rect 11658 4864 11722 4868
rect 11738 4924 11802 4928
rect 11738 4868 11742 4924
rect 11742 4868 11798 4924
rect 11798 4868 11802 4924
rect 11738 4864 11802 4868
rect 11818 4924 11882 4928
rect 11818 4868 11822 4924
rect 11822 4868 11878 4924
rect 11878 4868 11882 4924
rect 11818 4864 11882 4868
rect 18662 4924 18726 4928
rect 18662 4868 18666 4924
rect 18666 4868 18722 4924
rect 18722 4868 18726 4924
rect 18662 4864 18726 4868
rect 18742 4924 18806 4928
rect 18742 4868 18746 4924
rect 18746 4868 18802 4924
rect 18802 4868 18806 4924
rect 18742 4864 18806 4868
rect 18822 4924 18886 4928
rect 18822 4868 18826 4924
rect 18826 4868 18882 4924
rect 18882 4868 18886 4924
rect 18822 4864 18886 4868
rect 18902 4924 18966 4928
rect 18902 4868 18906 4924
rect 18906 4868 18962 4924
rect 18962 4868 18966 4924
rect 18902 4864 18966 4868
rect 25746 4924 25810 4928
rect 25746 4868 25750 4924
rect 25750 4868 25806 4924
rect 25806 4868 25810 4924
rect 25746 4864 25810 4868
rect 25826 4924 25890 4928
rect 25826 4868 25830 4924
rect 25830 4868 25886 4924
rect 25886 4868 25890 4924
rect 25826 4864 25890 4868
rect 25906 4924 25970 4928
rect 25906 4868 25910 4924
rect 25910 4868 25966 4924
rect 25966 4868 25970 4924
rect 25906 4864 25970 4868
rect 25986 4924 26050 4928
rect 25986 4868 25990 4924
rect 25990 4868 26046 4924
rect 26046 4868 26050 4924
rect 25986 4864 26050 4868
rect 8036 4380 8100 4384
rect 8036 4324 8040 4380
rect 8040 4324 8096 4380
rect 8096 4324 8100 4380
rect 8036 4320 8100 4324
rect 8116 4380 8180 4384
rect 8116 4324 8120 4380
rect 8120 4324 8176 4380
rect 8176 4324 8180 4380
rect 8116 4320 8180 4324
rect 8196 4380 8260 4384
rect 8196 4324 8200 4380
rect 8200 4324 8256 4380
rect 8256 4324 8260 4380
rect 8196 4320 8260 4324
rect 8276 4380 8340 4384
rect 8276 4324 8280 4380
rect 8280 4324 8336 4380
rect 8336 4324 8340 4380
rect 8276 4320 8340 4324
rect 15120 4380 15184 4384
rect 15120 4324 15124 4380
rect 15124 4324 15180 4380
rect 15180 4324 15184 4380
rect 15120 4320 15184 4324
rect 15200 4380 15264 4384
rect 15200 4324 15204 4380
rect 15204 4324 15260 4380
rect 15260 4324 15264 4380
rect 15200 4320 15264 4324
rect 15280 4380 15344 4384
rect 15280 4324 15284 4380
rect 15284 4324 15340 4380
rect 15340 4324 15344 4380
rect 15280 4320 15344 4324
rect 15360 4380 15424 4384
rect 15360 4324 15364 4380
rect 15364 4324 15420 4380
rect 15420 4324 15424 4380
rect 15360 4320 15424 4324
rect 22204 4380 22268 4384
rect 22204 4324 22208 4380
rect 22208 4324 22264 4380
rect 22264 4324 22268 4380
rect 22204 4320 22268 4324
rect 22284 4380 22348 4384
rect 22284 4324 22288 4380
rect 22288 4324 22344 4380
rect 22344 4324 22348 4380
rect 22284 4320 22348 4324
rect 22364 4380 22428 4384
rect 22364 4324 22368 4380
rect 22368 4324 22424 4380
rect 22424 4324 22428 4380
rect 22364 4320 22428 4324
rect 22444 4380 22508 4384
rect 22444 4324 22448 4380
rect 22448 4324 22504 4380
rect 22504 4324 22508 4380
rect 22444 4320 22508 4324
rect 29288 4380 29352 4384
rect 29288 4324 29292 4380
rect 29292 4324 29348 4380
rect 29348 4324 29352 4380
rect 29288 4320 29352 4324
rect 29368 4380 29432 4384
rect 29368 4324 29372 4380
rect 29372 4324 29428 4380
rect 29428 4324 29432 4380
rect 29368 4320 29432 4324
rect 29448 4380 29512 4384
rect 29448 4324 29452 4380
rect 29452 4324 29508 4380
rect 29508 4324 29512 4380
rect 29448 4320 29512 4324
rect 29528 4380 29592 4384
rect 29528 4324 29532 4380
rect 29532 4324 29588 4380
rect 29588 4324 29592 4380
rect 29528 4320 29592 4324
rect 4494 3836 4558 3840
rect 4494 3780 4498 3836
rect 4498 3780 4554 3836
rect 4554 3780 4558 3836
rect 4494 3776 4558 3780
rect 4574 3836 4638 3840
rect 4574 3780 4578 3836
rect 4578 3780 4634 3836
rect 4634 3780 4638 3836
rect 4574 3776 4638 3780
rect 4654 3836 4718 3840
rect 4654 3780 4658 3836
rect 4658 3780 4714 3836
rect 4714 3780 4718 3836
rect 4654 3776 4718 3780
rect 4734 3836 4798 3840
rect 4734 3780 4738 3836
rect 4738 3780 4794 3836
rect 4794 3780 4798 3836
rect 4734 3776 4798 3780
rect 11578 3836 11642 3840
rect 11578 3780 11582 3836
rect 11582 3780 11638 3836
rect 11638 3780 11642 3836
rect 11578 3776 11642 3780
rect 11658 3836 11722 3840
rect 11658 3780 11662 3836
rect 11662 3780 11718 3836
rect 11718 3780 11722 3836
rect 11658 3776 11722 3780
rect 11738 3836 11802 3840
rect 11738 3780 11742 3836
rect 11742 3780 11798 3836
rect 11798 3780 11802 3836
rect 11738 3776 11802 3780
rect 11818 3836 11882 3840
rect 11818 3780 11822 3836
rect 11822 3780 11878 3836
rect 11878 3780 11882 3836
rect 11818 3776 11882 3780
rect 18662 3836 18726 3840
rect 18662 3780 18666 3836
rect 18666 3780 18722 3836
rect 18722 3780 18726 3836
rect 18662 3776 18726 3780
rect 18742 3836 18806 3840
rect 18742 3780 18746 3836
rect 18746 3780 18802 3836
rect 18802 3780 18806 3836
rect 18742 3776 18806 3780
rect 18822 3836 18886 3840
rect 18822 3780 18826 3836
rect 18826 3780 18882 3836
rect 18882 3780 18886 3836
rect 18822 3776 18886 3780
rect 18902 3836 18966 3840
rect 18902 3780 18906 3836
rect 18906 3780 18962 3836
rect 18962 3780 18966 3836
rect 18902 3776 18966 3780
rect 25746 3836 25810 3840
rect 25746 3780 25750 3836
rect 25750 3780 25806 3836
rect 25806 3780 25810 3836
rect 25746 3776 25810 3780
rect 25826 3836 25890 3840
rect 25826 3780 25830 3836
rect 25830 3780 25886 3836
rect 25886 3780 25890 3836
rect 25826 3776 25890 3780
rect 25906 3836 25970 3840
rect 25906 3780 25910 3836
rect 25910 3780 25966 3836
rect 25966 3780 25970 3836
rect 25906 3776 25970 3780
rect 25986 3836 26050 3840
rect 25986 3780 25990 3836
rect 25990 3780 26046 3836
rect 26046 3780 26050 3836
rect 25986 3776 26050 3780
rect 8036 3292 8100 3296
rect 8036 3236 8040 3292
rect 8040 3236 8096 3292
rect 8096 3236 8100 3292
rect 8036 3232 8100 3236
rect 8116 3292 8180 3296
rect 8116 3236 8120 3292
rect 8120 3236 8176 3292
rect 8176 3236 8180 3292
rect 8116 3232 8180 3236
rect 8196 3292 8260 3296
rect 8196 3236 8200 3292
rect 8200 3236 8256 3292
rect 8256 3236 8260 3292
rect 8196 3232 8260 3236
rect 8276 3292 8340 3296
rect 8276 3236 8280 3292
rect 8280 3236 8336 3292
rect 8336 3236 8340 3292
rect 8276 3232 8340 3236
rect 15120 3292 15184 3296
rect 15120 3236 15124 3292
rect 15124 3236 15180 3292
rect 15180 3236 15184 3292
rect 15120 3232 15184 3236
rect 15200 3292 15264 3296
rect 15200 3236 15204 3292
rect 15204 3236 15260 3292
rect 15260 3236 15264 3292
rect 15200 3232 15264 3236
rect 15280 3292 15344 3296
rect 15280 3236 15284 3292
rect 15284 3236 15340 3292
rect 15340 3236 15344 3292
rect 15280 3232 15344 3236
rect 15360 3292 15424 3296
rect 15360 3236 15364 3292
rect 15364 3236 15420 3292
rect 15420 3236 15424 3292
rect 15360 3232 15424 3236
rect 22204 3292 22268 3296
rect 22204 3236 22208 3292
rect 22208 3236 22264 3292
rect 22264 3236 22268 3292
rect 22204 3232 22268 3236
rect 22284 3292 22348 3296
rect 22284 3236 22288 3292
rect 22288 3236 22344 3292
rect 22344 3236 22348 3292
rect 22284 3232 22348 3236
rect 22364 3292 22428 3296
rect 22364 3236 22368 3292
rect 22368 3236 22424 3292
rect 22424 3236 22428 3292
rect 22364 3232 22428 3236
rect 22444 3292 22508 3296
rect 22444 3236 22448 3292
rect 22448 3236 22504 3292
rect 22504 3236 22508 3292
rect 22444 3232 22508 3236
rect 29288 3292 29352 3296
rect 29288 3236 29292 3292
rect 29292 3236 29348 3292
rect 29348 3236 29352 3292
rect 29288 3232 29352 3236
rect 29368 3292 29432 3296
rect 29368 3236 29372 3292
rect 29372 3236 29428 3292
rect 29428 3236 29432 3292
rect 29368 3232 29432 3236
rect 29448 3292 29512 3296
rect 29448 3236 29452 3292
rect 29452 3236 29508 3292
rect 29508 3236 29512 3292
rect 29448 3232 29512 3236
rect 29528 3292 29592 3296
rect 29528 3236 29532 3292
rect 29532 3236 29588 3292
rect 29588 3236 29592 3292
rect 29528 3232 29592 3236
rect 4494 2748 4558 2752
rect 4494 2692 4498 2748
rect 4498 2692 4554 2748
rect 4554 2692 4558 2748
rect 4494 2688 4558 2692
rect 4574 2748 4638 2752
rect 4574 2692 4578 2748
rect 4578 2692 4634 2748
rect 4634 2692 4638 2748
rect 4574 2688 4638 2692
rect 4654 2748 4718 2752
rect 4654 2692 4658 2748
rect 4658 2692 4714 2748
rect 4714 2692 4718 2748
rect 4654 2688 4718 2692
rect 4734 2748 4798 2752
rect 4734 2692 4738 2748
rect 4738 2692 4794 2748
rect 4794 2692 4798 2748
rect 4734 2688 4798 2692
rect 11578 2748 11642 2752
rect 11578 2692 11582 2748
rect 11582 2692 11638 2748
rect 11638 2692 11642 2748
rect 11578 2688 11642 2692
rect 11658 2748 11722 2752
rect 11658 2692 11662 2748
rect 11662 2692 11718 2748
rect 11718 2692 11722 2748
rect 11658 2688 11722 2692
rect 11738 2748 11802 2752
rect 11738 2692 11742 2748
rect 11742 2692 11798 2748
rect 11798 2692 11802 2748
rect 11738 2688 11802 2692
rect 11818 2748 11882 2752
rect 11818 2692 11822 2748
rect 11822 2692 11878 2748
rect 11878 2692 11882 2748
rect 11818 2688 11882 2692
rect 18662 2748 18726 2752
rect 18662 2692 18666 2748
rect 18666 2692 18722 2748
rect 18722 2692 18726 2748
rect 18662 2688 18726 2692
rect 18742 2748 18806 2752
rect 18742 2692 18746 2748
rect 18746 2692 18802 2748
rect 18802 2692 18806 2748
rect 18742 2688 18806 2692
rect 18822 2748 18886 2752
rect 18822 2692 18826 2748
rect 18826 2692 18882 2748
rect 18882 2692 18886 2748
rect 18822 2688 18886 2692
rect 18902 2748 18966 2752
rect 18902 2692 18906 2748
rect 18906 2692 18962 2748
rect 18962 2692 18966 2748
rect 18902 2688 18966 2692
rect 25746 2748 25810 2752
rect 25746 2692 25750 2748
rect 25750 2692 25806 2748
rect 25806 2692 25810 2748
rect 25746 2688 25810 2692
rect 25826 2748 25890 2752
rect 25826 2692 25830 2748
rect 25830 2692 25886 2748
rect 25886 2692 25890 2748
rect 25826 2688 25890 2692
rect 25906 2748 25970 2752
rect 25906 2692 25910 2748
rect 25910 2692 25966 2748
rect 25966 2692 25970 2748
rect 25906 2688 25970 2692
rect 25986 2748 26050 2752
rect 25986 2692 25990 2748
rect 25990 2692 26046 2748
rect 26046 2692 26050 2748
rect 25986 2688 26050 2692
rect 8036 2204 8100 2208
rect 8036 2148 8040 2204
rect 8040 2148 8096 2204
rect 8096 2148 8100 2204
rect 8036 2144 8100 2148
rect 8116 2204 8180 2208
rect 8116 2148 8120 2204
rect 8120 2148 8176 2204
rect 8176 2148 8180 2204
rect 8116 2144 8180 2148
rect 8196 2204 8260 2208
rect 8196 2148 8200 2204
rect 8200 2148 8256 2204
rect 8256 2148 8260 2204
rect 8196 2144 8260 2148
rect 8276 2204 8340 2208
rect 8276 2148 8280 2204
rect 8280 2148 8336 2204
rect 8336 2148 8340 2204
rect 8276 2144 8340 2148
rect 15120 2204 15184 2208
rect 15120 2148 15124 2204
rect 15124 2148 15180 2204
rect 15180 2148 15184 2204
rect 15120 2144 15184 2148
rect 15200 2204 15264 2208
rect 15200 2148 15204 2204
rect 15204 2148 15260 2204
rect 15260 2148 15264 2204
rect 15200 2144 15264 2148
rect 15280 2204 15344 2208
rect 15280 2148 15284 2204
rect 15284 2148 15340 2204
rect 15340 2148 15344 2204
rect 15280 2144 15344 2148
rect 15360 2204 15424 2208
rect 15360 2148 15364 2204
rect 15364 2148 15420 2204
rect 15420 2148 15424 2204
rect 15360 2144 15424 2148
rect 22204 2204 22268 2208
rect 22204 2148 22208 2204
rect 22208 2148 22264 2204
rect 22264 2148 22268 2204
rect 22204 2144 22268 2148
rect 22284 2204 22348 2208
rect 22284 2148 22288 2204
rect 22288 2148 22344 2204
rect 22344 2148 22348 2204
rect 22284 2144 22348 2148
rect 22364 2204 22428 2208
rect 22364 2148 22368 2204
rect 22368 2148 22424 2204
rect 22424 2148 22428 2204
rect 22364 2144 22428 2148
rect 22444 2204 22508 2208
rect 22444 2148 22448 2204
rect 22448 2148 22504 2204
rect 22504 2148 22508 2204
rect 22444 2144 22508 2148
rect 29288 2204 29352 2208
rect 29288 2148 29292 2204
rect 29292 2148 29348 2204
rect 29348 2148 29352 2204
rect 29288 2144 29352 2148
rect 29368 2204 29432 2208
rect 29368 2148 29372 2204
rect 29372 2148 29428 2204
rect 29428 2148 29432 2204
rect 29368 2144 29432 2148
rect 29448 2204 29512 2208
rect 29448 2148 29452 2204
rect 29452 2148 29508 2204
rect 29508 2148 29512 2204
rect 29448 2144 29512 2148
rect 29528 2204 29592 2208
rect 29528 2148 29532 2204
rect 29532 2148 29588 2204
rect 29588 2148 29592 2204
rect 29528 2144 29592 2148
<< metal4 >>
rect 4486 29952 4806 30512
rect 4486 29888 4494 29952
rect 4558 29888 4574 29952
rect 4638 29888 4654 29952
rect 4718 29888 4734 29952
rect 4798 29888 4806 29952
rect 4486 28864 4806 29888
rect 4486 28800 4494 28864
rect 4558 28800 4574 28864
rect 4638 28800 4654 28864
rect 4718 28800 4734 28864
rect 4798 28800 4806 28864
rect 4486 27776 4806 28800
rect 4486 27712 4494 27776
rect 4558 27712 4574 27776
rect 4638 27712 4654 27776
rect 4718 27712 4734 27776
rect 4798 27712 4806 27776
rect 4486 26688 4806 27712
rect 4486 26624 4494 26688
rect 4558 26624 4574 26688
rect 4638 26624 4654 26688
rect 4718 26624 4734 26688
rect 4798 26624 4806 26688
rect 4486 25600 4806 26624
rect 4486 25536 4494 25600
rect 4558 25536 4574 25600
rect 4638 25536 4654 25600
rect 4718 25536 4734 25600
rect 4798 25536 4806 25600
rect 4486 24512 4806 25536
rect 4486 24448 4494 24512
rect 4558 24448 4574 24512
rect 4638 24448 4654 24512
rect 4718 24448 4734 24512
rect 4798 24448 4806 24512
rect 4486 23424 4806 24448
rect 4486 23360 4494 23424
rect 4558 23360 4574 23424
rect 4638 23360 4654 23424
rect 4718 23360 4734 23424
rect 4798 23360 4806 23424
rect 4486 22336 4806 23360
rect 4486 22272 4494 22336
rect 4558 22272 4574 22336
rect 4638 22272 4654 22336
rect 4718 22272 4734 22336
rect 4798 22272 4806 22336
rect 4486 21248 4806 22272
rect 4486 21184 4494 21248
rect 4558 21184 4574 21248
rect 4638 21184 4654 21248
rect 4718 21184 4734 21248
rect 4798 21184 4806 21248
rect 4486 20160 4806 21184
rect 4486 20096 4494 20160
rect 4558 20096 4574 20160
rect 4638 20096 4654 20160
rect 4718 20096 4734 20160
rect 4798 20096 4806 20160
rect 4486 19072 4806 20096
rect 4486 19008 4494 19072
rect 4558 19008 4574 19072
rect 4638 19008 4654 19072
rect 4718 19008 4734 19072
rect 4798 19008 4806 19072
rect 4486 17984 4806 19008
rect 4486 17920 4494 17984
rect 4558 17920 4574 17984
rect 4638 17920 4654 17984
rect 4718 17920 4734 17984
rect 4798 17920 4806 17984
rect 4486 16896 4806 17920
rect 4486 16832 4494 16896
rect 4558 16832 4574 16896
rect 4638 16832 4654 16896
rect 4718 16832 4734 16896
rect 4798 16832 4806 16896
rect 4486 15808 4806 16832
rect 4486 15744 4494 15808
rect 4558 15744 4574 15808
rect 4638 15744 4654 15808
rect 4718 15744 4734 15808
rect 4798 15744 4806 15808
rect 4486 14720 4806 15744
rect 4486 14656 4494 14720
rect 4558 14656 4574 14720
rect 4638 14656 4654 14720
rect 4718 14656 4734 14720
rect 4798 14656 4806 14720
rect 4486 13632 4806 14656
rect 4486 13568 4494 13632
rect 4558 13568 4574 13632
rect 4638 13568 4654 13632
rect 4718 13568 4734 13632
rect 4798 13568 4806 13632
rect 4486 12544 4806 13568
rect 4486 12480 4494 12544
rect 4558 12480 4574 12544
rect 4638 12480 4654 12544
rect 4718 12480 4734 12544
rect 4798 12480 4806 12544
rect 4486 11456 4806 12480
rect 4486 11392 4494 11456
rect 4558 11392 4574 11456
rect 4638 11392 4654 11456
rect 4718 11392 4734 11456
rect 4798 11392 4806 11456
rect 4486 10368 4806 11392
rect 4486 10304 4494 10368
rect 4558 10304 4574 10368
rect 4638 10304 4654 10368
rect 4718 10304 4734 10368
rect 4798 10304 4806 10368
rect 4486 9280 4806 10304
rect 4486 9216 4494 9280
rect 4558 9216 4574 9280
rect 4638 9216 4654 9280
rect 4718 9216 4734 9280
rect 4798 9216 4806 9280
rect 4486 8192 4806 9216
rect 4486 8128 4494 8192
rect 4558 8128 4574 8192
rect 4638 8128 4654 8192
rect 4718 8128 4734 8192
rect 4798 8128 4806 8192
rect 4486 7104 4806 8128
rect 4486 7040 4494 7104
rect 4558 7040 4574 7104
rect 4638 7040 4654 7104
rect 4718 7040 4734 7104
rect 4798 7040 4806 7104
rect 4486 6016 4806 7040
rect 4486 5952 4494 6016
rect 4558 5952 4574 6016
rect 4638 5952 4654 6016
rect 4718 5952 4734 6016
rect 4798 5952 4806 6016
rect 4486 4928 4806 5952
rect 4486 4864 4494 4928
rect 4558 4864 4574 4928
rect 4638 4864 4654 4928
rect 4718 4864 4734 4928
rect 4798 4864 4806 4928
rect 4486 3840 4806 4864
rect 4486 3776 4494 3840
rect 4558 3776 4574 3840
rect 4638 3776 4654 3840
rect 4718 3776 4734 3840
rect 4798 3776 4806 3840
rect 4486 2752 4806 3776
rect 4486 2688 4494 2752
rect 4558 2688 4574 2752
rect 4638 2688 4654 2752
rect 4718 2688 4734 2752
rect 4798 2688 4806 2752
rect 4486 2128 4806 2688
rect 8028 30496 8348 30512
rect 8028 30432 8036 30496
rect 8100 30432 8116 30496
rect 8180 30432 8196 30496
rect 8260 30432 8276 30496
rect 8340 30432 8348 30496
rect 8028 29408 8348 30432
rect 8028 29344 8036 29408
rect 8100 29344 8116 29408
rect 8180 29344 8196 29408
rect 8260 29344 8276 29408
rect 8340 29344 8348 29408
rect 8028 28320 8348 29344
rect 8028 28256 8036 28320
rect 8100 28256 8116 28320
rect 8180 28256 8196 28320
rect 8260 28256 8276 28320
rect 8340 28256 8348 28320
rect 8028 27232 8348 28256
rect 8028 27168 8036 27232
rect 8100 27168 8116 27232
rect 8180 27168 8196 27232
rect 8260 27168 8276 27232
rect 8340 27168 8348 27232
rect 8028 26144 8348 27168
rect 8028 26080 8036 26144
rect 8100 26080 8116 26144
rect 8180 26080 8196 26144
rect 8260 26080 8276 26144
rect 8340 26080 8348 26144
rect 8028 25056 8348 26080
rect 8028 24992 8036 25056
rect 8100 24992 8116 25056
rect 8180 24992 8196 25056
rect 8260 24992 8276 25056
rect 8340 24992 8348 25056
rect 8028 23968 8348 24992
rect 8028 23904 8036 23968
rect 8100 23904 8116 23968
rect 8180 23904 8196 23968
rect 8260 23904 8276 23968
rect 8340 23904 8348 23968
rect 8028 22880 8348 23904
rect 8028 22816 8036 22880
rect 8100 22816 8116 22880
rect 8180 22816 8196 22880
rect 8260 22816 8276 22880
rect 8340 22816 8348 22880
rect 8028 21792 8348 22816
rect 8028 21728 8036 21792
rect 8100 21728 8116 21792
rect 8180 21728 8196 21792
rect 8260 21728 8276 21792
rect 8340 21728 8348 21792
rect 8028 20704 8348 21728
rect 8028 20640 8036 20704
rect 8100 20640 8116 20704
rect 8180 20640 8196 20704
rect 8260 20640 8276 20704
rect 8340 20640 8348 20704
rect 8028 19616 8348 20640
rect 8028 19552 8036 19616
rect 8100 19552 8116 19616
rect 8180 19552 8196 19616
rect 8260 19552 8276 19616
rect 8340 19552 8348 19616
rect 8028 18528 8348 19552
rect 8028 18464 8036 18528
rect 8100 18464 8116 18528
rect 8180 18464 8196 18528
rect 8260 18464 8276 18528
rect 8340 18464 8348 18528
rect 8028 17440 8348 18464
rect 8028 17376 8036 17440
rect 8100 17376 8116 17440
rect 8180 17376 8196 17440
rect 8260 17376 8276 17440
rect 8340 17376 8348 17440
rect 8028 16352 8348 17376
rect 8028 16288 8036 16352
rect 8100 16288 8116 16352
rect 8180 16288 8196 16352
rect 8260 16288 8276 16352
rect 8340 16288 8348 16352
rect 8028 15264 8348 16288
rect 8028 15200 8036 15264
rect 8100 15200 8116 15264
rect 8180 15200 8196 15264
rect 8260 15200 8276 15264
rect 8340 15200 8348 15264
rect 8028 14176 8348 15200
rect 8028 14112 8036 14176
rect 8100 14112 8116 14176
rect 8180 14112 8196 14176
rect 8260 14112 8276 14176
rect 8340 14112 8348 14176
rect 8028 13088 8348 14112
rect 8028 13024 8036 13088
rect 8100 13024 8116 13088
rect 8180 13024 8196 13088
rect 8260 13024 8276 13088
rect 8340 13024 8348 13088
rect 8028 12000 8348 13024
rect 8028 11936 8036 12000
rect 8100 11936 8116 12000
rect 8180 11936 8196 12000
rect 8260 11936 8276 12000
rect 8340 11936 8348 12000
rect 8028 10912 8348 11936
rect 8028 10848 8036 10912
rect 8100 10848 8116 10912
rect 8180 10848 8196 10912
rect 8260 10848 8276 10912
rect 8340 10848 8348 10912
rect 8028 9824 8348 10848
rect 8028 9760 8036 9824
rect 8100 9760 8116 9824
rect 8180 9760 8196 9824
rect 8260 9760 8276 9824
rect 8340 9760 8348 9824
rect 8028 8736 8348 9760
rect 8028 8672 8036 8736
rect 8100 8672 8116 8736
rect 8180 8672 8196 8736
rect 8260 8672 8276 8736
rect 8340 8672 8348 8736
rect 8028 7648 8348 8672
rect 8028 7584 8036 7648
rect 8100 7584 8116 7648
rect 8180 7584 8196 7648
rect 8260 7584 8276 7648
rect 8340 7584 8348 7648
rect 8028 6560 8348 7584
rect 8028 6496 8036 6560
rect 8100 6496 8116 6560
rect 8180 6496 8196 6560
rect 8260 6496 8276 6560
rect 8340 6496 8348 6560
rect 8028 5472 8348 6496
rect 8028 5408 8036 5472
rect 8100 5408 8116 5472
rect 8180 5408 8196 5472
rect 8260 5408 8276 5472
rect 8340 5408 8348 5472
rect 8028 4384 8348 5408
rect 8028 4320 8036 4384
rect 8100 4320 8116 4384
rect 8180 4320 8196 4384
rect 8260 4320 8276 4384
rect 8340 4320 8348 4384
rect 8028 3296 8348 4320
rect 8028 3232 8036 3296
rect 8100 3232 8116 3296
rect 8180 3232 8196 3296
rect 8260 3232 8276 3296
rect 8340 3232 8348 3296
rect 8028 2208 8348 3232
rect 8028 2144 8036 2208
rect 8100 2144 8116 2208
rect 8180 2144 8196 2208
rect 8260 2144 8276 2208
rect 8340 2144 8348 2208
rect 8028 2128 8348 2144
rect 11570 29952 11890 30512
rect 11570 29888 11578 29952
rect 11642 29888 11658 29952
rect 11722 29888 11738 29952
rect 11802 29888 11818 29952
rect 11882 29888 11890 29952
rect 11570 28864 11890 29888
rect 11570 28800 11578 28864
rect 11642 28800 11658 28864
rect 11722 28800 11738 28864
rect 11802 28800 11818 28864
rect 11882 28800 11890 28864
rect 11570 27776 11890 28800
rect 11570 27712 11578 27776
rect 11642 27712 11658 27776
rect 11722 27712 11738 27776
rect 11802 27712 11818 27776
rect 11882 27712 11890 27776
rect 11570 26688 11890 27712
rect 11570 26624 11578 26688
rect 11642 26624 11658 26688
rect 11722 26624 11738 26688
rect 11802 26624 11818 26688
rect 11882 26624 11890 26688
rect 11570 25600 11890 26624
rect 11570 25536 11578 25600
rect 11642 25536 11658 25600
rect 11722 25536 11738 25600
rect 11802 25536 11818 25600
rect 11882 25536 11890 25600
rect 11570 24512 11890 25536
rect 11570 24448 11578 24512
rect 11642 24448 11658 24512
rect 11722 24448 11738 24512
rect 11802 24448 11818 24512
rect 11882 24448 11890 24512
rect 11570 23424 11890 24448
rect 11570 23360 11578 23424
rect 11642 23360 11658 23424
rect 11722 23360 11738 23424
rect 11802 23360 11818 23424
rect 11882 23360 11890 23424
rect 11570 22336 11890 23360
rect 11570 22272 11578 22336
rect 11642 22272 11658 22336
rect 11722 22272 11738 22336
rect 11802 22272 11818 22336
rect 11882 22272 11890 22336
rect 11570 21248 11890 22272
rect 11570 21184 11578 21248
rect 11642 21184 11658 21248
rect 11722 21184 11738 21248
rect 11802 21184 11818 21248
rect 11882 21184 11890 21248
rect 11570 20160 11890 21184
rect 11570 20096 11578 20160
rect 11642 20096 11658 20160
rect 11722 20096 11738 20160
rect 11802 20096 11818 20160
rect 11882 20096 11890 20160
rect 11570 19072 11890 20096
rect 11570 19008 11578 19072
rect 11642 19008 11658 19072
rect 11722 19008 11738 19072
rect 11802 19008 11818 19072
rect 11882 19008 11890 19072
rect 11570 17984 11890 19008
rect 11570 17920 11578 17984
rect 11642 17920 11658 17984
rect 11722 17920 11738 17984
rect 11802 17920 11818 17984
rect 11882 17920 11890 17984
rect 11570 16896 11890 17920
rect 11570 16832 11578 16896
rect 11642 16832 11658 16896
rect 11722 16832 11738 16896
rect 11802 16832 11818 16896
rect 11882 16832 11890 16896
rect 11570 15808 11890 16832
rect 11570 15744 11578 15808
rect 11642 15744 11658 15808
rect 11722 15744 11738 15808
rect 11802 15744 11818 15808
rect 11882 15744 11890 15808
rect 11570 14720 11890 15744
rect 11570 14656 11578 14720
rect 11642 14656 11658 14720
rect 11722 14656 11738 14720
rect 11802 14656 11818 14720
rect 11882 14656 11890 14720
rect 11570 13632 11890 14656
rect 11570 13568 11578 13632
rect 11642 13568 11658 13632
rect 11722 13568 11738 13632
rect 11802 13568 11818 13632
rect 11882 13568 11890 13632
rect 11570 12544 11890 13568
rect 11570 12480 11578 12544
rect 11642 12480 11658 12544
rect 11722 12480 11738 12544
rect 11802 12480 11818 12544
rect 11882 12480 11890 12544
rect 11570 11456 11890 12480
rect 11570 11392 11578 11456
rect 11642 11392 11658 11456
rect 11722 11392 11738 11456
rect 11802 11392 11818 11456
rect 11882 11392 11890 11456
rect 11570 10368 11890 11392
rect 11570 10304 11578 10368
rect 11642 10304 11658 10368
rect 11722 10304 11738 10368
rect 11802 10304 11818 10368
rect 11882 10304 11890 10368
rect 11570 9280 11890 10304
rect 11570 9216 11578 9280
rect 11642 9216 11658 9280
rect 11722 9216 11738 9280
rect 11802 9216 11818 9280
rect 11882 9216 11890 9280
rect 11570 8192 11890 9216
rect 11570 8128 11578 8192
rect 11642 8128 11658 8192
rect 11722 8128 11738 8192
rect 11802 8128 11818 8192
rect 11882 8128 11890 8192
rect 11570 7104 11890 8128
rect 11570 7040 11578 7104
rect 11642 7040 11658 7104
rect 11722 7040 11738 7104
rect 11802 7040 11818 7104
rect 11882 7040 11890 7104
rect 11570 6016 11890 7040
rect 11570 5952 11578 6016
rect 11642 5952 11658 6016
rect 11722 5952 11738 6016
rect 11802 5952 11818 6016
rect 11882 5952 11890 6016
rect 11570 4928 11890 5952
rect 11570 4864 11578 4928
rect 11642 4864 11658 4928
rect 11722 4864 11738 4928
rect 11802 4864 11818 4928
rect 11882 4864 11890 4928
rect 11570 3840 11890 4864
rect 11570 3776 11578 3840
rect 11642 3776 11658 3840
rect 11722 3776 11738 3840
rect 11802 3776 11818 3840
rect 11882 3776 11890 3840
rect 11570 2752 11890 3776
rect 11570 2688 11578 2752
rect 11642 2688 11658 2752
rect 11722 2688 11738 2752
rect 11802 2688 11818 2752
rect 11882 2688 11890 2752
rect 11570 2128 11890 2688
rect 15112 30496 15432 30512
rect 15112 30432 15120 30496
rect 15184 30432 15200 30496
rect 15264 30432 15280 30496
rect 15344 30432 15360 30496
rect 15424 30432 15432 30496
rect 15112 29408 15432 30432
rect 15112 29344 15120 29408
rect 15184 29344 15200 29408
rect 15264 29344 15280 29408
rect 15344 29344 15360 29408
rect 15424 29344 15432 29408
rect 15112 28320 15432 29344
rect 15112 28256 15120 28320
rect 15184 28256 15200 28320
rect 15264 28256 15280 28320
rect 15344 28256 15360 28320
rect 15424 28256 15432 28320
rect 15112 27232 15432 28256
rect 15112 27168 15120 27232
rect 15184 27168 15200 27232
rect 15264 27168 15280 27232
rect 15344 27168 15360 27232
rect 15424 27168 15432 27232
rect 15112 26144 15432 27168
rect 15112 26080 15120 26144
rect 15184 26080 15200 26144
rect 15264 26080 15280 26144
rect 15344 26080 15360 26144
rect 15424 26080 15432 26144
rect 15112 25056 15432 26080
rect 15112 24992 15120 25056
rect 15184 24992 15200 25056
rect 15264 24992 15280 25056
rect 15344 24992 15360 25056
rect 15424 24992 15432 25056
rect 15112 23968 15432 24992
rect 15112 23904 15120 23968
rect 15184 23904 15200 23968
rect 15264 23904 15280 23968
rect 15344 23904 15360 23968
rect 15424 23904 15432 23968
rect 15112 22880 15432 23904
rect 15112 22816 15120 22880
rect 15184 22816 15200 22880
rect 15264 22816 15280 22880
rect 15344 22816 15360 22880
rect 15424 22816 15432 22880
rect 15112 21792 15432 22816
rect 15112 21728 15120 21792
rect 15184 21728 15200 21792
rect 15264 21728 15280 21792
rect 15344 21728 15360 21792
rect 15424 21728 15432 21792
rect 15112 20704 15432 21728
rect 15112 20640 15120 20704
rect 15184 20640 15200 20704
rect 15264 20640 15280 20704
rect 15344 20640 15360 20704
rect 15424 20640 15432 20704
rect 15112 19616 15432 20640
rect 15112 19552 15120 19616
rect 15184 19552 15200 19616
rect 15264 19552 15280 19616
rect 15344 19552 15360 19616
rect 15424 19552 15432 19616
rect 15112 18528 15432 19552
rect 15112 18464 15120 18528
rect 15184 18464 15200 18528
rect 15264 18464 15280 18528
rect 15344 18464 15360 18528
rect 15424 18464 15432 18528
rect 15112 17440 15432 18464
rect 15112 17376 15120 17440
rect 15184 17376 15200 17440
rect 15264 17376 15280 17440
rect 15344 17376 15360 17440
rect 15424 17376 15432 17440
rect 15112 16352 15432 17376
rect 15112 16288 15120 16352
rect 15184 16288 15200 16352
rect 15264 16288 15280 16352
rect 15344 16288 15360 16352
rect 15424 16288 15432 16352
rect 15112 15264 15432 16288
rect 15112 15200 15120 15264
rect 15184 15200 15200 15264
rect 15264 15200 15280 15264
rect 15344 15200 15360 15264
rect 15424 15200 15432 15264
rect 15112 14176 15432 15200
rect 15112 14112 15120 14176
rect 15184 14112 15200 14176
rect 15264 14112 15280 14176
rect 15344 14112 15360 14176
rect 15424 14112 15432 14176
rect 15112 13088 15432 14112
rect 15112 13024 15120 13088
rect 15184 13024 15200 13088
rect 15264 13024 15280 13088
rect 15344 13024 15360 13088
rect 15424 13024 15432 13088
rect 15112 12000 15432 13024
rect 15112 11936 15120 12000
rect 15184 11936 15200 12000
rect 15264 11936 15280 12000
rect 15344 11936 15360 12000
rect 15424 11936 15432 12000
rect 15112 10912 15432 11936
rect 15112 10848 15120 10912
rect 15184 10848 15200 10912
rect 15264 10848 15280 10912
rect 15344 10848 15360 10912
rect 15424 10848 15432 10912
rect 15112 9824 15432 10848
rect 15112 9760 15120 9824
rect 15184 9760 15200 9824
rect 15264 9760 15280 9824
rect 15344 9760 15360 9824
rect 15424 9760 15432 9824
rect 15112 8736 15432 9760
rect 15112 8672 15120 8736
rect 15184 8672 15200 8736
rect 15264 8672 15280 8736
rect 15344 8672 15360 8736
rect 15424 8672 15432 8736
rect 15112 7648 15432 8672
rect 15112 7584 15120 7648
rect 15184 7584 15200 7648
rect 15264 7584 15280 7648
rect 15344 7584 15360 7648
rect 15424 7584 15432 7648
rect 15112 6560 15432 7584
rect 15112 6496 15120 6560
rect 15184 6496 15200 6560
rect 15264 6496 15280 6560
rect 15344 6496 15360 6560
rect 15424 6496 15432 6560
rect 15112 5472 15432 6496
rect 15112 5408 15120 5472
rect 15184 5408 15200 5472
rect 15264 5408 15280 5472
rect 15344 5408 15360 5472
rect 15424 5408 15432 5472
rect 15112 4384 15432 5408
rect 15112 4320 15120 4384
rect 15184 4320 15200 4384
rect 15264 4320 15280 4384
rect 15344 4320 15360 4384
rect 15424 4320 15432 4384
rect 15112 3296 15432 4320
rect 15112 3232 15120 3296
rect 15184 3232 15200 3296
rect 15264 3232 15280 3296
rect 15344 3232 15360 3296
rect 15424 3232 15432 3296
rect 15112 2208 15432 3232
rect 15112 2144 15120 2208
rect 15184 2144 15200 2208
rect 15264 2144 15280 2208
rect 15344 2144 15360 2208
rect 15424 2144 15432 2208
rect 15112 2128 15432 2144
rect 18654 29952 18974 30512
rect 18654 29888 18662 29952
rect 18726 29888 18742 29952
rect 18806 29888 18822 29952
rect 18886 29888 18902 29952
rect 18966 29888 18974 29952
rect 18654 28864 18974 29888
rect 18654 28800 18662 28864
rect 18726 28800 18742 28864
rect 18806 28800 18822 28864
rect 18886 28800 18902 28864
rect 18966 28800 18974 28864
rect 18654 27776 18974 28800
rect 18654 27712 18662 27776
rect 18726 27712 18742 27776
rect 18806 27712 18822 27776
rect 18886 27712 18902 27776
rect 18966 27712 18974 27776
rect 18654 26688 18974 27712
rect 18654 26624 18662 26688
rect 18726 26624 18742 26688
rect 18806 26624 18822 26688
rect 18886 26624 18902 26688
rect 18966 26624 18974 26688
rect 18654 25600 18974 26624
rect 18654 25536 18662 25600
rect 18726 25536 18742 25600
rect 18806 25536 18822 25600
rect 18886 25536 18902 25600
rect 18966 25536 18974 25600
rect 18654 24512 18974 25536
rect 18654 24448 18662 24512
rect 18726 24448 18742 24512
rect 18806 24448 18822 24512
rect 18886 24448 18902 24512
rect 18966 24448 18974 24512
rect 18654 23424 18974 24448
rect 18654 23360 18662 23424
rect 18726 23360 18742 23424
rect 18806 23360 18822 23424
rect 18886 23360 18902 23424
rect 18966 23360 18974 23424
rect 18654 22336 18974 23360
rect 22196 30496 22516 30512
rect 22196 30432 22204 30496
rect 22268 30432 22284 30496
rect 22348 30432 22364 30496
rect 22428 30432 22444 30496
rect 22508 30432 22516 30496
rect 22196 29408 22516 30432
rect 22196 29344 22204 29408
rect 22268 29344 22284 29408
rect 22348 29344 22364 29408
rect 22428 29344 22444 29408
rect 22508 29344 22516 29408
rect 22196 28320 22516 29344
rect 22196 28256 22204 28320
rect 22268 28256 22284 28320
rect 22348 28256 22364 28320
rect 22428 28256 22444 28320
rect 22508 28256 22516 28320
rect 22196 27232 22516 28256
rect 22196 27168 22204 27232
rect 22268 27168 22284 27232
rect 22348 27168 22364 27232
rect 22428 27168 22444 27232
rect 22508 27168 22516 27232
rect 22196 26144 22516 27168
rect 25738 29952 26058 30512
rect 25738 29888 25746 29952
rect 25810 29888 25826 29952
rect 25890 29888 25906 29952
rect 25970 29888 25986 29952
rect 26050 29888 26058 29952
rect 25738 28864 26058 29888
rect 29280 30496 29600 30512
rect 29280 30432 29288 30496
rect 29352 30432 29368 30496
rect 29432 30432 29448 30496
rect 29512 30432 29528 30496
rect 29592 30432 29600 30496
rect 29280 29408 29600 30432
rect 29280 29344 29288 29408
rect 29352 29344 29368 29408
rect 29432 29344 29448 29408
rect 29512 29344 29528 29408
rect 29592 29344 29600 29408
rect 27843 29340 27909 29341
rect 27843 29276 27844 29340
rect 27908 29276 27909 29340
rect 27843 29275 27909 29276
rect 25738 28800 25746 28864
rect 25810 28800 25826 28864
rect 25890 28800 25906 28864
rect 25970 28800 25986 28864
rect 26050 28800 26058 28864
rect 25738 27776 26058 28800
rect 25738 27712 25746 27776
rect 25810 27712 25826 27776
rect 25890 27712 25906 27776
rect 25970 27712 25986 27776
rect 26050 27712 26058 27776
rect 25738 26688 26058 27712
rect 25738 26624 25746 26688
rect 25810 26624 25826 26688
rect 25890 26624 25906 26688
rect 25970 26624 25986 26688
rect 26050 26624 26058 26688
rect 22691 26348 22757 26349
rect 22691 26284 22692 26348
rect 22756 26284 22757 26348
rect 22691 26283 22757 26284
rect 22196 26080 22204 26144
rect 22268 26080 22284 26144
rect 22348 26080 22364 26144
rect 22428 26080 22444 26144
rect 22508 26080 22516 26144
rect 22196 25056 22516 26080
rect 22196 24992 22204 25056
rect 22268 24992 22284 25056
rect 22348 24992 22364 25056
rect 22428 24992 22444 25056
rect 22508 24992 22516 25056
rect 22196 23968 22516 24992
rect 22196 23904 22204 23968
rect 22268 23904 22284 23968
rect 22348 23904 22364 23968
rect 22428 23904 22444 23968
rect 22508 23904 22516 23968
rect 21035 22948 21101 22949
rect 21035 22884 21036 22948
rect 21100 22884 21101 22948
rect 21035 22883 21101 22884
rect 18654 22272 18662 22336
rect 18726 22272 18742 22336
rect 18806 22272 18822 22336
rect 18886 22272 18902 22336
rect 18966 22272 18974 22336
rect 18654 21248 18974 22272
rect 18654 21184 18662 21248
rect 18726 21184 18742 21248
rect 18806 21184 18822 21248
rect 18886 21184 18902 21248
rect 18966 21184 18974 21248
rect 18654 20160 18974 21184
rect 18654 20096 18662 20160
rect 18726 20096 18742 20160
rect 18806 20096 18822 20160
rect 18886 20096 18902 20160
rect 18966 20096 18974 20160
rect 18654 19072 18974 20096
rect 18654 19008 18662 19072
rect 18726 19008 18742 19072
rect 18806 19008 18822 19072
rect 18886 19008 18902 19072
rect 18966 19008 18974 19072
rect 18654 17984 18974 19008
rect 18654 17920 18662 17984
rect 18726 17920 18742 17984
rect 18806 17920 18822 17984
rect 18886 17920 18902 17984
rect 18966 17920 18974 17984
rect 18654 16896 18974 17920
rect 18654 16832 18662 16896
rect 18726 16832 18742 16896
rect 18806 16832 18822 16896
rect 18886 16832 18902 16896
rect 18966 16832 18974 16896
rect 18654 15808 18974 16832
rect 20667 16692 20733 16693
rect 20667 16628 20668 16692
rect 20732 16628 20733 16692
rect 20667 16627 20733 16628
rect 18654 15744 18662 15808
rect 18726 15744 18742 15808
rect 18806 15744 18822 15808
rect 18886 15744 18902 15808
rect 18966 15744 18974 15808
rect 18654 14720 18974 15744
rect 18654 14656 18662 14720
rect 18726 14656 18742 14720
rect 18806 14656 18822 14720
rect 18886 14656 18902 14720
rect 18966 14656 18974 14720
rect 18654 13632 18974 14656
rect 18654 13568 18662 13632
rect 18726 13568 18742 13632
rect 18806 13568 18822 13632
rect 18886 13568 18902 13632
rect 18966 13568 18974 13632
rect 18654 12544 18974 13568
rect 18654 12480 18662 12544
rect 18726 12480 18742 12544
rect 18806 12480 18822 12544
rect 18886 12480 18902 12544
rect 18966 12480 18974 12544
rect 18654 11456 18974 12480
rect 20670 12205 20730 16627
rect 21038 13021 21098 22883
rect 22196 22880 22516 23904
rect 22196 22816 22204 22880
rect 22268 22816 22284 22880
rect 22348 22816 22364 22880
rect 22428 22816 22444 22880
rect 22508 22816 22516 22880
rect 22196 21792 22516 22816
rect 22196 21728 22204 21792
rect 22268 21728 22284 21792
rect 22348 21728 22364 21792
rect 22428 21728 22444 21792
rect 22508 21728 22516 21792
rect 22196 20704 22516 21728
rect 22196 20640 22204 20704
rect 22268 20640 22284 20704
rect 22348 20640 22364 20704
rect 22428 20640 22444 20704
rect 22508 20640 22516 20704
rect 22196 19616 22516 20640
rect 22196 19552 22204 19616
rect 22268 19552 22284 19616
rect 22348 19552 22364 19616
rect 22428 19552 22444 19616
rect 22508 19552 22516 19616
rect 22196 18528 22516 19552
rect 22196 18464 22204 18528
rect 22268 18464 22284 18528
rect 22348 18464 22364 18528
rect 22428 18464 22444 18528
rect 22508 18464 22516 18528
rect 22196 17440 22516 18464
rect 22196 17376 22204 17440
rect 22268 17376 22284 17440
rect 22348 17376 22364 17440
rect 22428 17376 22444 17440
rect 22508 17376 22516 17440
rect 22196 16352 22516 17376
rect 22196 16288 22204 16352
rect 22268 16288 22284 16352
rect 22348 16288 22364 16352
rect 22428 16288 22444 16352
rect 22508 16288 22516 16352
rect 22196 15264 22516 16288
rect 22196 15200 22204 15264
rect 22268 15200 22284 15264
rect 22348 15200 22364 15264
rect 22428 15200 22444 15264
rect 22508 15200 22516 15264
rect 22196 14176 22516 15200
rect 22196 14112 22204 14176
rect 22268 14112 22284 14176
rect 22348 14112 22364 14176
rect 22428 14112 22444 14176
rect 22508 14112 22516 14176
rect 22196 13088 22516 14112
rect 22196 13024 22204 13088
rect 22268 13024 22284 13088
rect 22348 13024 22364 13088
rect 22428 13024 22444 13088
rect 22508 13024 22516 13088
rect 21035 13020 21101 13021
rect 21035 12956 21036 13020
rect 21100 12956 21101 13020
rect 21035 12955 21101 12956
rect 20667 12204 20733 12205
rect 20667 12140 20668 12204
rect 20732 12140 20733 12204
rect 20667 12139 20733 12140
rect 18654 11392 18662 11456
rect 18726 11392 18742 11456
rect 18806 11392 18822 11456
rect 18886 11392 18902 11456
rect 18966 11392 18974 11456
rect 18654 10368 18974 11392
rect 18654 10304 18662 10368
rect 18726 10304 18742 10368
rect 18806 10304 18822 10368
rect 18886 10304 18902 10368
rect 18966 10304 18974 10368
rect 18654 9280 18974 10304
rect 18654 9216 18662 9280
rect 18726 9216 18742 9280
rect 18806 9216 18822 9280
rect 18886 9216 18902 9280
rect 18966 9216 18974 9280
rect 18654 8192 18974 9216
rect 18654 8128 18662 8192
rect 18726 8128 18742 8192
rect 18806 8128 18822 8192
rect 18886 8128 18902 8192
rect 18966 8128 18974 8192
rect 18654 7104 18974 8128
rect 18654 7040 18662 7104
rect 18726 7040 18742 7104
rect 18806 7040 18822 7104
rect 18886 7040 18902 7104
rect 18966 7040 18974 7104
rect 18654 6016 18974 7040
rect 18654 5952 18662 6016
rect 18726 5952 18742 6016
rect 18806 5952 18822 6016
rect 18886 5952 18902 6016
rect 18966 5952 18974 6016
rect 18654 4928 18974 5952
rect 18654 4864 18662 4928
rect 18726 4864 18742 4928
rect 18806 4864 18822 4928
rect 18886 4864 18902 4928
rect 18966 4864 18974 4928
rect 18654 3840 18974 4864
rect 18654 3776 18662 3840
rect 18726 3776 18742 3840
rect 18806 3776 18822 3840
rect 18886 3776 18902 3840
rect 18966 3776 18974 3840
rect 18654 2752 18974 3776
rect 18654 2688 18662 2752
rect 18726 2688 18742 2752
rect 18806 2688 18822 2752
rect 18886 2688 18902 2752
rect 18966 2688 18974 2752
rect 18654 2128 18974 2688
rect 22196 12000 22516 13024
rect 22196 11936 22204 12000
rect 22268 11936 22284 12000
rect 22348 11936 22364 12000
rect 22428 11936 22444 12000
rect 22508 11936 22516 12000
rect 22196 10912 22516 11936
rect 22196 10848 22204 10912
rect 22268 10848 22284 10912
rect 22348 10848 22364 10912
rect 22428 10848 22444 10912
rect 22508 10848 22516 10912
rect 22196 9824 22516 10848
rect 22196 9760 22204 9824
rect 22268 9760 22284 9824
rect 22348 9760 22364 9824
rect 22428 9760 22444 9824
rect 22508 9760 22516 9824
rect 22196 8736 22516 9760
rect 22196 8672 22204 8736
rect 22268 8672 22284 8736
rect 22348 8672 22364 8736
rect 22428 8672 22444 8736
rect 22508 8672 22516 8736
rect 22196 7648 22516 8672
rect 22694 7853 22754 26283
rect 25738 25600 26058 26624
rect 25738 25536 25746 25600
rect 25810 25536 25826 25600
rect 25890 25536 25906 25600
rect 25970 25536 25986 25600
rect 26050 25536 26058 25600
rect 25738 24512 26058 25536
rect 25738 24448 25746 24512
rect 25810 24448 25826 24512
rect 25890 24448 25906 24512
rect 25970 24448 25986 24512
rect 26050 24448 26058 24512
rect 25738 23424 26058 24448
rect 25738 23360 25746 23424
rect 25810 23360 25826 23424
rect 25890 23360 25906 23424
rect 25970 23360 25986 23424
rect 26050 23360 26058 23424
rect 25738 22336 26058 23360
rect 25738 22272 25746 22336
rect 25810 22272 25826 22336
rect 25890 22272 25906 22336
rect 25970 22272 25986 22336
rect 26050 22272 26058 22336
rect 25738 21248 26058 22272
rect 25738 21184 25746 21248
rect 25810 21184 25826 21248
rect 25890 21184 25906 21248
rect 25970 21184 25986 21248
rect 26050 21184 26058 21248
rect 25738 20160 26058 21184
rect 25738 20096 25746 20160
rect 25810 20096 25826 20160
rect 25890 20096 25906 20160
rect 25970 20096 25986 20160
rect 26050 20096 26058 20160
rect 25738 19072 26058 20096
rect 25738 19008 25746 19072
rect 25810 19008 25826 19072
rect 25890 19008 25906 19072
rect 25970 19008 25986 19072
rect 26050 19008 26058 19072
rect 25738 17984 26058 19008
rect 25738 17920 25746 17984
rect 25810 17920 25826 17984
rect 25890 17920 25906 17984
rect 25970 17920 25986 17984
rect 26050 17920 26058 17984
rect 25738 16896 26058 17920
rect 25738 16832 25746 16896
rect 25810 16832 25826 16896
rect 25890 16832 25906 16896
rect 25970 16832 25986 16896
rect 26050 16832 26058 16896
rect 25738 15808 26058 16832
rect 25738 15744 25746 15808
rect 25810 15744 25826 15808
rect 25890 15744 25906 15808
rect 25970 15744 25986 15808
rect 26050 15744 26058 15808
rect 25738 14720 26058 15744
rect 25738 14656 25746 14720
rect 25810 14656 25826 14720
rect 25890 14656 25906 14720
rect 25970 14656 25986 14720
rect 26050 14656 26058 14720
rect 25738 13632 26058 14656
rect 25738 13568 25746 13632
rect 25810 13568 25826 13632
rect 25890 13568 25906 13632
rect 25970 13568 25986 13632
rect 26050 13568 26058 13632
rect 25738 12544 26058 13568
rect 25738 12480 25746 12544
rect 25810 12480 25826 12544
rect 25890 12480 25906 12544
rect 25970 12480 25986 12544
rect 26050 12480 26058 12544
rect 25738 11456 26058 12480
rect 25738 11392 25746 11456
rect 25810 11392 25826 11456
rect 25890 11392 25906 11456
rect 25970 11392 25986 11456
rect 26050 11392 26058 11456
rect 25738 10368 26058 11392
rect 25738 10304 25746 10368
rect 25810 10304 25826 10368
rect 25890 10304 25906 10368
rect 25970 10304 25986 10368
rect 26050 10304 26058 10368
rect 25738 9280 26058 10304
rect 25738 9216 25746 9280
rect 25810 9216 25826 9280
rect 25890 9216 25906 9280
rect 25970 9216 25986 9280
rect 26050 9216 26058 9280
rect 25738 8192 26058 9216
rect 25738 8128 25746 8192
rect 25810 8128 25826 8192
rect 25890 8128 25906 8192
rect 25970 8128 25986 8192
rect 26050 8128 26058 8192
rect 22691 7852 22757 7853
rect 22691 7788 22692 7852
rect 22756 7788 22757 7852
rect 22691 7787 22757 7788
rect 22196 7584 22204 7648
rect 22268 7584 22284 7648
rect 22348 7584 22364 7648
rect 22428 7584 22444 7648
rect 22508 7584 22516 7648
rect 22196 6560 22516 7584
rect 22196 6496 22204 6560
rect 22268 6496 22284 6560
rect 22348 6496 22364 6560
rect 22428 6496 22444 6560
rect 22508 6496 22516 6560
rect 22196 5472 22516 6496
rect 22196 5408 22204 5472
rect 22268 5408 22284 5472
rect 22348 5408 22364 5472
rect 22428 5408 22444 5472
rect 22508 5408 22516 5472
rect 22196 4384 22516 5408
rect 22196 4320 22204 4384
rect 22268 4320 22284 4384
rect 22348 4320 22364 4384
rect 22428 4320 22444 4384
rect 22508 4320 22516 4384
rect 22196 3296 22516 4320
rect 22196 3232 22204 3296
rect 22268 3232 22284 3296
rect 22348 3232 22364 3296
rect 22428 3232 22444 3296
rect 22508 3232 22516 3296
rect 22196 2208 22516 3232
rect 22196 2144 22204 2208
rect 22268 2144 22284 2208
rect 22348 2144 22364 2208
rect 22428 2144 22444 2208
rect 22508 2144 22516 2208
rect 22196 2128 22516 2144
rect 25738 7104 26058 8128
rect 25738 7040 25746 7104
rect 25810 7040 25826 7104
rect 25890 7040 25906 7104
rect 25970 7040 25986 7104
rect 26050 7040 26058 7104
rect 25738 6016 26058 7040
rect 25738 5952 25746 6016
rect 25810 5952 25826 6016
rect 25890 5952 25906 6016
rect 25970 5952 25986 6016
rect 26050 5952 26058 6016
rect 25738 4928 26058 5952
rect 27846 5133 27906 29275
rect 29280 28320 29600 29344
rect 29280 28256 29288 28320
rect 29352 28256 29368 28320
rect 29432 28256 29448 28320
rect 29512 28256 29528 28320
rect 29592 28256 29600 28320
rect 29280 27232 29600 28256
rect 29280 27168 29288 27232
rect 29352 27168 29368 27232
rect 29432 27168 29448 27232
rect 29512 27168 29528 27232
rect 29592 27168 29600 27232
rect 29280 26144 29600 27168
rect 29280 26080 29288 26144
rect 29352 26080 29368 26144
rect 29432 26080 29448 26144
rect 29512 26080 29528 26144
rect 29592 26080 29600 26144
rect 29280 25056 29600 26080
rect 29280 24992 29288 25056
rect 29352 24992 29368 25056
rect 29432 24992 29448 25056
rect 29512 24992 29528 25056
rect 29592 24992 29600 25056
rect 29280 23968 29600 24992
rect 29280 23904 29288 23968
rect 29352 23904 29368 23968
rect 29432 23904 29448 23968
rect 29512 23904 29528 23968
rect 29592 23904 29600 23968
rect 29280 22880 29600 23904
rect 29280 22816 29288 22880
rect 29352 22816 29368 22880
rect 29432 22816 29448 22880
rect 29512 22816 29528 22880
rect 29592 22816 29600 22880
rect 29280 21792 29600 22816
rect 29280 21728 29288 21792
rect 29352 21728 29368 21792
rect 29432 21728 29448 21792
rect 29512 21728 29528 21792
rect 29592 21728 29600 21792
rect 29280 20704 29600 21728
rect 29280 20640 29288 20704
rect 29352 20640 29368 20704
rect 29432 20640 29448 20704
rect 29512 20640 29528 20704
rect 29592 20640 29600 20704
rect 29280 19616 29600 20640
rect 29280 19552 29288 19616
rect 29352 19552 29368 19616
rect 29432 19552 29448 19616
rect 29512 19552 29528 19616
rect 29592 19552 29600 19616
rect 29280 18528 29600 19552
rect 29280 18464 29288 18528
rect 29352 18464 29368 18528
rect 29432 18464 29448 18528
rect 29512 18464 29528 18528
rect 29592 18464 29600 18528
rect 29280 17440 29600 18464
rect 29280 17376 29288 17440
rect 29352 17376 29368 17440
rect 29432 17376 29448 17440
rect 29512 17376 29528 17440
rect 29592 17376 29600 17440
rect 29280 16352 29600 17376
rect 29280 16288 29288 16352
rect 29352 16288 29368 16352
rect 29432 16288 29448 16352
rect 29512 16288 29528 16352
rect 29592 16288 29600 16352
rect 29280 15264 29600 16288
rect 29280 15200 29288 15264
rect 29352 15200 29368 15264
rect 29432 15200 29448 15264
rect 29512 15200 29528 15264
rect 29592 15200 29600 15264
rect 29280 14176 29600 15200
rect 29280 14112 29288 14176
rect 29352 14112 29368 14176
rect 29432 14112 29448 14176
rect 29512 14112 29528 14176
rect 29592 14112 29600 14176
rect 29280 13088 29600 14112
rect 29280 13024 29288 13088
rect 29352 13024 29368 13088
rect 29432 13024 29448 13088
rect 29512 13024 29528 13088
rect 29592 13024 29600 13088
rect 29280 12000 29600 13024
rect 29280 11936 29288 12000
rect 29352 11936 29368 12000
rect 29432 11936 29448 12000
rect 29512 11936 29528 12000
rect 29592 11936 29600 12000
rect 29280 10912 29600 11936
rect 29280 10848 29288 10912
rect 29352 10848 29368 10912
rect 29432 10848 29448 10912
rect 29512 10848 29528 10912
rect 29592 10848 29600 10912
rect 29280 9824 29600 10848
rect 29280 9760 29288 9824
rect 29352 9760 29368 9824
rect 29432 9760 29448 9824
rect 29512 9760 29528 9824
rect 29592 9760 29600 9824
rect 29280 8736 29600 9760
rect 29280 8672 29288 8736
rect 29352 8672 29368 8736
rect 29432 8672 29448 8736
rect 29512 8672 29528 8736
rect 29592 8672 29600 8736
rect 29280 7648 29600 8672
rect 29280 7584 29288 7648
rect 29352 7584 29368 7648
rect 29432 7584 29448 7648
rect 29512 7584 29528 7648
rect 29592 7584 29600 7648
rect 29280 6560 29600 7584
rect 29280 6496 29288 6560
rect 29352 6496 29368 6560
rect 29432 6496 29448 6560
rect 29512 6496 29528 6560
rect 29592 6496 29600 6560
rect 29280 5472 29600 6496
rect 29280 5408 29288 5472
rect 29352 5408 29368 5472
rect 29432 5408 29448 5472
rect 29512 5408 29528 5472
rect 29592 5408 29600 5472
rect 27843 5132 27909 5133
rect 27843 5068 27844 5132
rect 27908 5068 27909 5132
rect 27843 5067 27909 5068
rect 25738 4864 25746 4928
rect 25810 4864 25826 4928
rect 25890 4864 25906 4928
rect 25970 4864 25986 4928
rect 26050 4864 26058 4928
rect 25738 3840 26058 4864
rect 25738 3776 25746 3840
rect 25810 3776 25826 3840
rect 25890 3776 25906 3840
rect 25970 3776 25986 3840
rect 26050 3776 26058 3840
rect 25738 2752 26058 3776
rect 25738 2688 25746 2752
rect 25810 2688 25826 2752
rect 25890 2688 25906 2752
rect 25970 2688 25986 2752
rect 26050 2688 26058 2752
rect 25738 2128 26058 2688
rect 29280 4384 29600 5408
rect 29280 4320 29288 4384
rect 29352 4320 29368 4384
rect 29432 4320 29448 4384
rect 29512 4320 29528 4384
rect 29592 4320 29600 4384
rect 29280 3296 29600 4320
rect 29280 3232 29288 3296
rect 29352 3232 29368 3296
rect 29432 3232 29448 3296
rect 29512 3232 29528 3296
rect 29592 3232 29600 3296
rect 29280 2208 29600 3232
rect 29280 2144 29288 2208
rect 29352 2144 29368 2208
rect 29432 2144 29448 2208
rect 29512 2144 29528 2208
rect 29592 2144 29600 2208
rect 29280 2128 29600 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__A opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19412 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__A
timestamp 1649977179
transform 1 0 18584 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__B
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__D
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__C
timestamp 1649977179
transform -1 0 26220 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__D
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__A
timestamp 1649977179
transform -1 0 25668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__A
timestamp 1649977179
transform -1 0 18768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__B
timestamp 1649977179
transform 1 0 19688 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__C
timestamp 1649977179
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__D
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A
timestamp 1649977179
transform 1 0 16560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__B
timestamp 1649977179
transform 1 0 17756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__C
timestamp 1649977179
transform -1 0 20332 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__D
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A
timestamp 1649977179
transform -1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__B
timestamp 1649977179
transform -1 0 20884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__A
timestamp 1649977179
transform -1 0 22724 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__A1
timestamp 1649977179
transform 1 0 20056 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__B1
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__C1
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__A1
timestamp 1649977179
transform 1 0 21160 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__A
timestamp 1649977179
transform -1 0 27692 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A
timestamp 1649977179
transform -1 0 26864 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__C
timestamp 1649977179
transform 1 0 25944 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__D
timestamp 1649977179
transform 1 0 24288 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__A
timestamp 1649977179
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A
timestamp 1649977179
transform 1 0 13524 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__A
timestamp 1649977179
transform -1 0 20240 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__B
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__C
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A1
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__S
timestamp 1649977179
transform -1 0 20148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A0
timestamp 1649977179
transform 1 0 19136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A1
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__S
timestamp 1649977179
transform 1 0 18584 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A
timestamp 1649977179
transform 1 0 20148 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__S
timestamp 1649977179
transform 1 0 18768 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__A0
timestamp 1649977179
transform -1 0 16468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__A1
timestamp 1649977179
transform 1 0 16836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__S
timestamp 1649977179
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A0
timestamp 1649977179
transform 1 0 15456 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A1
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__S
timestamp 1649977179
transform 1 0 17848 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__S
timestamp 1649977179
transform 1 0 17480 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__A
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__B1
timestamp 1649977179
transform -1 0 21252 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A
timestamp 1649977179
transform 1 0 15640 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__A0
timestamp 1649977179
transform 1 0 20608 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__A1
timestamp 1649977179
transform -1 0 21988 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__S
timestamp 1649977179
transform 1 0 20056 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__A
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__B
timestamp 1649977179
transform -1 0 20516 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A1
timestamp 1649977179
transform -1 0 21068 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A2
timestamp 1649977179
transform 1 0 19780 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__C1
timestamp 1649977179
transform 1 0 20516 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__A1
timestamp 1649977179
transform 1 0 19228 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A0
timestamp 1649977179
transform 1 0 16008 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A1
timestamp 1649977179
transform 1 0 15456 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__S
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A
timestamp 1649977179
transform -1 0 27876 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A0
timestamp 1649977179
transform 1 0 20148 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A1
timestamp 1649977179
transform 1 0 19044 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__S
timestamp 1649977179
transform 1 0 19596 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__S
timestamp 1649977179
transform 1 0 17756 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__A
timestamp 1649977179
transform -1 0 23460 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__B
timestamp 1649977179
transform 1 0 23920 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A1
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A2
timestamp 1649977179
transform 1 0 23460 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__B2
timestamp 1649977179
transform 1 0 23644 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A1
timestamp 1649977179
transform 1 0 18768 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__A2
timestamp 1649977179
transform 1 0 26312 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__B
timestamp 1649977179
transform 1 0 23276 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B
timestamp 1649977179
transform -1 0 21436 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A1
timestamp 1649977179
transform -1 0 23920 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A
timestamp 1649977179
transform 1 0 25024 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A2_N
timestamp 1649977179
transform -1 0 25208 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A
timestamp 1649977179
transform 1 0 14076 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1649977179
transform -1 0 23184 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__B
timestamp 1649977179
transform 1 0 22356 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A
timestamp 1649977179
transform 1 0 22264 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 1649977179
transform 1 0 23368 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B
timestamp 1649977179
transform 1 0 22356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A1
timestamp 1649977179
transform 1 0 21804 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__B
timestamp 1649977179
transform 1 0 21160 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A1
timestamp 1649977179
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A2
timestamp 1649977179
transform 1 0 20884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A
timestamp 1649977179
transform 1 0 24288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B
timestamp 1649977179
transform 1 0 23552 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A2
timestamp 1649977179
transform -1 0 20884 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__S
timestamp 1649977179
transform 1 0 19320 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1649977179
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__B
timestamp 1649977179
transform 1 0 13064 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A0
timestamp 1649977179
transform 1 0 21160 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A1
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A2
timestamp 1649977179
transform 1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A3
timestamp 1649977179
transform 1 0 23000 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__S1
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A0
timestamp 1649977179
transform 1 0 26312 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A1
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A2
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A3
timestamp 1649977179
transform 1 0 26036 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__S1
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1649977179
transform 1 0 23644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B
timestamp 1649977179
transform 1 0 24656 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1649977179
transform 1 0 23736 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A1
timestamp 1649977179
transform -1 0 23552 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A2
timestamp 1649977179
transform -1 0 23736 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__B
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1649977179
transform 1 0 13892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A
timestamp 1649977179
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 1649977179
transform -1 0 23000 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A1
timestamp 1649977179
transform -1 0 21344 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A
timestamp 1649977179
transform 1 0 20332 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A1
timestamp 1649977179
transform -1 0 20884 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B
timestamp 1649977179
transform 1 0 21160 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B
timestamp 1649977179
transform 1 0 21252 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A1
timestamp 1649977179
transform -1 0 21620 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A2
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B1
timestamp 1649977179
transform -1 0 22724 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__C1
timestamp 1649977179
transform 1 0 21988 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1649977179
transform 1 0 22356 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__B
timestamp 1649977179
transform 1 0 20700 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A2
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__B1
timestamp 1649977179
transform 1 0 20148 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A1
timestamp 1649977179
transform -1 0 20792 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B1
timestamp 1649977179
transform 1 0 23092 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B2
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A2
timestamp 1649977179
transform 1 0 17940 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A3
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1649977179
transform 1 0 13432 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B
timestamp 1649977179
transform 1 0 14076 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1649977179
transform 1 0 14812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B
timestamp 1649977179
transform 1 0 16192 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A
timestamp 1649977179
transform -1 0 17664 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A1
timestamp 1649977179
transform -1 0 17204 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A
timestamp 1649977179
transform 1 0 12420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1649977179
transform 1 0 11224 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A2
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__B1
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__C1
timestamp 1649977179
transform 1 0 17204 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A1
timestamp 1649977179
transform -1 0 16376 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A2
timestamp 1649977179
transform 1 0 16744 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B2
timestamp 1649977179
transform 1 0 15640 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__S
timestamp 1649977179
transform 1 0 18032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A1
timestamp 1649977179
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B1
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__C1
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__S
timestamp 1649977179
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A1
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A0
timestamp 1649977179
transform 1 0 26036 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A1
timestamp 1649977179
transform 1 0 22724 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1
timestamp 1649977179
transform 1 0 17664 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A3
timestamp 1649977179
transform -1 0 18400 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B2
timestamp 1649977179
transform 1 0 18308 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A
timestamp 1649977179
transform -1 0 9844 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__B
timestamp 1649977179
transform -1 0 11224 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A
timestamp 1649977179
transform 1 0 10856 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B
timestamp 1649977179
transform -1 0 9936 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A
timestamp 1649977179
transform 1 0 12144 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B
timestamp 1649977179
transform 1 0 12696 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1
timestamp 1649977179
transform 1 0 10856 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A2
timestamp 1649977179
transform -1 0 9568 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B1
timestamp 1649977179
transform 1 0 10304 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A1
timestamp 1649977179
transform 1 0 12788 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__C1
timestamp 1649977179
transform 1 0 13156 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A1
timestamp 1649977179
transform 1 0 13064 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A2
timestamp 1649977179
transform 1 0 10212 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B
timestamp 1649977179
transform 1 0 13432 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A1
timestamp 1649977179
transform 1 0 17296 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A
timestamp 1649977179
transform 1 0 14444 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A1
timestamp 1649977179
transform 1 0 13892 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__S
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__S
timestamp 1649977179
transform 1 0 17848 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A0
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A1
timestamp 1649977179
transform -1 0 27692 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A2
timestamp 1649977179
transform -1 0 28796 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A3
timestamp 1649977179
transform 1 0 27232 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__S1
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A0
timestamp 1649977179
transform -1 0 17480 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A1
timestamp 1649977179
transform 1 0 16008 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__S
timestamp 1649977179
transform 1 0 17664 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A1
timestamp 1649977179
transform 1 0 21160 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A2
timestamp 1649977179
transform 1 0 20148 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A1
timestamp 1649977179
transform 1 0 18216 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A0
timestamp 1649977179
transform 1 0 27968 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A1
timestamp 1649977179
transform 1 0 27784 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__S
timestamp 1649977179
transform -1 0 27140 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A
timestamp 1649977179
transform 1 0 23736 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A
timestamp 1649977179
transform 1 0 17848 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B
timestamp 1649977179
transform 1 0 18400 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A0
timestamp 1649977179
transform 1 0 28520 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A1
timestamp 1649977179
transform 1 0 28336 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1649977179
transform 1 0 19320 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A
timestamp 1649977179
transform 1 0 9200 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B
timestamp 1649977179
transform 1 0 8372 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A
timestamp 1649977179
transform 1 0 7544 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B
timestamp 1649977179
transform -1 0 8280 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B
timestamp 1649977179
transform 1 0 12420 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A
timestamp 1649977179
transform 1 0 5152 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A
timestamp 1649977179
transform 1 0 12420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A1
timestamp 1649977179
transform 1 0 10672 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A2
timestamp 1649977179
transform -1 0 9752 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B2
timestamp 1649977179
transform -1 0 9384 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A1
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A2
timestamp 1649977179
transform 1 0 12052 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B1
timestamp 1649977179
transform 1 0 11040 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__C1
timestamp 1649977179
transform 1 0 10304 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A1
timestamp 1649977179
transform 1 0 8280 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A1
timestamp 1649977179
transform -1 0 8096 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A2
timestamp 1649977179
transform -1 0 8464 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A
timestamp 1649977179
transform 1 0 8740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A
timestamp 1649977179
transform 1 0 10488 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B
timestamp 1649977179
transform 1 0 11408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A
timestamp 1649977179
transform 1 0 6716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B
timestamp 1649977179
transform 1 0 7912 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A2
timestamp 1649977179
transform -1 0 7084 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__B
timestamp 1649977179
transform -1 0 5796 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1649977179
transform 1 0 6164 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A0
timestamp 1649977179
transform -1 0 28336 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A1
timestamp 1649977179
transform -1 0 28796 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A
timestamp 1649977179
transform 1 0 9568 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B
timestamp 1649977179
transform 1 0 9292 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B1
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1649977179
transform -1 0 12144 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A0
timestamp 1649977179
transform 1 0 10672 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A1
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A1
timestamp 1649977179
transform 1 0 7728 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A2
timestamp 1649977179
transform -1 0 10764 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B1
timestamp 1649977179
transform -1 0 8464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A1
timestamp 1649977179
transform 1 0 8648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A2
timestamp 1649977179
transform 1 0 10120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A
timestamp 1649977179
transform 1 0 8188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A
timestamp 1649977179
transform 1 0 8280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__B
timestamp 1649977179
transform 1 0 9108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A
timestamp 1649977179
transform 1 0 8188 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B
timestamp 1649977179
transform 1 0 8280 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A1
timestamp 1649977179
transform -1 0 5888 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A2
timestamp 1649977179
transform -1 0 5336 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A
timestamp 1649977179
transform -1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__B
timestamp 1649977179
transform 1 0 6532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A1
timestamp 1649977179
transform -1 0 7084 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A2
timestamp 1649977179
transform 1 0 8188 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1649977179
transform -1 0 5888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A0
timestamp 1649977179
transform 1 0 27232 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A1
timestamp 1649977179
transform 1 0 28244 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A0
timestamp 1649977179
transform -1 0 23644 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A
timestamp 1649977179
transform 1 0 5152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__B
timestamp 1649977179
transform 1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A1
timestamp 1649977179
transform 1 0 8004 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A2
timestamp 1649977179
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__B1
timestamp 1649977179
transform 1 0 10304 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A1
timestamp 1649977179
transform -1 0 10396 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__C1
timestamp 1649977179
transform 1 0 11960 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A1_N
timestamp 1649977179
transform 1 0 9108 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A2_N
timestamp 1649977179
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A1
timestamp 1649977179
transform 1 0 11500 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A1
timestamp 1649977179
transform -1 0 4784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B
timestamp 1649977179
transform 1 0 8280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A
timestamp 1649977179
transform 1 0 6992 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B
timestamp 1649977179
transform -1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A0
timestamp 1649977179
transform 1 0 26312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A1
timestamp 1649977179
transform 1 0 26864 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__S
timestamp 1649977179
transform 1 0 28244 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A1
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A2
timestamp 1649977179
transform 1 0 10488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B1
timestamp 1649977179
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__C1
timestamp 1649977179
transform 1 0 10396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1649977179
transform 1 0 9108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__C
timestamp 1649977179
transform 1 0 9936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A1
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A2
timestamp 1649977179
transform -1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A1
timestamp 1649977179
transform 1 0 12052 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A
timestamp 1649977179
transform 1 0 1932 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A1
timestamp 1649977179
transform 1 0 3220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A
timestamp 1649977179
transform 1 0 1656 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__C1
timestamp 1649977179
transform 1 0 4600 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A1
timestamp 1649977179
transform 1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1649977179
transform 1 0 9108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B
timestamp 1649977179
transform 1 0 9568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B
timestamp 1649977179
transform -1 0 9384 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1649977179
transform 1 0 5704 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__B
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A2
timestamp 1649977179
transform -1 0 5612 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__B
timestamp 1649977179
transform 1 0 4692 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 1649977179
transform 1 0 5520 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A0
timestamp 1649977179
transform 1 0 26864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A1
timestamp 1649977179
transform 1 0 26312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__S
timestamp 1649977179
transform -1 0 28796 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1649977179
transform 1 0 12052 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A2
timestamp 1649977179
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A3
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__B1
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1649977179
transform 1 0 21804 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A1
timestamp 1649977179
transform 1 0 10672 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A2
timestamp 1649977179
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__B1
timestamp 1649977179
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A1
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A2
timestamp 1649977179
transform 1 0 10764 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__B1
timestamp 1649977179
transform 1 0 12052 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__B1
timestamp 1649977179
transform 1 0 14996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A1
timestamp 1649977179
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A
timestamp 1649977179
transform 1 0 7912 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1649977179
transform 1 0 6532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A
timestamp 1649977179
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A0
timestamp 1649977179
transform -1 0 28704 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A1
timestamp 1649977179
transform 1 0 26036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__S
timestamp 1649977179
transform 1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__B
timestamp 1649977179
transform 1 0 23092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A1
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A2
timestamp 1649977179
transform -1 0 9476 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__B1
timestamp 1649977179
transform 1 0 9752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__C1
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__B
timestamp 1649977179
transform 1 0 10304 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__C
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A1
timestamp 1649977179
transform 1 0 10856 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A2
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__B1
timestamp 1649977179
transform 1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A1
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A1
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1649977179
transform 1 0 10120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__B
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1649977179
transform 1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__B
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1649977179
transform 1 0 7636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1649977179
transform 1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A2
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A1
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A2
timestamp 1649977179
transform -1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A
timestamp 1649977179
transform 1 0 7176 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B
timestamp 1649977179
transform 1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A0
timestamp 1649977179
transform 1 0 26312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__S
timestamp 1649977179
transform -1 0 27692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A1
timestamp 1649977179
transform 1 0 17388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A2
timestamp 1649977179
transform 1 0 17940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A0
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A1
timestamp 1649977179
transform 1 0 11040 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A1
timestamp 1649977179
transform 1 0 11408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A1
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A2
timestamp 1649977179
transform 1 0 12696 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B1
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1649977179
transform 1 0 8280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1649977179
transform 1 0 6440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A2
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1649977179
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B
timestamp 1649977179
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A
timestamp 1649977179
transform 1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__B
timestamp 1649977179
transform 1 0 9936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__B1
timestamp 1649977179
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A1
timestamp 1649977179
transform 1 0 27876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A2
timestamp 1649977179
transform 1 0 27140 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A
timestamp 1649977179
transform -1 0 26036 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A1
timestamp 1649977179
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A2
timestamp 1649977179
transform -1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B1
timestamp 1649977179
transform 1 0 9476 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A1
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A2
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__B2
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__C1
timestamp 1649977179
transform 1 0 11684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A1
timestamp 1649977179
transform -1 0 11224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A
timestamp 1649977179
transform -1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A2
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__B
timestamp 1649977179
transform -1 0 5888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__B1
timestamp 1649977179
transform 1 0 5612 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B
timestamp 1649977179
transform -1 0 13064 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A0
timestamp 1649977179
transform 1 0 27876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A1
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__S
timestamp 1649977179
transform -1 0 28796 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B
timestamp 1649977179
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1649977179
transform 1 0 14628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A1
timestamp 1649977179
transform -1 0 11960 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__B1
timestamp 1649977179
transform -1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A1
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A2
timestamp 1649977179
transform 1 0 11684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B1
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1649977179
transform 1 0 12144 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A2
timestamp 1649977179
transform 1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1
timestamp 1649977179
transform 1 0 10856 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B1
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A1
timestamp 1649977179
transform -1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A2
timestamp 1649977179
transform 1 0 14628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B1
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B
timestamp 1649977179
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A
timestamp 1649977179
transform 1 0 16560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__B
timestamp 1649977179
transform 1 0 17112 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A
timestamp 1649977179
transform 1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A2
timestamp 1649977179
transform 1 0 16192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B
timestamp 1649977179
transform 1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1649977179
transform 1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A1
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A2
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B1
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__C1
timestamp 1649977179
transform 1 0 15640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__B
timestamp 1649977179
transform 1 0 15364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A1
timestamp 1649977179
transform 1 0 15824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A2
timestamp 1649977179
transform 1 0 17112 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__B2
timestamp 1649977179
transform 1 0 15272 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__C1
timestamp 1649977179
transform 1 0 16560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A1
timestamp 1649977179
transform -1 0 14628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A
timestamp 1649977179
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A
timestamp 1649977179
transform 1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A
timestamp 1649977179
transform 1 0 20976 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__B1
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A
timestamp 1649977179
transform 1 0 16744 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A
timestamp 1649977179
transform -1 0 19688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A2
timestamp 1649977179
transform 1 0 17756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A1
timestamp 1649977179
transform -1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A1
timestamp 1649977179
transform 1 0 21160 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A2
timestamp 1649977179
transform 1 0 17756 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__B1
timestamp 1649977179
transform -1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__C1
timestamp 1649977179
transform -1 0 17848 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A2
timestamp 1649977179
transform 1 0 20424 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__B2
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__C1
timestamp 1649977179
transform -1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1649977179
transform 1 0 24748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__S
timestamp 1649977179
transform -1 0 25944 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A
timestamp 1649977179
transform 1 0 16928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A1
timestamp 1649977179
transform 1 0 18032 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1649977179
transform 1 0 21160 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1649977179
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__B
timestamp 1649977179
transform 1 0 23184 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__B
timestamp 1649977179
transform 1 0 24104 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A
timestamp 1649977179
transform 1 0 21804 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A1
timestamp 1649977179
transform 1 0 23092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A1
timestamp 1649977179
transform 1 0 25024 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A1
timestamp 1649977179
transform 1 0 20424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A2
timestamp 1649977179
transform 1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__B1
timestamp 1649977179
transform -1 0 20056 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__C1
timestamp 1649977179
transform -1 0 19780 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A1
timestamp 1649977179
transform 1 0 23552 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A2
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A3
timestamp 1649977179
transform -1 0 23092 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__B1
timestamp 1649977179
transform 1 0 23460 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1649977179
transform -1 0 23184 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A1
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A2
timestamp 1649977179
transform 1 0 24656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A
timestamp 1649977179
transform -1 0 2944 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__B
timestamp 1649977179
transform 1 0 2392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A
timestamp 1649977179
transform 1 0 2760 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__B
timestamp 1649977179
transform 1 0 10120 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1649977179
transform -1 0 9384 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__B
timestamp 1649977179
transform 1 0 9568 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A
timestamp 1649977179
transform 1 0 2392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B
timestamp 1649977179
transform 1 0 2760 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__B2
timestamp 1649977179
transform 1 0 20976 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1649977179
transform -1 0 26128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A1
timestamp 1649977179
transform -1 0 24564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A1
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__B1
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__B1
timestamp 1649977179
transform -1 0 21988 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A1
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A
timestamp 1649977179
transform 1 0 2576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__A
timestamp 1649977179
transform -1 0 3956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__B
timestamp 1649977179
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A
timestamp 1649977179
transform 1 0 9200 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__B
timestamp 1649977179
transform 1 0 10488 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__C
timestamp 1649977179
transform 1 0 9936 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__D
timestamp 1649977179
transform -1 0 10212 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A
timestamp 1649977179
transform -1 0 8188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__B
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__C
timestamp 1649977179
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__D
timestamp 1649977179
transform 1 0 2944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__A
timestamp 1649977179
transform -1 0 24932 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A
timestamp 1649977179
transform -1 0 23552 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A
timestamp 1649977179
transform 1 0 21988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A1
timestamp 1649977179
transform -1 0 24564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A2
timestamp 1649977179
transform -1 0 23920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A
timestamp 1649977179
transform 1 0 2852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 17020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 19412 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 28796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 1656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 28796 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 28796 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 2668 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 28796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 28796 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 27416 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 28796 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 1748 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 1748 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 15180 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 2208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 22908 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 1564 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 28060 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 28796 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 19964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 24564 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 24840 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 28060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 1564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 28796 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 27140 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 21344 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 6808 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 13616 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 3220 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 20056 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output39_A
timestamp 1649977179
transform -1 0 2300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output40_A
timestamp 1649977179
transform 1 0 27508 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output42_A
timestamp 1649977179
transform -1 0 28152 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output43_A
timestamp 1649977179
transform -1 0 27324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output44_A
timestamp 1649977179
transform 1 0 11500 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output45_A
timestamp 1649977179
transform -1 0 27876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output48_A
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output50_A
timestamp 1649977179
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output51_A
timestamp 1649977179
transform 1 0 28244 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output52_A
timestamp 1649977179
transform 1 0 26312 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output55_A
timestamp 1649977179
transform -1 0 21988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output58_A
timestamp 1649977179
transform -1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35
timestamp 1649977179
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61
timestamp 1649977179
transform 1 0 6716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1649977179
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1649977179
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154
timestamp 1649977179
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1649977179
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_177
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1649977179
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_207
timestamp 1649977179
transform 1 0 20148 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_213
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1649977179
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_229
timestamp 1649977179
transform 1 0 22172 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1649977179
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1649977179
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_266
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1649977179
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1649977179
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_296
timestamp 1649977179
transform 1 0 28336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_7
timestamp 1649977179
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1649977179
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_99
timestamp 1649977179
transform 1 0 10212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_119
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_128
timestamp 1649977179
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_136
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1649977179
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_153
timestamp 1649977179
transform 1 0 15180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1649977179
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_186
timestamp 1649977179
transform 1 0 18216 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_214
timestamp 1649977179
transform 1 0 20792 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_227
timestamp 1649977179
transform 1 0 21988 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_239
timestamp 1649977179
transform 1 0 23092 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_244
timestamp 1649977179
transform 1 0 23552 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_256
timestamp 1649977179
transform 1 0 24656 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_268
timestamp 1649977179
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_285
timestamp 1649977179
transform 1 0 27324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_301
timestamp 1649977179
transform 1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19
timestamp 1649977179
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1649977179
transform 1 0 12052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_126
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_148
timestamp 1649977179
transform 1 0 14720 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_161
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1649977179
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_183
timestamp 1649977179
transform 1 0 17940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1649977179
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_211
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_217
timestamp 1649977179
transform 1 0 21068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_225
timestamp 1649977179
transform 1 0 21804 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_232
timestamp 1649977179
transform 1 0 22448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_236
timestamp 1649977179
transform 1 0 22816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1649977179
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1649977179
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_255
timestamp 1649977179
transform 1 0 24564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_267
timestamp 1649977179
transform 1 0 25668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_279
timestamp 1649977179
transform 1 0 26772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_293
timestamp 1649977179
transform 1 0 28060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1649977179
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_21
timestamp 1649977179
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_33
timestamp 1649977179
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_45
timestamp 1649977179
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_102
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_116
timestamp 1649977179
transform 1 0 11776 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_122
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_132
timestamp 1649977179
transform 1 0 13248 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_140
timestamp 1649977179
transform 1 0 13984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1649977179
transform 1 0 15456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1649977179
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1649977179
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1649977179
transform 1 0 17572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_189
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_196
timestamp 1649977179
transform 1 0 19136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_202
timestamp 1649977179
transform 1 0 19688 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_210
timestamp 1649977179
transform 1 0 20424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1649977179
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_231
timestamp 1649977179
transform 1 0 22356 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_246
timestamp 1649977179
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_253
timestamp 1649977179
transform 1 0 24380 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_259
timestamp 1649977179
transform 1 0 24932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_271
timestamp 1649977179
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_301
timestamp 1649977179
transform 1 0 28796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1649977179
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1649977179
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_69
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1649977179
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_103
timestamp 1649977179
transform 1 0 10580 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_147
timestamp 1649977179
transform 1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1649977179
transform 1 0 15272 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_160
timestamp 1649977179
transform 1 0 15824 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_166
timestamp 1649977179
transform 1 0 16376 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_178
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_183
timestamp 1649977179
transform 1 0 17940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_203
timestamp 1649977179
transform 1 0 19780 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_212
timestamp 1649977179
transform 1 0 20608 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_218
timestamp 1649977179
transform 1 0 21160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_226
timestamp 1649977179
transform 1 0 21896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_229
timestamp 1649977179
transform 1 0 22172 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_236
timestamp 1649977179
transform 1 0 22816 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1649977179
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_255
timestamp 1649977179
transform 1 0 24564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_267
timestamp 1649977179
transform 1 0 25668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_279
timestamp 1649977179
transform 1 0 26772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_291
timestamp 1649977179
transform 1 0 27876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_303
timestamp 1649977179
transform 1 0 28980 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_47
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_61
timestamp 1649977179
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_67
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_77
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_89
timestamp 1649977179
transform 1 0 9292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1649977179
transform 1 0 9844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_98
timestamp 1649977179
transform 1 0 10120 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_139
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_157
timestamp 1649977179
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1649977179
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_183
timestamp 1649977179
transform 1 0 17940 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1649977179
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_192
timestamp 1649977179
transform 1 0 18768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_198
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_204
timestamp 1649977179
transform 1 0 19872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1649977179
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_233
timestamp 1649977179
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_252
timestamp 1649977179
transform 1 0 24288 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_258
timestamp 1649977179
transform 1 0 24840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_270
timestamp 1649977179
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1649977179
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_301
timestamp 1649977179
transform 1 0 28796 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_5
timestamp 1649977179
transform 1 0 1564 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_17
timestamp 1649977179
transform 1 0 2668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1649977179
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_47
timestamp 1649977179
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_54
timestamp 1649977179
transform 1 0 6072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_61
timestamp 1649977179
transform 1 0 6716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_68
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_89
timestamp 1649977179
transform 1 0 9292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_101
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_104
timestamp 1649977179
transform 1 0 10672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_110
timestamp 1649977179
transform 1 0 11224 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1649977179
transform 1 0 11960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_129
timestamp 1649977179
transform 1 0 12972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_143
timestamp 1649977179
transform 1 0 14260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1649977179
transform 1 0 14812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_155
timestamp 1649977179
transform 1 0 15364 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1649977179
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1649977179
transform 1 0 16744 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_176
timestamp 1649977179
transform 1 0 17296 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1649977179
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_200
timestamp 1649977179
transform 1 0 19504 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_206
timestamp 1649977179
transform 1 0 20056 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_212
timestamp 1649977179
transform 1 0 20608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_227
timestamp 1649977179
transform 1 0 21988 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_235
timestamp 1649977179
transform 1 0 22724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1649977179
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_293
timestamp 1649977179
transform 1 0 28060 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_7
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_19
timestamp 1649977179
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_31
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_37
timestamp 1649977179
transform 1 0 4508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_40
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_61
timestamp 1649977179
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_68
timestamp 1649977179
transform 1 0 7360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_75
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_87
timestamp 1649977179
transform 1 0 9108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1649977179
transform 1 0 11960 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_127
timestamp 1649977179
transform 1 0 12788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_134
timestamp 1649977179
transform 1 0 13432 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1649977179
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_148
timestamp 1649977179
transform 1 0 14720 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_174
timestamp 1649977179
transform 1 0 17112 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1649977179
transform 1 0 17848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_190
timestamp 1649977179
transform 1 0 18584 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_197
timestamp 1649977179
transform 1 0 19228 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_203
timestamp 1649977179
transform 1 0 19780 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_212
timestamp 1649977179
transform 1 0 20608 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1649977179
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_230
timestamp 1649977179
transform 1 0 22264 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_236
timestamp 1649977179
transform 1 0 22816 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_242
timestamp 1649977179
transform 1 0 23368 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_252
timestamp 1649977179
transform 1 0 24288 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_256
timestamp 1649977179
transform 1 0 24656 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_259
timestamp 1649977179
transform 1 0 24932 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_267
timestamp 1649977179
transform 1 0 25668 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_270
timestamp 1649977179
transform 1 0 25944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1649977179
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_283
timestamp 1649977179
transform 1 0 27140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_289
timestamp 1649977179
transform 1 0 27692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_295
timestamp 1649977179
transform 1 0 28244 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_301
timestamp 1649977179
transform 1 0 28796 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_36
timestamp 1649977179
transform 1 0 4416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_45
timestamp 1649977179
transform 1 0 5244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_57
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_63
timestamp 1649977179
transform 1 0 6900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_67
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_73
timestamp 1649977179
transform 1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_94
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_106
timestamp 1649977179
transform 1 0 10856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_117
timestamp 1649977179
transform 1 0 11868 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_127
timestamp 1649977179
transform 1 0 12788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_134
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_146
timestamp 1649977179
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_152
timestamp 1649977179
transform 1 0 15088 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_156
timestamp 1649977179
transform 1 0 15456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_173
timestamp 1649977179
transform 1 0 17020 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_179
timestamp 1649977179
transform 1 0 17572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_205
timestamp 1649977179
transform 1 0 19964 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_214
timestamp 1649977179
transform 1 0 20792 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_220
timestamp 1649977179
transform 1 0 21344 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_226
timestamp 1649977179
transform 1 0 21896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1649977179
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_239
timestamp 1649977179
transform 1 0 23092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1649977179
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_255
timestamp 1649977179
transform 1 0 24564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_268
timestamp 1649977179
transform 1 0 25760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1649977179
transform 1 0 26496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_286
timestamp 1649977179
transform 1 0 27416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_299
timestamp 1649977179
transform 1 0 28612 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_60
timestamp 1649977179
transform 1 0 6624 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_70
timestamp 1649977179
transform 1 0 7544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1649977179
transform 1 0 8280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_89
timestamp 1649977179
transform 1 0 9292 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_96
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1649977179
transform 1 0 11868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_135
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_141
timestamp 1649977179
transform 1 0 14076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_147
timestamp 1649977179
transform 1 0 14628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_153
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_156
timestamp 1649977179
transform 1 0 15456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_182
timestamp 1649977179
transform 1 0 17848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_186
timestamp 1649977179
transform 1 0 18216 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_195
timestamp 1649977179
transform 1 0 19044 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_207
timestamp 1649977179
transform 1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_213
timestamp 1649977179
transform 1 0 20700 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1649977179
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_227
timestamp 1649977179
transform 1 0 21988 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_231
timestamp 1649977179
transform 1 0 22356 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_246
timestamp 1649977179
transform 1 0 23736 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_258
timestamp 1649977179
transform 1 0 24840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_266
timestamp 1649977179
transform 1 0 25576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_271
timestamp 1649977179
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_285
timestamp 1649977179
transform 1 0 27324 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_301
timestamp 1649977179
transform 1 0 28796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_5
timestamp 1649977179
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_14
timestamp 1649977179
transform 1 0 2392 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_22
timestamp 1649977179
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_37
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1649977179
transform 1 0 5336 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_56
timestamp 1649977179
transform 1 0 6256 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_68
timestamp 1649977179
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_92
timestamp 1649977179
transform 1 0 9568 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1649977179
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_111
timestamp 1649977179
transform 1 0 11316 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_117
timestamp 1649977179
transform 1 0 11868 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_125
timestamp 1649977179
transform 1 0 12604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp 1649977179
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_143
timestamp 1649977179
transform 1 0 14260 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_152
timestamp 1649977179
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1649977179
transform 1 0 16192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_176
timestamp 1649977179
transform 1 0 17296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_180
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_183
timestamp 1649977179
transform 1 0 17940 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1649977179
transform 1 0 19504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_206
timestamp 1649977179
transform 1 0 20056 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_212
timestamp 1649977179
transform 1 0 20608 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_220
timestamp 1649977179
transform 1 0 21344 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_239
timestamp 1649977179
transform 1 0 23092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_255
timestamp 1649977179
transform 1 0 24564 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_267
timestamp 1649977179
transform 1 0 25668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_279
timestamp 1649977179
transform 1 0 26772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_292
timestamp 1649977179
transform 1 0 27968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_296
timestamp 1649977179
transform 1 0 28336 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp 1649977179
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_20
timestamp 1649977179
transform 1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_26
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_45
timestamp 1649977179
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_59
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_67
timestamp 1649977179
transform 1 0 7268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1649977179
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1649977179
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_115
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_127
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_131
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1649977179
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_151
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 1649977179
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_186
timestamp 1649977179
transform 1 0 18216 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_198
timestamp 1649977179
transform 1 0 19320 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_213
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_234
timestamp 1649977179
transform 1 0 22632 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_240
timestamp 1649977179
transform 1 0 23184 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_246
timestamp 1649977179
transform 1 0 23736 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_258
timestamp 1649977179
transform 1 0 24840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_271
timestamp 1649977179
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_290
timestamp 1649977179
transform 1 0 27784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_302
timestamp 1649977179
transform 1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_16
timestamp 1649977179
transform 1 0 2576 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_31
timestamp 1649977179
transform 1 0 3956 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_42
timestamp 1649977179
transform 1 0 4968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_51
timestamp 1649977179
transform 1 0 5796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_57
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_60
timestamp 1649977179
transform 1 0 6624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_71
timestamp 1649977179
transform 1 0 7636 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_94
timestamp 1649977179
transform 1 0 9752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_100
timestamp 1649977179
transform 1 0 10304 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_122
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_130
timestamp 1649977179
transform 1 0 13064 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1649977179
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1649977179
transform 1 0 15272 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_160
timestamp 1649977179
transform 1 0 15824 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_174
timestamp 1649977179
transform 1 0 17112 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_183
timestamp 1649977179
transform 1 0 17940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_217
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_220
timestamp 1649977179
transform 1 0 21344 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_232
timestamp 1649977179
transform 1 0 22448 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_240
timestamp 1649977179
transform 1 0 23184 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_246
timestamp 1649977179
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_268
timestamp 1649977179
transform 1 0 25760 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_280
timestamp 1649977179
transform 1 0 26864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_285
timestamp 1649977179
transform 1 0 27324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_293
timestamp 1649977179
transform 1 0 28060 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_16
timestamp 1649977179
transform 1 0 2576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_25
timestamp 1649977179
transform 1 0 3404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_31
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_38
timestamp 1649977179
transform 1 0 4600 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1649977179
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_63
timestamp 1649977179
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_68
timestamp 1649977179
transform 1 0 7360 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_80
timestamp 1649977179
transform 1 0 8464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_91
timestamp 1649977179
transform 1 0 9476 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_115
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1649977179
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_135
timestamp 1649977179
transform 1 0 13524 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_143
timestamp 1649977179
transform 1 0 14260 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_146
timestamp 1649977179
transform 1 0 14536 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_155
timestamp 1649977179
transform 1 0 15364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_173
timestamp 1649977179
transform 1 0 17020 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_186
timestamp 1649977179
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_192
timestamp 1649977179
transform 1 0 18768 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_198
timestamp 1649977179
transform 1 0 19320 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_206
timestamp 1649977179
transform 1 0 20056 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_211
timestamp 1649977179
transform 1 0 20516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_227
timestamp 1649977179
transform 1 0 21988 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_233
timestamp 1649977179
transform 1 0 22540 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1649977179
transform 1 0 23092 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_248
timestamp 1649977179
transform 1 0 23920 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1649977179
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_258
timestamp 1649977179
transform 1 0 24840 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_267
timestamp 1649977179
transform 1 0 25668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_291
timestamp 1649977179
transform 1 0 27876 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_301
timestamp 1649977179
transform 1 0 28796 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_18
timestamp 1649977179
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1649977179
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_88
timestamp 1649977179
transform 1 0 9200 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_108
timestamp 1649977179
transform 1 0 11040 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_114
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1649977179
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_143
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_149
timestamp 1649977179
transform 1 0 14812 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_161
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_167
timestamp 1649977179
transform 1 0 16468 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_173
timestamp 1649977179
transform 1 0 17020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_186
timestamp 1649977179
transform 1 0 18216 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_199
timestamp 1649977179
transform 1 0 19412 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1649977179
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_216
timestamp 1649977179
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_226
timestamp 1649977179
transform 1 0 21896 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_235
timestamp 1649977179
transform 1 0 22724 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_239
timestamp 1649977179
transform 1 0 23092 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1649977179
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_266
timestamp 1649977179
transform 1 0 25576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_272
timestamp 1649977179
transform 1 0 26128 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_285
timestamp 1649977179
transform 1 0 27324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_298
timestamp 1649977179
transform 1 0 28520 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_304
timestamp 1649977179
transform 1 0 29072 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_7
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_13
timestamp 1649977179
transform 1 0 2300 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_16
timestamp 1649977179
transform 1 0 2576 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_28
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_43
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_59
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_71
timestamp 1649977179
transform 1 0 7636 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_95
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1649977179
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_115
timestamp 1649977179
transform 1 0 11684 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_123
timestamp 1649977179
transform 1 0 12420 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_128
timestamp 1649977179
transform 1 0 12880 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_141
timestamp 1649977179
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_147
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_178
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_189
timestamp 1649977179
transform 1 0 18492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_197
timestamp 1649977179
transform 1 0 19228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_207
timestamp 1649977179
transform 1 0 20148 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_211
timestamp 1649977179
transform 1 0 20516 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_229
timestamp 1649977179
transform 1 0 22172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_236
timestamp 1649977179
transform 1 0 22816 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_246
timestamp 1649977179
transform 1 0 23736 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_253
timestamp 1649977179
transform 1 0 24380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_257
timestamp 1649977179
transform 1 0 24748 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_267
timestamp 1649977179
transform 1 0 25668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_284
timestamp 1649977179
transform 1 0 27232 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_292
timestamp 1649977179
transform 1 0 27968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_304
timestamp 1649977179
transform 1 0 29072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_14
timestamp 1649977179
transform 1 0 2392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1649977179
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp 1649977179
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_39
timestamp 1649977179
transform 1 0 4692 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_51
timestamp 1649977179
transform 1 0 5796 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_63
timestamp 1649977179
transform 1 0 6900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1649977179
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1649977179
transform 1 0 9200 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_94
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1649977179
transform 1 0 10488 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_108
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_114
timestamp 1649977179
transform 1 0 11592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_117
timestamp 1649977179
transform 1 0 11868 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_125
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_148
timestamp 1649977179
transform 1 0 14720 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_160
timestamp 1649977179
transform 1 0 15824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1649977179
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1649977179
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_203
timestamp 1649977179
transform 1 0 19780 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1649977179
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_227
timestamp 1649977179
transform 1 0 21988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_235
timestamp 1649977179
transform 1 0 22724 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_241
timestamp 1649977179
transform 1 0 23276 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1649977179
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_255
timestamp 1649977179
transform 1 0 24564 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_267
timestamp 1649977179
transform 1 0 25668 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_279
timestamp 1649977179
transform 1 0 26772 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_291
timestamp 1649977179
transform 1 0 27876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_303
timestamp 1649977179
transform 1 0 28980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1649977179
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1649977179
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_35
timestamp 1649977179
transform 1 0 4324 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 1649977179
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_59
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_70
timestamp 1649977179
transform 1 0 7544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_76
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_90
timestamp 1649977179
transform 1 0 9384 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_96
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_102
timestamp 1649977179
transform 1 0 10488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_118
timestamp 1649977179
transform 1 0 11960 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_124
timestamp 1649977179
transform 1 0 12512 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_133
timestamp 1649977179
transform 1 0 13340 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_139
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_147
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_180
timestamp 1649977179
transform 1 0 17664 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1649977179
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_207
timestamp 1649977179
transform 1 0 20148 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1649977179
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_233
timestamp 1649977179
transform 1 0 22540 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1649977179
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_250
timestamp 1649977179
transform 1 0 24104 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_299
timestamp 1649977179
transform 1 0 28612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_16
timestamp 1649977179
transform 1 0 2576 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_39
timestamp 1649977179
transform 1 0 4692 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_47
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_55
timestamp 1649977179
transform 1 0 6164 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_61
timestamp 1649977179
transform 1 0 6716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp 1649977179
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1649977179
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_91
timestamp 1649977179
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_103
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_107
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1649977179
transform 1 0 11684 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_132
timestamp 1649977179
transform 1 0 13248 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_145
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_156
timestamp 1649977179
transform 1 0 15456 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_170
timestamp 1649977179
transform 1 0 16744 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_178
timestamp 1649977179
transform 1 0 17480 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_183
timestamp 1649977179
transform 1 0 17940 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1649977179
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_208
timestamp 1649977179
transform 1 0 20240 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_216
timestamp 1649977179
transform 1 0 20976 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_220
timestamp 1649977179
transform 1 0 21344 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_232
timestamp 1649977179
transform 1 0 22448 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_244
timestamp 1649977179
transform 1 0 23552 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_257
timestamp 1649977179
transform 1 0 24748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_267
timestamp 1649977179
transform 1 0 25668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_273
timestamp 1649977179
transform 1 0 26220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_281
timestamp 1649977179
transform 1 0 26956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_294
timestamp 1649977179
transform 1 0 28152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_300
timestamp 1649977179
transform 1 0 28704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_304
timestamp 1649977179
transform 1 0 29072 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_47
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1649977179
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_59
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_70
timestamp 1649977179
transform 1 0 7544 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_74
timestamp 1649977179
transform 1 0 7912 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_87
timestamp 1649977179
transform 1 0 9108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_95
timestamp 1649977179
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_99
timestamp 1649977179
transform 1 0 10212 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1649977179
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_119
timestamp 1649977179
transform 1 0 12052 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_127
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1649977179
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_145
timestamp 1649977179
transform 1 0 14444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_153
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1649977179
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_173
timestamp 1649977179
transform 1 0 17020 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1649977179
transform 1 0 17572 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 1649977179
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_202
timestamp 1649977179
transform 1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1649977179
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_212
timestamp 1649977179
transform 1 0 20608 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1649977179
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_244
timestamp 1649977179
transform 1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_251
timestamp 1649977179
transform 1 0 24196 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_265
timestamp 1649977179
transform 1 0 25484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1649977179
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_301
timestamp 1649977179
transform 1 0 28796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_7
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_13
timestamp 1649977179
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1649977179
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_71
timestamp 1649977179
transform 1 0 7636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1649977179
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1649977179
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1649977179
transform 1 0 9752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_98
timestamp 1649977179
transform 1 0 10120 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_101
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_113
timestamp 1649977179
transform 1 0 11500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_128
timestamp 1649977179
transform 1 0 12880 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_161
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_173
timestamp 1649977179
transform 1 0 17020 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_185
timestamp 1649977179
transform 1 0 18124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1649977179
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_199
timestamp 1649977179
transform 1 0 19412 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_215
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_222
timestamp 1649977179
transform 1 0 21528 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_234
timestamp 1649977179
transform 1 0 22632 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_242
timestamp 1649977179
transform 1 0 23368 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1649977179
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_256
timestamp 1649977179
transform 1 0 24656 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_262
timestamp 1649977179
transform 1 0 25208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_269
timestamp 1649977179
transform 1 0 25852 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_278
timestamp 1649977179
transform 1 0 26680 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_286
timestamp 1649977179
transform 1 0 27416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_291
timestamp 1649977179
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_297
timestamp 1649977179
transform 1 0 28428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_14
timestamp 1649977179
transform 1 0 2392 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_26
timestamp 1649977179
transform 1 0 3496 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_29
timestamp 1649977179
transform 1 0 3772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_36
timestamp 1649977179
transform 1 0 4416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_42
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_46
timestamp 1649977179
transform 1 0 5336 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1649977179
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1649977179
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_65
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_71
timestamp 1649977179
transform 1 0 7636 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_83
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_89
timestamp 1649977179
transform 1 0 9292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_115
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_121
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_127
timestamp 1649977179
transform 1 0 12788 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_139
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_151
timestamp 1649977179
transform 1 0 14996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_155
timestamp 1649977179
transform 1 0 15364 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1649977179
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_216
timestamp 1649977179
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_240
timestamp 1649977179
transform 1 0 23184 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_248
timestamp 1649977179
transform 1 0 23920 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_259
timestamp 1649977179
transform 1 0 24932 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_271
timestamp 1649977179
transform 1 0 26036 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_285
timestamp 1649977179
transform 1 0 27324 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_290
timestamp 1649977179
transform 1 0 27784 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_296
timestamp 1649977179
transform 1 0 28336 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_301
timestamp 1649977179
transform 1 0 28796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1649977179
transform 1 0 2392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1649977179
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_39
timestamp 1649977179
transform 1 0 4692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_47
timestamp 1649977179
transform 1 0 5428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_60
timestamp 1649977179
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_64
timestamp 1649977179
transform 1 0 6992 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_71
timestamp 1649977179
transform 1 0 7636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_92
timestamp 1649977179
transform 1 0 9568 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_105
timestamp 1649977179
transform 1 0 10764 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1649977179
transform 1 0 11684 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_148
timestamp 1649977179
transform 1 0 14720 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_178
timestamp 1649977179
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_205
timestamp 1649977179
transform 1 0 19964 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_216
timestamp 1649977179
transform 1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_225
timestamp 1649977179
transform 1 0 21804 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_237
timestamp 1649977179
transform 1 0 22908 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_241
timestamp 1649977179
transform 1 0 23276 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1649977179
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_261
timestamp 1649977179
transform 1 0 25116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_273
timestamp 1649977179
transform 1 0 26220 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_276
timestamp 1649977179
transform 1 0 26496 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_282
timestamp 1649977179
transform 1 0 27048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_295
timestamp 1649977179
transform 1 0 28244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1649977179
transform 1 0 3864 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_48
timestamp 1649977179
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_65
timestamp 1649977179
transform 1 0 7084 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_75
timestamp 1649977179
transform 1 0 8004 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_89
timestamp 1649977179
transform 1 0 9292 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_100
timestamp 1649977179
transform 1 0 10304 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1649977179
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_119
timestamp 1649977179
transform 1 0 12052 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1649977179
transform 1 0 13156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_147
timestamp 1649977179
transform 1 0 14628 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_153
timestamp 1649977179
transform 1 0 15180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1649977179
transform 1 0 17572 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1649977179
transform 1 0 18400 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_194
timestamp 1649977179
transform 1 0 18952 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_202
timestamp 1649977179
transform 1 0 19688 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_207
timestamp 1649977179
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1649977179
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_259
timestamp 1649977179
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_271
timestamp 1649977179
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_290
timestamp 1649977179
transform 1 0 27784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_298
timestamp 1649977179
transform 1 0 28520 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_304
timestamp 1649977179
transform 1 0 29072 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_35
timestamp 1649977179
transform 1 0 4324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_47
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_50
timestamp 1649977179
transform 1 0 5704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_54
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_100
timestamp 1649977179
transform 1 0 10304 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_106
timestamp 1649977179
transform 1 0 10856 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_112
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_118
timestamp 1649977179
transform 1 0 11960 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_149
timestamp 1649977179
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_159
timestamp 1649977179
transform 1 0 15732 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_175
timestamp 1649977179
transform 1 0 17204 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_181
timestamp 1649977179
transform 1 0 17756 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_187
timestamp 1649977179
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_199
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_207
timestamp 1649977179
transform 1 0 20148 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_211
timestamp 1649977179
transform 1 0 20516 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_223
timestamp 1649977179
transform 1 0 21620 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_241
timestamp 1649977179
transform 1 0 23276 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1649977179
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_271
timestamp 1649977179
transform 1 0 26036 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1649977179
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1649977179
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_12
timestamp 1649977179
transform 1 0 2208 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_24
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_28
timestamp 1649977179
transform 1 0 3680 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1649977179
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1649977179
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_73
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_79
timestamp 1649977179
transform 1 0 8372 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_89
timestamp 1649977179
transform 1 0 9292 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_95
timestamp 1649977179
transform 1 0 9844 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_98
timestamp 1649977179
transform 1 0 10120 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1649977179
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_120
timestamp 1649977179
transform 1 0 12144 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_126
timestamp 1649977179
transform 1 0 12696 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_131
timestamp 1649977179
transform 1 0 13156 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_140
timestamp 1649977179
transform 1 0 13984 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_146
timestamp 1649977179
transform 1 0 14536 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_156
timestamp 1649977179
transform 1 0 15456 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_178
timestamp 1649977179
transform 1 0 17480 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_184
timestamp 1649977179
transform 1 0 18032 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1649977179
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_200
timestamp 1649977179
transform 1 0 19504 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_206
timestamp 1649977179
transform 1 0 20056 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_216
timestamp 1649977179
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_227
timestamp 1649977179
transform 1 0 21988 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_238
timestamp 1649977179
transform 1 0 23000 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_244
timestamp 1649977179
transform 1 0 23552 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_259
timestamp 1649977179
transform 1 0 24932 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_271
timestamp 1649977179
transform 1 0 26036 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_290
timestamp 1649977179
transform 1 0 27784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_298
timestamp 1649977179
transform 1 0 28520 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_304
timestamp 1649977179
transform 1 0 29072 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_14
timestamp 1649977179
transform 1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_20
timestamp 1649977179
transform 1 0 2944 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_45
timestamp 1649977179
transform 1 0 5244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_57
timestamp 1649977179
transform 1 0 6348 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1649977179
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_72
timestamp 1649977179
transform 1 0 7728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1649977179
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_96
timestamp 1649977179
transform 1 0 9936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_102
timestamp 1649977179
transform 1 0 10488 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_110
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_119
timestamp 1649977179
transform 1 0 12052 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_131
timestamp 1649977179
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_152
timestamp 1649977179
transform 1 0 15088 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_164
timestamp 1649977179
transform 1 0 16192 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1649977179
transform 1 0 17296 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1649977179
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_186
timestamp 1649977179
transform 1 0 18216 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_201
timestamp 1649977179
transform 1 0 19596 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_207
timestamp 1649977179
transform 1 0 20148 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_227
timestamp 1649977179
transform 1 0 21988 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1649977179
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_266
timestamp 1649977179
transform 1 0 25576 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1649977179
transform 1 0 26312 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_284
timestamp 1649977179
transform 1 0 27232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_292
timestamp 1649977179
transform 1 0 27968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_296
timestamp 1649977179
transform 1 0 28336 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_14
timestamp 1649977179
transform 1 0 2392 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_26
timestamp 1649977179
transform 1 0 3496 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_38
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_41
timestamp 1649977179
transform 1 0 4876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_49
timestamp 1649977179
transform 1 0 5612 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_59
timestamp 1649977179
transform 1 0 6532 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_63
timestamp 1649977179
transform 1 0 6900 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_66
timestamp 1649977179
transform 1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_73
timestamp 1649977179
transform 1 0 7820 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_87
timestamp 1649977179
transform 1 0 9108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_98
timestamp 1649977179
transform 1 0 10120 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_104
timestamp 1649977179
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_122
timestamp 1649977179
transform 1 0 12328 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_130
timestamp 1649977179
transform 1 0 13064 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_171
timestamp 1649977179
transform 1 0 16836 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_183
timestamp 1649977179
transform 1 0 17940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_195
timestamp 1649977179
transform 1 0 19044 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_210
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_231
timestamp 1649977179
transform 1 0 22356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_235
timestamp 1649977179
transform 1 0 22724 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_243
timestamp 1649977179
transform 1 0 23460 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_255
timestamp 1649977179
transform 1 0 24564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_267
timestamp 1649977179
transform 1 0 25668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_286
timestamp 1649977179
transform 1 0 27416 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_294
timestamp 1649977179
transform 1 0 28152 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_297
timestamp 1649977179
transform 1 0 28428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_43
timestamp 1649977179
transform 1 0 5060 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_60
timestamp 1649977179
transform 1 0 6624 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_71
timestamp 1649977179
transform 1 0 7636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1649977179
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_115
timestamp 1649977179
transform 1 0 11684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_127
timestamp 1649977179
transform 1 0 12788 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_135
timestamp 1649977179
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_146
timestamp 1649977179
transform 1 0 14536 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_154
timestamp 1649977179
transform 1 0 15272 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_158
timestamp 1649977179
transform 1 0 15640 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_178
timestamp 1649977179
transform 1 0 17480 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_184
timestamp 1649977179
transform 1 0 18032 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_226
timestamp 1649977179
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_232
timestamp 1649977179
transform 1 0 22448 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_244
timestamp 1649977179
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_260
timestamp 1649977179
transform 1 0 25024 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_266
timestamp 1649977179
transform 1 0 25576 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_276
timestamp 1649977179
transform 1 0 26496 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_282
timestamp 1649977179
transform 1 0 27048 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_295
timestamp 1649977179
transform 1 0 28244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_13
timestamp 1649977179
transform 1 0 2300 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_25
timestamp 1649977179
transform 1 0 3404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_29
timestamp 1649977179
transform 1 0 3772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_37
timestamp 1649977179
transform 1 0 4508 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1649977179
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_64
timestamp 1649977179
transform 1 0 6992 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_70
timestamp 1649977179
transform 1 0 7544 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_74
timestamp 1649977179
transform 1 0 7912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_80
timestamp 1649977179
transform 1 0 8464 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_86
timestamp 1649977179
transform 1 0 9016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_89
timestamp 1649977179
transform 1 0 9292 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_97
timestamp 1649977179
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_103
timestamp 1649977179
transform 1 0 10580 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_121
timestamp 1649977179
transform 1 0 12236 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_133
timestamp 1649977179
transform 1 0 13340 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_141
timestamp 1649977179
transform 1 0 14076 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_152
timestamp 1649977179
transform 1 0 15088 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1649977179
transform 1 0 15824 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_176
timestamp 1649977179
transform 1 0 17296 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_182
timestamp 1649977179
transform 1 0 17848 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_188
timestamp 1649977179
transform 1 0 18400 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_200
timestamp 1649977179
transform 1 0 19504 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_204
timestamp 1649977179
transform 1 0 19872 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_207
timestamp 1649977179
transform 1 0 20148 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1649977179
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_248
timestamp 1649977179
transform 1 0 23920 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_260
timestamp 1649977179
transform 1 0 25024 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1649977179
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_285
timestamp 1649977179
transform 1 0 27324 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_296
timestamp 1649977179
transform 1 0 28336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_304
timestamp 1649977179
transform 1 0 29072 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_8
timestamp 1649977179
transform 1 0 1840 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_16
timestamp 1649977179
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_37
timestamp 1649977179
transform 1 0 4508 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp 1649977179
transform 1 0 4784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_46
timestamp 1649977179
transform 1 0 5336 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_57
timestamp 1649977179
transform 1 0 6348 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_68
timestamp 1649977179
transform 1 0 7360 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_74
timestamp 1649977179
transform 1 0 7912 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1649977179
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_92
timestamp 1649977179
transform 1 0 9568 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_98
timestamp 1649977179
transform 1 0 10120 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_101
timestamp 1649977179
transform 1 0 10396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_113
timestamp 1649977179
transform 1 0 11500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_125
timestamp 1649977179
transform 1 0 12604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1649977179
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_144
timestamp 1649977179
transform 1 0 14352 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_178
timestamp 1649977179
transform 1 0 17480 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1649977179
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_205
timestamp 1649977179
transform 1 0 19964 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1649977179
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_226
timestamp 1649977179
transform 1 0 21896 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_238
timestamp 1649977179
transform 1 0 23000 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1649977179
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_256
timestamp 1649977179
transform 1 0 24656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_268
timestamp 1649977179
transform 1 0 25760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_281
timestamp 1649977179
transform 1 0 26956 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_294
timestamp 1649977179
transform 1 0 28152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1649977179
transform 1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_25
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_29
timestamp 1649977179
transform 1 0 3772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_34
timestamp 1649977179
transform 1 0 4232 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_40
timestamp 1649977179
transform 1 0 4784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_46
timestamp 1649977179
transform 1 0 5336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1649977179
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_65
timestamp 1649977179
transform 1 0 7084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_71
timestamp 1649977179
transform 1 0 7636 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1649977179
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_88
timestamp 1649977179
transform 1 0 9200 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_100
timestamp 1649977179
transform 1 0 10304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1649977179
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_133
timestamp 1649977179
transform 1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_141
timestamp 1649977179
transform 1 0 14076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_153
timestamp 1649977179
transform 1 0 15180 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1649977179
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1649977179
transform 1 0 16928 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1649977179
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_184
timestamp 1649977179
transform 1 0 18032 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_196
timestamp 1649977179
transform 1 0 19136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_200
timestamp 1649977179
transform 1 0 19504 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_213
timestamp 1649977179
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1649977179
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_244
timestamp 1649977179
transform 1 0 23552 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1649977179
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_285
timestamp 1649977179
transform 1 0 27324 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_295
timestamp 1649977179
transform 1 0 28244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_301
timestamp 1649977179
transform 1 0 28796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_14
timestamp 1649977179
transform 1 0 2392 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1649977179
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_38
timestamp 1649977179
transform 1 0 4600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_48
timestamp 1649977179
transform 1 0 5520 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_59
timestamp 1649977179
transform 1 0 6532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_69
timestamp 1649977179
transform 1 0 7452 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1649977179
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_89
timestamp 1649977179
transform 1 0 9292 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1649977179
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_108
timestamp 1649977179
transform 1 0 11040 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1649977179
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_120
timestamp 1649977179
transform 1 0 12144 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_126
timestamp 1649977179
transform 1 0 12696 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_148
timestamp 1649977179
transform 1 0 14720 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1649977179
transform 1 0 15640 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_164
timestamp 1649977179
transform 1 0 16192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_199
timestamp 1649977179
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_227
timestamp 1649977179
transform 1 0 21988 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_237
timestamp 1649977179
transform 1 0 22908 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1649977179
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_275
timestamp 1649977179
transform 1 0 26404 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_283
timestamp 1649977179
transform 1 0 27140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_286
timestamp 1649977179
transform 1 0 27416 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_296
timestamp 1649977179
transform 1 0 28336 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_304
timestamp 1649977179
transform 1 0 29072 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_11
timestamp 1649977179
transform 1 0 2116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_17
timestamp 1649977179
transform 1 0 2668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_21
timestamp 1649977179
transform 1 0 3036 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_30
timestamp 1649977179
transform 1 0 3864 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_36
timestamp 1649977179
transform 1 0 4416 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_40
timestamp 1649977179
transform 1 0 4784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_48
timestamp 1649977179
transform 1 0 5520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1649977179
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_59
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1649977179
transform 1 0 7636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_77
timestamp 1649977179
transform 1 0 8188 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1649977179
transform 1 0 9016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_90
timestamp 1649977179
transform 1 0 9384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_98
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_104
timestamp 1649977179
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_117
timestamp 1649977179
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_120
timestamp 1649977179
transform 1 0 12144 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_124
timestamp 1649977179
transform 1 0 12512 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_131
timestamp 1649977179
transform 1 0 13156 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_146
timestamp 1649977179
transform 1 0 14536 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_158
timestamp 1649977179
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1649977179
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_171
timestamp 1649977179
transform 1 0 16836 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_185
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_207
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_227
timestamp 1649977179
transform 1 0 21988 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_235
timestamp 1649977179
transform 1 0 22724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1649977179
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_244
timestamp 1649977179
transform 1 0 23552 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_247
timestamp 1649977179
transform 1 0 23828 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_256
timestamp 1649977179
transform 1 0 24656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_269
timestamp 1649977179
transform 1 0 25852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1649977179
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_283
timestamp 1649977179
transform 1 0 27140 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_291
timestamp 1649977179
transform 1 0 27876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_297
timestamp 1649977179
transform 1 0 28428 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_61
timestamp 1649977179
transform 1 0 6716 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_69
timestamp 1649977179
transform 1 0 7452 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_74
timestamp 1649977179
transform 1 0 7912 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1649977179
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_96
timestamp 1649977179
transform 1 0 9936 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_108
timestamp 1649977179
transform 1 0 11040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_118
timestamp 1649977179
transform 1 0 11960 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_122
timestamp 1649977179
transform 1 0 12328 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_126
timestamp 1649977179
transform 1 0 12696 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1649977179
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_149
timestamp 1649977179
transform 1 0 14812 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_161
timestamp 1649977179
transform 1 0 15916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_169
timestamp 1649977179
transform 1 0 16652 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_173
timestamp 1649977179
transform 1 0 17020 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_183
timestamp 1649977179
transform 1 0 17940 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1649977179
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_199
timestamp 1649977179
transform 1 0 19412 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_211
timestamp 1649977179
transform 1 0 20516 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_216
timestamp 1649977179
transform 1 0 20976 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_222
timestamp 1649977179
transform 1 0 21528 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_229
timestamp 1649977179
transform 1 0 22172 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_235
timestamp 1649977179
transform 1 0 22724 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_241
timestamp 1649977179
transform 1 0 23276 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_258
timestamp 1649977179
transform 1 0 24840 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_264
timestamp 1649977179
transform 1 0 25392 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_267
timestamp 1649977179
transform 1 0 25668 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_275
timestamp 1649977179
transform 1 0 26404 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_300
timestamp 1649977179
transform 1 0 28704 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_304
timestamp 1649977179
transform 1 0 29072 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_11
timestamp 1649977179
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_16
timestamp 1649977179
transform 1 0 2576 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_22
timestamp 1649977179
transform 1 0 3128 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_30
timestamp 1649977179
transform 1 0 3864 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_84
timestamp 1649977179
transform 1 0 8832 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_96
timestamp 1649977179
transform 1 0 9936 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_102
timestamp 1649977179
transform 1 0 10488 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1649977179
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_115
timestamp 1649977179
transform 1 0 11684 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_123
timestamp 1649977179
transform 1 0 12420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_128
timestamp 1649977179
transform 1 0 12880 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_135
timestamp 1649977179
transform 1 0 13524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_148
timestamp 1649977179
transform 1 0 14720 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_160
timestamp 1649977179
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1649977179
transform 1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_191
timestamp 1649977179
transform 1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_197
timestamp 1649977179
transform 1 0 19228 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_203
timestamp 1649977179
transform 1 0 19780 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1649977179
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_213
timestamp 1649977179
transform 1 0 20700 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_227
timestamp 1649977179
transform 1 0 21988 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_231
timestamp 1649977179
transform 1 0 22356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_245
timestamp 1649977179
transform 1 0 23644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_253
timestamp 1649977179
transform 1 0 24380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_267
timestamp 1649977179
transform 1 0 25668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_290
timestamp 1649977179
transform 1 0 27784 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_296
timestamp 1649977179
transform 1 0 28336 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1649977179
transform 1 0 28796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_14
timestamp 1649977179
transform 1 0 2392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1649977179
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_32
timestamp 1649977179
transform 1 0 4048 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_44
timestamp 1649977179
transform 1 0 5152 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_56
timestamp 1649977179
transform 1 0 6256 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_60
timestamp 1649977179
transform 1 0 6624 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_63
timestamp 1649977179
transform 1 0 6900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_70
timestamp 1649977179
transform 1 0 7544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_76
timestamp 1649977179
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_89
timestamp 1649977179
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1649977179
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_105
timestamp 1649977179
transform 1 0 10764 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_111
timestamp 1649977179
transform 1 0 11316 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1649977179
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_129
timestamp 1649977179
transform 1 0 12972 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_132
timestamp 1649977179
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_151
timestamp 1649977179
transform 1 0 14996 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_163
timestamp 1649977179
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_175
timestamp 1649977179
transform 1 0 17204 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_179
timestamp 1649977179
transform 1 0 17572 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1649977179
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_206
timestamp 1649977179
transform 1 0 20056 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_210
timestamp 1649977179
transform 1 0 20424 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_232
timestamp 1649977179
transform 1 0 22448 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_255
timestamp 1649977179
transform 1 0 24564 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_267
timestamp 1649977179
transform 1 0 25668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_273
timestamp 1649977179
transform 1 0 26220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_279
timestamp 1649977179
transform 1 0 26772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_296
timestamp 1649977179
transform 1 0 28336 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_304
timestamp 1649977179
transform 1 0 29072 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_8
timestamp 1649977179
transform 1 0 1840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_25
timestamp 1649977179
transform 1 0 3404 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_35
timestamp 1649977179
transform 1 0 4324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_47
timestamp 1649977179
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_64
timestamp 1649977179
transform 1 0 6992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_71
timestamp 1649977179
transform 1 0 7636 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_79
timestamp 1649977179
transform 1 0 8372 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_85
timestamp 1649977179
transform 1 0 8924 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_91
timestamp 1649977179
transform 1 0 9476 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_94
timestamp 1649977179
transform 1 0 9752 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_100
timestamp 1649977179
transform 1 0 10304 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_106
timestamp 1649977179
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_123
timestamp 1649977179
transform 1 0 12420 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_131
timestamp 1649977179
transform 1 0 13156 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_143
timestamp 1649977179
transform 1 0 14260 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_154
timestamp 1649977179
transform 1 0 15272 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1649977179
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_174
timestamp 1649977179
transform 1 0 17112 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_180
timestamp 1649977179
transform 1 0 17664 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_183
timestamp 1649977179
transform 1 0 17940 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_199
timestamp 1649977179
transform 1 0 19412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_208
timestamp 1649977179
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_214
timestamp 1649977179
transform 1 0 20792 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1649977179
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_229
timestamp 1649977179
transform 1 0 22172 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_240
timestamp 1649977179
transform 1 0 23184 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_246
timestamp 1649977179
transform 1 0 23736 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_252
timestamp 1649977179
transform 1 0 24288 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_258
timestamp 1649977179
transform 1 0 24840 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_267
timestamp 1649977179
transform 1 0 25668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_283
timestamp 1649977179
transform 1 0 27140 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_297
timestamp 1649977179
transform 1 0 28428 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_5
timestamp 1649977179
transform 1 0 1564 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_17
timestamp 1649977179
transform 1 0 2668 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1649977179
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_40
timestamp 1649977179
transform 1 0 4784 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_48
timestamp 1649977179
transform 1 0 5520 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_51
timestamp 1649977179
transform 1 0 5796 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_59
timestamp 1649977179
transform 1 0 6532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_90
timestamp 1649977179
transform 1 0 9384 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_100
timestamp 1649977179
transform 1 0 10304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_112
timestamp 1649977179
transform 1 0 11408 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_126
timestamp 1649977179
transform 1 0 12696 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_134
timestamp 1649977179
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_145
timestamp 1649977179
transform 1 0 14444 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_161
timestamp 1649977179
transform 1 0 15916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_174
timestamp 1649977179
transform 1 0 17112 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1649977179
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_205
timestamp 1649977179
transform 1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_219
timestamp 1649977179
transform 1 0 21252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_231
timestamp 1649977179
transform 1 0 22356 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_237
timestamp 1649977179
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_243
timestamp 1649977179
transform 1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_266
timestamp 1649977179
transform 1 0 25576 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_272
timestamp 1649977179
transform 1 0 26128 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_33
timestamp 1649977179
transform 1 0 4140 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_40
timestamp 1649977179
transform 1 0 4784 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1649977179
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_63
timestamp 1649977179
transform 1 0 6900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_74
timestamp 1649977179
transform 1 0 7912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_78
timestamp 1649977179
transform 1 0 8280 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_88
timestamp 1649977179
transform 1 0 9200 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_100
timestamp 1649977179
transform 1 0 10304 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_106
timestamp 1649977179
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_115
timestamp 1649977179
transform 1 0 11684 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_121
timestamp 1649977179
transform 1 0 12236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_130
timestamp 1649977179
transform 1 0 13064 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_139
timestamp 1649977179
transform 1 0 13892 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1649977179
transform 1 0 15272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_160
timestamp 1649977179
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_177
timestamp 1649977179
transform 1 0 17388 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_189
timestamp 1649977179
transform 1 0 18492 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_199
timestamp 1649977179
transform 1 0 19412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_211
timestamp 1649977179
transform 1 0 20516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_227
timestamp 1649977179
transform 1 0 21988 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_231
timestamp 1649977179
transform 1 0 22356 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_238
timestamp 1649977179
transform 1 0 23000 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_244
timestamp 1649977179
transform 1 0 23552 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_250
timestamp 1649977179
transform 1 0 24104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_254
timestamp 1649977179
transform 1 0 24472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_263
timestamp 1649977179
transform 1 0 25300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_271
timestamp 1649977179
transform 1 0 26036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_283
timestamp 1649977179
transform 1 0 27140 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_289
timestamp 1649977179
transform 1 0 27692 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_292
timestamp 1649977179
transform 1 0 27968 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_296
timestamp 1649977179
transform 1 0 28336 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_301
timestamp 1649977179
transform 1 0 28796 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_5
timestamp 1649977179
transform 1 0 1564 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_17
timestamp 1649977179
transform 1 0 2668 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1649977179
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_33
timestamp 1649977179
transform 1 0 4140 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_37
timestamp 1649977179
transform 1 0 4508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_44
timestamp 1649977179
transform 1 0 5152 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_51
timestamp 1649977179
transform 1 0 5796 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_69
timestamp 1649977179
transform 1 0 7452 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_72
timestamp 1649977179
transform 1 0 7728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_78
timestamp 1649977179
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_92
timestamp 1649977179
transform 1 0 9568 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_104
timestamp 1649977179
transform 1 0 10672 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_110
timestamp 1649977179
transform 1 0 11224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_119
timestamp 1649977179
transform 1 0 12052 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_125
timestamp 1649977179
transform 1 0 12604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_137
timestamp 1649977179
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_151
timestamp 1649977179
transform 1 0 14996 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_163
timestamp 1649977179
transform 1 0 16100 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_175
timestamp 1649977179
transform 1 0 17204 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_187
timestamp 1649977179
transform 1 0 18308 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1649977179
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_207
timestamp 1649977179
transform 1 0 20148 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_213
timestamp 1649977179
transform 1 0 20700 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_219
timestamp 1649977179
transform 1 0 21252 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_223
timestamp 1649977179
transform 1 0 21620 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_229
timestamp 1649977179
transform 1 0 22172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_241
timestamp 1649977179
transform 1 0 23276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1649977179
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_257
timestamp 1649977179
transform 1 0 24748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_266
timestamp 1649977179
transform 1 0 25576 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_274
timestamp 1649977179
transform 1 0 26312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_280
timestamp 1649977179
transform 1 0 26864 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_286
timestamp 1649977179
transform 1 0 27416 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1649977179
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_298
timestamp 1649977179
transform 1 0 28520 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_7
timestamp 1649977179
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_19
timestamp 1649977179
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_31
timestamp 1649977179
transform 1 0 3956 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_42
timestamp 1649977179
transform 1 0 4968 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1649977179
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_71
timestamp 1649977179
transform 1 0 7636 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_78
timestamp 1649977179
transform 1 0 8280 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_86
timestamp 1649977179
transform 1 0 9016 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_90
timestamp 1649977179
transform 1 0 9384 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_98
timestamp 1649977179
transform 1 0 10120 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_102
timestamp 1649977179
transform 1 0 10488 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1649977179
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_121
timestamp 1649977179
transform 1 0 12236 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_135
timestamp 1649977179
transform 1 0 13524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_142
timestamp 1649977179
transform 1 0 14168 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_148
timestamp 1649977179
transform 1 0 14720 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_151
timestamp 1649977179
transform 1 0 14996 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_163
timestamp 1649977179
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_189
timestamp 1649977179
transform 1 0 18492 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_194
timestamp 1649977179
transform 1 0 18952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_198
timestamp 1649977179
transform 1 0 19320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_201
timestamp 1649977179
transform 1 0 19596 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_207
timestamp 1649977179
transform 1 0 20148 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_219
timestamp 1649977179
transform 1 0 21252 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_227
timestamp 1649977179
transform 1 0 21988 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_231
timestamp 1649977179
transform 1 0 22356 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_243
timestamp 1649977179
transform 1 0 23460 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_251
timestamp 1649977179
transform 1 0 24196 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_254
timestamp 1649977179
transform 1 0 24472 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_270
timestamp 1649977179
transform 1 0 25944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1649977179
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_283
timestamp 1649977179
transform 1 0 27140 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_289
timestamp 1649977179
transform 1 0 27692 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_295
timestamp 1649977179
transform 1 0 28244 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_298
timestamp 1649977179
transform 1 0 28520 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_304
timestamp 1649977179
transform 1 0 29072 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_39
timestamp 1649977179
transform 1 0 4692 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_46
timestamp 1649977179
transform 1 0 5336 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_58
timestamp 1649977179
transform 1 0 6440 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_64
timestamp 1649977179
transform 1 0 6992 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_69
timestamp 1649977179
transform 1 0 7452 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1649977179
transform 1 0 8280 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_88
timestamp 1649977179
transform 1 0 9200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_94
timestamp 1649977179
transform 1 0 9752 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_106
timestamp 1649977179
transform 1 0 10856 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_112
timestamp 1649977179
transform 1 0 11408 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_122
timestamp 1649977179
transform 1 0 12328 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_128
timestamp 1649977179
transform 1 0 12880 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1649977179
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_143
timestamp 1649977179
transform 1 0 14260 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_151
timestamp 1649977179
transform 1 0 14996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_160
timestamp 1649977179
transform 1 0 15824 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_166
timestamp 1649977179
transform 1 0 16376 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_172
timestamp 1649977179
transform 1 0 16928 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_178
timestamp 1649977179
transform 1 0 17480 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_184
timestamp 1649977179
transform 1 0 18032 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1649977179
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_203
timestamp 1649977179
transform 1 0 19780 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_215
timestamp 1649977179
transform 1 0 20884 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_225
timestamp 1649977179
transform 1 0 21804 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_229
timestamp 1649977179
transform 1 0 22172 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_234
timestamp 1649977179
transform 1 0 22632 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_242
timestamp 1649977179
transform 1 0 23368 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_258
timestamp 1649977179
transform 1 0 24840 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_274
timestamp 1649977179
transform 1 0 26312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_283
timestamp 1649977179
transform 1 0 27140 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_291
timestamp 1649977179
transform 1 0 27876 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_294
timestamp 1649977179
transform 1 0 28152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_300
timestamp 1649977179
transform 1 0 28704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_304
timestamp 1649977179
transform 1 0 29072 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_40
timestamp 1649977179
transform 1 0 4784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1649977179
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_67
timestamp 1649977179
transform 1 0 7268 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_78
timestamp 1649977179
transform 1 0 8280 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_85
timestamp 1649977179
transform 1 0 8924 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_91
timestamp 1649977179
transform 1 0 9476 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_99
timestamp 1649977179
transform 1 0 10212 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_102
timestamp 1649977179
transform 1 0 10488 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1649977179
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_118
timestamp 1649977179
transform 1 0 11960 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_126
timestamp 1649977179
transform 1 0 12696 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_129
timestamp 1649977179
transform 1 0 12972 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_138
timestamp 1649977179
transform 1 0 13800 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_147
timestamp 1649977179
transform 1 0 14628 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_159
timestamp 1649977179
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_171
timestamp 1649977179
transform 1 0 16836 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_177
timestamp 1649977179
transform 1 0 17388 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_183
timestamp 1649977179
transform 1 0 17940 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_189
timestamp 1649977179
transform 1 0 18492 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_204
timestamp 1649977179
transform 1 0 19872 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_212
timestamp 1649977179
transform 1 0 20608 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_216
timestamp 1649977179
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_227
timestamp 1649977179
transform 1 0 21988 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_233
timestamp 1649977179
transform 1 0 22540 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_247
timestamp 1649977179
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_259
timestamp 1649977179
transform 1 0 24932 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_265
timestamp 1649977179
transform 1 0 25484 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1649977179
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_289
timestamp 1649977179
transform 1 0 27692 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_295
timestamp 1649977179
transform 1 0 28244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_301
timestamp 1649977179
transform 1 0 28796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_7
timestamp 1649977179
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1649977179
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_44
timestamp 1649977179
transform 1 0 5152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_51
timestamp 1649977179
transform 1 0 5796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_57
timestamp 1649977179
transform 1 0 6348 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_63
timestamp 1649977179
transform 1 0 6900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_74
timestamp 1649977179
transform 1 0 7912 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1649977179
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1649977179
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_92
timestamp 1649977179
transform 1 0 9568 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_103
timestamp 1649977179
transform 1 0 10580 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_114
timestamp 1649977179
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_125
timestamp 1649977179
transform 1 0 12604 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1649977179
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_146
timestamp 1649977179
transform 1 0 14536 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_152
timestamp 1649977179
transform 1 0 15088 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_160
timestamp 1649977179
transform 1 0 15824 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_166
timestamp 1649977179
transform 1 0 16376 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_175
timestamp 1649977179
transform 1 0 17204 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_183
timestamp 1649977179
transform 1 0 17940 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1649977179
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_206
timestamp 1649977179
transform 1 0 20056 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_217
timestamp 1649977179
transform 1 0 21068 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_223
timestamp 1649977179
transform 1 0 21620 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_229
timestamp 1649977179
transform 1 0 22172 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_235
timestamp 1649977179
transform 1 0 22724 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_241
timestamp 1649977179
transform 1 0 23276 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1649977179
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_256
timestamp 1649977179
transform 1 0 24656 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_264
timestamp 1649977179
transform 1 0 25392 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_272
timestamp 1649977179
transform 1 0 26128 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_284
timestamp 1649977179
transform 1 0 27232 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_292
timestamp 1649977179
transform 1 0 27968 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_13
timestamp 1649977179
transform 1 0 2300 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_25
timestamp 1649977179
transform 1 0 3404 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_37
timestamp 1649977179
transform 1 0 4508 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_43
timestamp 1649977179
transform 1 0 5060 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_46
timestamp 1649977179
transform 1 0 5336 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1649977179
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_65
timestamp 1649977179
transform 1 0 7084 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_74
timestamp 1649977179
transform 1 0 7912 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_80
timestamp 1649977179
transform 1 0 8464 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_92
timestamp 1649977179
transform 1 0 9568 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_95
timestamp 1649977179
transform 1 0 9844 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_101
timestamp 1649977179
transform 1 0 10396 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1649977179
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_120
timestamp 1649977179
transform 1 0 12144 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_127
timestamp 1649977179
transform 1 0 12788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_133
timestamp 1649977179
transform 1 0 13340 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_143
timestamp 1649977179
transform 1 0 14260 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_151
timestamp 1649977179
transform 1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_160
timestamp 1649977179
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_176
timestamp 1649977179
transform 1 0 17296 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_182
timestamp 1649977179
transform 1 0 17848 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_188
timestamp 1649977179
transform 1 0 18400 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_199
timestamp 1649977179
transform 1 0 19412 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_211
timestamp 1649977179
transform 1 0 20516 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1649977179
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_227
timestamp 1649977179
transform 1 0 21988 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_231
timestamp 1649977179
transform 1 0 22356 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_236
timestamp 1649977179
transform 1 0 22816 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_248
timestamp 1649977179
transform 1 0 23920 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_262
timestamp 1649977179
transform 1 0 25208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1649977179
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 1649977179
transform 1 0 28796 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_73
timestamp 1649977179
transform 1 0 7820 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_76
timestamp 1649977179
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_90
timestamp 1649977179
transform 1 0 9384 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_96
timestamp 1649977179
transform 1 0 9936 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_105
timestamp 1649977179
transform 1 0 10764 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_114
timestamp 1649977179
transform 1 0 11592 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_122
timestamp 1649977179
transform 1 0 12328 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_126
timestamp 1649977179
transform 1 0 12696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_132
timestamp 1649977179
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_152
timestamp 1649977179
transform 1 0 15088 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_160
timestamp 1649977179
transform 1 0 15824 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_166
timestamp 1649977179
transform 1 0 16376 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_172
timestamp 1649977179
transform 1 0 16928 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_184
timestamp 1649977179
transform 1 0 18032 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_208
timestamp 1649977179
transform 1 0 20240 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_219
timestamp 1649977179
transform 1 0 21252 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_229
timestamp 1649977179
transform 1 0 22172 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_241
timestamp 1649977179
transform 1 0 23276 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1649977179
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_267
timestamp 1649977179
transform 1 0 25668 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_279
timestamp 1649977179
transform 1 0 26772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_291
timestamp 1649977179
transform 1 0 27876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_303
timestamp 1649977179
transform 1 0 28980 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_74
timestamp 1649977179
transform 1 0 7912 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_82
timestamp 1649977179
transform 1 0 8648 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_91
timestamp 1649977179
transform 1 0 9476 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_99
timestamp 1649977179
transform 1 0 10212 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1649977179
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_124
timestamp 1649977179
transform 1 0 12512 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_135
timestamp 1649977179
transform 1 0 13524 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_141
timestamp 1649977179
transform 1 0 14076 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_147
timestamp 1649977179
transform 1 0 14628 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_171
timestamp 1649977179
transform 1 0 16836 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_183
timestamp 1649977179
transform 1 0 17940 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_191
timestamp 1649977179
transform 1 0 18676 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_197
timestamp 1649977179
transform 1 0 19228 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_208
timestamp 1649977179
transform 1 0 20240 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_214
timestamp 1649977179
transform 1 0 20792 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1649977179
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_234
timestamp 1649977179
transform 1 0 22632 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_245
timestamp 1649977179
transform 1 0 23644 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_256
timestamp 1649977179
transform 1 0 24656 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_262
timestamp 1649977179
transform 1 0 25208 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1649977179
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_289
timestamp 1649977179
transform 1 0 27692 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_301
timestamp 1649977179
transform 1 0 28796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_7
timestamp 1649977179
transform 1 0 1748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1649977179
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_49
timestamp 1649977179
transform 1 0 5612 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_58
timestamp 1649977179
transform 1 0 6440 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_67
timestamp 1649977179
transform 1 0 7268 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_75
timestamp 1649977179
transform 1 0 8004 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_79
timestamp 1649977179
transform 1 0 8372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_92
timestamp 1649977179
transform 1 0 9568 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_98
timestamp 1649977179
transform 1 0 10120 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_104
timestamp 1649977179
transform 1 0 10672 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_110
timestamp 1649977179
transform 1 0 11224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_131
timestamp 1649977179
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1649977179
transform 1 0 14444 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_156
timestamp 1649977179
transform 1 0 15456 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_160
timestamp 1649977179
transform 1 0 15824 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_166
timestamp 1649977179
transform 1 0 16376 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_174
timestamp 1649977179
transform 1 0 17112 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_178
timestamp 1649977179
transform 1 0 17480 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_188
timestamp 1649977179
transform 1 0 18400 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_203
timestamp 1649977179
transform 1 0 19780 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_215
timestamp 1649977179
transform 1 0 20884 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_225
timestamp 1649977179
transform 1 0 21804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_243
timestamp 1649977179
transform 1 0 23460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_256
timestamp 1649977179
transform 1 0 24656 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_262
timestamp 1649977179
transform 1 0 25208 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_274
timestamp 1649977179
transform 1 0 26312 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_286
timestamp 1649977179
transform 1 0 27416 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_298
timestamp 1649977179
transform 1 0 28520 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_304
timestamp 1649977179
transform 1 0 29072 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_11
timestamp 1649977179
transform 1 0 2116 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_17
timestamp 1649977179
transform 1 0 2668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_29
timestamp 1649977179
transform 1 0 3772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_41
timestamp 1649977179
transform 1 0 4876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1649977179
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_64
timestamp 1649977179
transform 1 0 6992 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_77
timestamp 1649977179
transform 1 0 8188 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_88
timestamp 1649977179
transform 1 0 9200 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_94
timestamp 1649977179
transform 1 0 9752 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_100
timestamp 1649977179
transform 1 0 10304 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_121
timestamp 1649977179
transform 1 0 12236 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_133
timestamp 1649977179
transform 1 0 13340 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_145
timestamp 1649977179
transform 1 0 14444 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_160
timestamp 1649977179
transform 1 0 15824 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_176
timestamp 1649977179
transform 1 0 17296 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_184
timestamp 1649977179
transform 1 0 18032 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_198
timestamp 1649977179
transform 1 0 19320 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_211
timestamp 1649977179
transform 1 0 20516 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1649977179
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_232
timestamp 1649977179
transform 1 0 22448 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_242
timestamp 1649977179
transform 1 0 23368 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_248
timestamp 1649977179
transform 1 0 23920 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_260
timestamp 1649977179
transform 1 0 25024 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1649977179
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_297
timestamp 1649977179
transform 1 0 28428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_7
timestamp 1649977179
transform 1 0 1748 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_17
timestamp 1649977179
transform 1 0 2668 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1649977179
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_90
timestamp 1649977179
transform 1 0 9384 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_102
timestamp 1649977179
transform 1 0 10488 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_110
timestamp 1649977179
transform 1 0 11224 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_115
timestamp 1649977179
transform 1 0 11684 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_128
timestamp 1649977179
transform 1 0 12880 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_169
timestamp 1649977179
transform 1 0 16652 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_175
timestamp 1649977179
transform 1 0 17204 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_179
timestamp 1649977179
transform 1 0 17572 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_185
timestamp 1649977179
transform 1 0 18124 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_191
timestamp 1649977179
transform 1 0 18676 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_203
timestamp 1649977179
transform 1 0 19780 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_206
timestamp 1649977179
transform 1 0 20056 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_218
timestamp 1649977179
transform 1 0 21160 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_232
timestamp 1649977179
transform 1 0 22448 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_238
timestamp 1649977179
transform 1 0 23000 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1649977179
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_255
timestamp 1649977179
transform 1 0 24564 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_267
timestamp 1649977179
transform 1 0 25668 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_279
timestamp 1649977179
transform 1 0 26772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_283
timestamp 1649977179
transform 1 0 27140 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_289
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_301
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_13
timestamp 1649977179
transform 1 0 2300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_23
timestamp 1649977179
transform 1 0 3220 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_29
timestamp 1649977179
transform 1 0 3772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_41
timestamp 1649977179
transform 1 0 4876 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp 1649977179
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_62
timestamp 1649977179
transform 1 0 6808 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_72
timestamp 1649977179
transform 1 0 7728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_85
timestamp 1649977179
transform 1 0 8924 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_91
timestamp 1649977179
transform 1 0 9476 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_103
timestamp 1649977179
transform 1 0 10580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_119
timestamp 1649977179
transform 1 0 12052 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_131
timestamp 1649977179
transform 1 0 13156 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_136
timestamp 1649977179
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_145
timestamp 1649977179
transform 1 0 14444 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_153
timestamp 1649977179
transform 1 0 15180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_163
timestamp 1649977179
transform 1 0 16100 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_177
timestamp 1649977179
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_180
timestamp 1649977179
transform 1 0 17664 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_184
timestamp 1649977179
transform 1 0 18032 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_189
timestamp 1649977179
transform 1 0 18492 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_195
timestamp 1649977179
transform 1 0 19044 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_199
timestamp 1649977179
transform 1 0 19412 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_210
timestamp 1649977179
transform 1 0 20424 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1649977179
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_231
timestamp 1649977179
transform 1 0 22356 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_243
timestamp 1649977179
transform 1 0 23460 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_251
timestamp 1649977179
transform 1 0 24196 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_253
timestamp 1649977179
transform 1 0 24380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_259
timestamp 1649977179
transform 1 0 24932 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_271
timestamp 1649977179
transform 1 0 26036 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1649977179
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_285
timestamp 1649977179
transform 1 0 27324 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_301
timestamp 1649977179
transform 1 0 28796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 29440 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 29440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 29440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 29440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 29440 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 29440 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 29440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 29440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 29440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 29440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 29440 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 29440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 29440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 29440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 29440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 29440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 29440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 29440 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 29440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 29440 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 29440 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 29440 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 29440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 29440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 29440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 29440 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 29440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 29440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 29440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 29440 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 29440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 29440 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 29440 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 29440 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 29440 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 29440 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 29440 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 29440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 29440 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 29440 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 29440 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 29440 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 29440 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 29440 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 29440 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 29440 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 29440 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 29440 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 3680 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 8832 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 24288 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _0578_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19596 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0579_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19596 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0580_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24932 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0581_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 25668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0582_
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0583_
timestamp 1649977179
transform 1 0 17940 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0584_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18676 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0585_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0586_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22080 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0587_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19688 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _0588_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0589_
timestamp 1649977179
transform -1 0 21160 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0590_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23000 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _0591_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22448 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _0592_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25944 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0593_
timestamp 1649977179
transform -1 0 26036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0594_
timestamp 1649977179
transform -1 0 25576 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand4b_2  _0595_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 25576 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _0596_
timestamp 1649977179
transform -1 0 21160 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0597_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20976 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0598_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19964 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _0599_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0600_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17848 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _0601_
timestamp 1649977179
transform 1 0 12788 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0602_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19688 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _0603_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18400 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_4  _0604_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21620 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0605_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19320 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0606_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18492 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0607_
timestamp 1649977179
transform 1 0 17388 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0608_
timestamp 1649977179
transform -1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _0609_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0610_
timestamp 1649977179
transform 1 0 17848 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0611_
timestamp 1649977179
transform 1 0 16744 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0612_
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0613_
timestamp 1649977179
transform -1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0614_
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0615_
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0616_
timestamp 1649977179
transform 1 0 16652 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0617_
timestamp 1649977179
transform -1 0 16284 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0618_
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0619_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0620_
timestamp 1649977179
transform 1 0 14444 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0621_
timestamp 1649977179
transform 1 0 14628 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0622_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 25300 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0623_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0624_
timestamp 1649977179
transform -1 0 14444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0625_
timestamp 1649977179
transform -1 0 13892 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0626_
timestamp 1649977179
transform -1 0 13064 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0627_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17112 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0628_
timestamp 1649977179
transform 1 0 21252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0629_
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _0630_
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0631_
timestamp 1649977179
transform -1 0 19412 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0632_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0633_
timestamp 1649977179
transform 1 0 18216 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1649977179
transform 1 0 16560 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0635_
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0636_
timestamp 1649977179
transform 1 0 27968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0637_
timestamp 1649977179
transform 1 0 17848 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0638_
timestamp 1649977179
transform -1 0 17388 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0639_
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _0640_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17112 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _0641_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25576 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0642_
timestamp 1649977179
transform 1 0 21804 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0643_
timestamp 1649977179
transform 1 0 27876 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0644_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25668 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _0645_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23920 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0646_
timestamp 1649977179
transform 1 0 21712 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0647_
timestamp 1649977179
transform -1 0 24840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0648_
timestamp 1649977179
transform -1 0 26312 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _0649_
timestamp 1649977179
transform 1 0 24288 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0650_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22448 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0651_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0652_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0653_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27140 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0654_
timestamp 1649977179
transform -1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _0655_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25208 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _0656_
timestamp 1649977179
transform -1 0 22908 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0657_
timestamp 1649977179
transform -1 0 22632 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0658_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0659_
timestamp 1649977179
transform -1 0 24656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0660_
timestamp 1649977179
transform 1 0 22908 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0662_
timestamp 1649977179
transform 1 0 21896 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0663_
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0664_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15732 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0665_
timestamp 1649977179
transform 1 0 17940 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0666_
timestamp 1649977179
transform -1 0 13432 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0667_
timestamp 1649977179
transform -1 0 23644 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0668_
timestamp 1649977179
transform -1 0 22724 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0669_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22172 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0670_
timestamp 1649977179
transform 1 0 21620 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0671_
timestamp 1649977179
transform -1 0 23000 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0672_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20792 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0673_
timestamp 1649977179
transform 1 0 20516 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _0674_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0675_
timestamp 1649977179
transform -1 0 23920 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _0676_
timestamp 1649977179
transform -1 0 21436 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0677_
timestamp 1649977179
transform 1 0 19872 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0678_
timestamp 1649977179
transform 1 0 12788 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0679_
timestamp 1649977179
transform -1 0 13524 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _0680_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22448 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _0681_
timestamp 1649977179
transform -1 0 21068 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0682_
timestamp 1649977179
transform 1 0 4876 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0683_
timestamp 1649977179
transform -1 0 28704 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _0684_
timestamp 1649977179
transform -1 0 20976 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0685_
timestamp 1649977179
transform -1 0 12880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0686_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13892 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0687_
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0688_
timestamp 1649977179
transform 1 0 24196 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0689_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 25116 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _0690_
timestamp 1649977179
transform -1 0 23184 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0691_
timestamp 1649977179
transform 1 0 23368 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0692_
timestamp 1649977179
transform -1 0 23552 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0693_
timestamp 1649977179
transform -1 0 19964 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0694_
timestamp 1649977179
transform -1 0 14536 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0695_
timestamp 1649977179
transform 1 0 15456 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0696_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15456 0 1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_4  _0697_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17664 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0698_
timestamp 1649977179
transform 1 0 19688 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0699_
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__or2b_1  _0700_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22816 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0701_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21896 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _0702_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18124 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0703_
timestamp 1649977179
transform 1 0 19688 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0704_
timestamp 1649977179
transform -1 0 24656 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0705_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0706_
timestamp 1649977179
transform -1 0 20240 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0707_
timestamp 1649977179
transform -1 0 21344 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0708_
timestamp 1649977179
transform 1 0 19320 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0709_
timestamp 1649977179
transform -1 0 20976 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0710_
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0711_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19872 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0712_
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0713_
timestamp 1649977179
transform 1 0 20424 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0714_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20608 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0715_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20516 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0716_
timestamp 1649977179
transform 1 0 19596 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0717_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0718_
timestamp 1649977179
transform 1 0 18124 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0719_
timestamp 1649977179
transform -1 0 14076 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_4  _0720_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 25668 0 1 27200
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_1  _0721_
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1649977179
transform 1 0 14352 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0723_
timestamp 1649977179
transform 1 0 15364 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0724_
timestamp 1649977179
transform 1 0 15364 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0725_
timestamp 1649977179
transform -1 0 18124 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0726_
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0727_
timestamp 1649977179
transform -1 0 15824 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0728_
timestamp 1649977179
transform 1 0 12972 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0729_
timestamp 1649977179
transform 1 0 10304 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0730_
timestamp 1649977179
transform -1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0731_
timestamp 1649977179
transform -1 0 15824 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0732_
timestamp 1649977179
transform -1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0733_
timestamp 1649977179
transform -1 0 18308 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0734_
timestamp 1649977179
transform 1 0 16376 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0735_
timestamp 1649977179
transform 1 0 14260 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0736_
timestamp 1649977179
transform -1 0 16652 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0737_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17940 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1649977179
transform 1 0 15456 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _0739_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0740_
timestamp 1649977179
transform -1 0 14996 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0741_
timestamp 1649977179
transform -1 0 15916 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1649977179
transform -1 0 23644 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0743_
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0744_
timestamp 1649977179
transform -1 0 23460 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0745_
timestamp 1649977179
transform -1 0 19412 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0746_
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1649977179
transform -1 0 23644 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0748_
timestamp 1649977179
transform -1 0 22816 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0749_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16468 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0750_
timestamp 1649977179
transform -1 0 16376 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0751_
timestamp 1649977179
transform -1 0 22172 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0752_
timestamp 1649977179
transform -1 0 11040 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0753_
timestamp 1649977179
transform -1 0 11592 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0754_
timestamp 1649977179
transform 1 0 10304 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0755_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11592 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a311o_1  _0756_
timestamp 1649977179
transform 1 0 18032 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0757_
timestamp 1649977179
transform -1 0 12788 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0758_
timestamp 1649977179
transform 1 0 11592 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0759_
timestamp 1649977179
transform -1 0 11960 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0760_
timestamp 1649977179
transform 1 0 9936 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0761_
timestamp 1649977179
transform 1 0 11960 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0762_
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0763_
timestamp 1649977179
transform -1 0 13800 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0764_
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0765_
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 1649977179
transform 1 0 12512 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0767_
timestamp 1649977179
transform -1 0 12696 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0768_
timestamp 1649977179
transform -1 0 13524 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0770_
timestamp 1649977179
transform -1 0 21252 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0771_
timestamp 1649977179
transform 1 0 17848 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0772_
timestamp 1649977179
transform -1 0 15272 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _0773_
timestamp 1649977179
transform -1 0 28796 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0774_
timestamp 1649977179
transform 1 0 16652 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _0775_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0776_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0777_
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0778_
timestamp 1649977179
transform -1 0 15272 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0780_
timestamp 1649977179
transform -1 0 26404 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_4  _0781_
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1649977179
transform 1 0 25024 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0783_
timestamp 1649977179
transform -1 0 17480 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0784_
timestamp 1649977179
transform -1 0 15088 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0785_
timestamp 1649977179
transform 1 0 14536 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 1649977179
transform 1 0 27508 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0787_
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0788_
timestamp 1649977179
transform -1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1649977179
transform 1 0 24748 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _0790_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _0791_
timestamp 1649977179
transform -1 0 23276 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0792_
timestamp 1649977179
transform 1 0 12604 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0793_
timestamp 1649977179
transform -1 0 9200 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0794_
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0795_
timestamp 1649977179
transform 1 0 9108 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0796_
timestamp 1649977179
transform -1 0 12052 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0797_
timestamp 1649977179
transform 1 0 4508 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0798_
timestamp 1649977179
transform -1 0 5152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0799_
timestamp 1649977179
transform -1 0 5796 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0800_
timestamp 1649977179
transform -1 0 5336 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0801_
timestamp 1649977179
transform 1 0 5152 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0802_
timestamp 1649977179
transform -1 0 5152 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0803_
timestamp 1649977179
transform 1 0 10948 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0804_
timestamp 1649977179
transform 1 0 7820 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0805_
timestamp 1649977179
transform 1 0 8004 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0806_
timestamp 1649977179
transform 1 0 12144 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0807_
timestamp 1649977179
transform -1 0 14720 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0808_
timestamp 1649977179
transform 1 0 11868 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _0809_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9752 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0810_
timestamp 1649977179
transform 1 0 9568 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _0811_
timestamp 1649977179
transform 1 0 10120 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _0812_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11408 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0813_
timestamp 1649977179
transform 1 0 7636 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _0814_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6992 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1649977179
transform -1 0 6992 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0816_
timestamp 1649977179
transform -1 0 11040 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0817_
timestamp 1649977179
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0818_
timestamp 1649977179
transform -1 0 7636 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0819_
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0820_
timestamp 1649977179
transform -1 0 6532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1649977179
transform -1 0 5428 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0822_
timestamp 1649977179
transform 1 0 4324 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0823_
timestamp 1649977179
transform 1 0 4140 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1649977179
transform 1 0 5520 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1649977179
transform 1 0 27324 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0826_
timestamp 1649977179
transform -1 0 27324 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp 1649977179
transform 1 0 26128 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0828_
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _0829_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23092 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0830_
timestamp 1649977179
transform -1 0 8924 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0831_
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0832_
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0833_
timestamp 1649977179
transform -1 0 7268 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0834_
timestamp 1649977179
transform 1 0 11408 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0835_
timestamp 1649977179
transform -1 0 10212 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0836_
timestamp 1649977179
transform 1 0 9292 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0837_
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0838_
timestamp 1649977179
transform -1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0839_
timestamp 1649977179
transform 1 0 12420 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0840_
timestamp 1649977179
transform -1 0 9936 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0841_
timestamp 1649977179
transform -1 0 7912 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0842_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7912 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0844_
timestamp 1649977179
transform -1 0 9568 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0845_
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0846_
timestamp 1649977179
transform -1 0 9200 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _0847_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4968 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0848_
timestamp 1649977179
transform -1 0 6532 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0849_
timestamp 1649977179
transform -1 0 4784 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 1649977179
transform -1 0 4508 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0851_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4232 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0852_
timestamp 1649977179
transform 1 0 3772 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0853_
timestamp 1649977179
transform 1 0 3220 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0854_
timestamp 1649977179
transform -1 0 8188 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _0855_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7452 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0856_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7636 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0857_
timestamp 1649977179
transform -1 0 7084 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1649977179
transform 1 0 27416 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0859_
timestamp 1649977179
transform -1 0 27968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 1649977179
transform 1 0 26404 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp 1649977179
transform 1 0 22632 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0862_
timestamp 1649977179
transform 1 0 12604 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0863_
timestamp 1649977179
transform -1 0 15088 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0864_
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0865_
timestamp 1649977179
transform 1 0 9476 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0866_
timestamp 1649977179
transform -1 0 11040 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0867_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9660 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0868_
timestamp 1649977179
transform -1 0 10304 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0869_
timestamp 1649977179
transform 1 0 11592 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0870_
timestamp 1649977179
transform 1 0 10764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0871_
timestamp 1649977179
transform 1 0 5704 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0872_
timestamp 1649977179
transform 1 0 5612 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0873_
timestamp 1649977179
transform -1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1649977179
transform -1 0 8464 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1649977179
transform -1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0876_
timestamp 1649977179
transform 1 0 6716 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0877_
timestamp 1649977179
transform 1 0 3864 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0878_
timestamp 1649977179
transform 1 0 28152 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0879_
timestamp 1649977179
transform -1 0 28244 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0880_
timestamp 1649977179
transform -1 0 28520 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0881_
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0882_
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0883_
timestamp 1649977179
transform 1 0 24104 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0884_
timestamp 1649977179
transform -1 0 14352 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0885_
timestamp 1649977179
transform 1 0 12880 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0886_
timestamp 1649977179
transform -1 0 13708 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0887_
timestamp 1649977179
transform -1 0 10028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0888_
timestamp 1649977179
transform -1 0 9936 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _0889_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9476 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0890_
timestamp 1649977179
transform 1 0 11592 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0891_
timestamp 1649977179
transform 1 0 11500 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1649977179
transform -1 0 1932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0893_
timestamp 1649977179
transform -1 0 2852 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0894_
timestamp 1649977179
transform -1 0 2576 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0895_
timestamp 1649977179
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0896_
timestamp 1649977179
transform -1 0 4232 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0897_
timestamp 1649977179
transform 1 0 3864 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_2  _0898_
timestamp 1649977179
transform 1 0 4140 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0899_
timestamp 1649977179
transform 1 0 9108 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0900_
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0901_
timestamp 1649977179
transform -1 0 9292 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0902_
timestamp 1649977179
transform -1 0 6624 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0903_
timestamp 1649977179
transform -1 0 7636 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0904_
timestamp 1649977179
transform -1 0 7084 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0906_
timestamp 1649977179
transform 1 0 5060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0907_
timestamp 1649977179
transform -1 0 4692 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0908_
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1649977179
transform -1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0910_
timestamp 1649977179
transform 1 0 2760 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _0911_
timestamp 1649977179
transform -1 0 3864 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1649977179
transform 1 0 4232 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0913_
timestamp 1649977179
transform -1 0 4784 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0914_
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0915_
timestamp 1649977179
transform -1 0 4324 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0916_
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0917_
timestamp 1649977179
transform 1 0 27416 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0918_
timestamp 1649977179
transform -1 0 27784 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0919_
timestamp 1649977179
transform 1 0 27140 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0921_
timestamp 1649977179
transform 1 0 24104 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0924_
timestamp 1649977179
transform -1 0 10672 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0925_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22908 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0926_
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0927_
timestamp 1649977179
transform -1 0 10764 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0928_
timestamp 1649977179
transform -1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0929_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_2  _0930_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13524 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _0931_
timestamp 1649977179
transform 1 0 6532 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0932_
timestamp 1649977179
transform 1 0 6164 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _0933_
timestamp 1649977179
transform 1 0 7912 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0934_
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0935_
timestamp 1649977179
transform -1 0 7544 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0936_
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0937_
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0938_
timestamp 1649977179
transform 1 0 6900 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0939_
timestamp 1649977179
transform -1 0 25024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 1649977179
transform 1 0 27324 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0941_
timestamp 1649977179
transform 1 0 27508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 1649977179
transform 1 0 27232 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0943_
timestamp 1649977179
transform -1 0 26680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0944_
timestamp 1649977179
transform -1 0 24656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0945_
timestamp 1649977179
transform -1 0 23920 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0946_
timestamp 1649977179
transform 1 0 24196 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0947_
timestamp 1649977179
transform 1 0 9844 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0948_
timestamp 1649977179
transform -1 0 11960 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0949_
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0950_
timestamp 1649977179
transform 1 0 12604 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0951_
timestamp 1649977179
transform 1 0 12052 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1649977179
transform -1 0 5888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0953_
timestamp 1649977179
transform 1 0 5060 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0954_
timestamp 1649977179
transform -1 0 6164 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0955_
timestamp 1649977179
transform -1 0 5060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0956_
timestamp 1649977179
transform -1 0 5060 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0957_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0958_
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0959_
timestamp 1649977179
transform 1 0 10304 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0960_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7728 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1649977179
transform 1 0 6808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0962_
timestamp 1649977179
transform -1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0963_
timestamp 1649977179
transform -1 0 9108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0964_
timestamp 1649977179
transform -1 0 9476 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0965_
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1649977179
transform -1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0967_
timestamp 1649977179
transform 1 0 6808 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0968_
timestamp 1649977179
transform 1 0 5796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0969_
timestamp 1649977179
transform 1 0 4140 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0970_
timestamp 1649977179
transform 1 0 4140 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0972_
timestamp 1649977179
transform 1 0 4508 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0973_
timestamp 1649977179
transform 1 0 4600 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0974_
timestamp 1649977179
transform 1 0 5336 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0975_
timestamp 1649977179
transform -1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0976_
timestamp 1649977179
transform 1 0 7728 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0977_
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0978_
timestamp 1649977179
transform -1 0 27416 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0979_
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0980_
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0981_
timestamp 1649977179
transform 1 0 24932 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0982_
timestamp 1649977179
transform -1 0 24380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0983_
timestamp 1649977179
transform -1 0 17020 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 1649977179
transform -1 0 13616 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0985_
timestamp 1649977179
transform -1 0 11040 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _0986_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11040 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _0987_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14076 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0988_
timestamp 1649977179
transform -1 0 14720 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0989_
timestamp 1649977179
transform -1 0 8464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0990_
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0991_
timestamp 1649977179
transform 1 0 6992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_4  _0993_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _0994_
timestamp 1649977179
transform -1 0 10488 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0995_
timestamp 1649977179
transform 1 0 10120 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_1  _0996_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0997_
timestamp 1649977179
transform -1 0 8280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0998_
timestamp 1649977179
transform -1 0 9292 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0999_
timestamp 1649977179
transform -1 0 27876 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1000_
timestamp 1649977179
transform -1 0 27968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1001_
timestamp 1649977179
transform 1 0 27232 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1002_
timestamp 1649977179
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1003_
timestamp 1649977179
transform -1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1649977179
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1005_
timestamp 1649977179
transform -1 0 25116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1006_
timestamp 1649977179
transform 1 0 11868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1007_
timestamp 1649977179
transform -1 0 13984 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1008_
timestamp 1649977179
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1009_
timestamp 1649977179
transform 1 0 10028 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1010_
timestamp 1649977179
transform 1 0 10304 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1011_
timestamp 1649977179
transform -1 0 11868 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1012_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1013_
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1649977179
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1649977179
transform -1 0 8004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1016_
timestamp 1649977179
transform -1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1017_
timestamp 1649977179
transform -1 0 7268 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 1649977179
transform -1 0 6716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1019_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5336 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1020_
timestamp 1649977179
transform -1 0 5428 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1021_
timestamp 1649977179
transform 1 0 5704 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1022_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1023_
timestamp 1649977179
transform -1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1024_
timestamp 1649977179
transform 1 0 13432 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1025_
timestamp 1649977179
transform 1 0 27784 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1026_
timestamp 1649977179
transform -1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1027_
timestamp 1649977179
transform 1 0 27140 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp 1649977179
transform 1 0 24840 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1029_
timestamp 1649977179
transform -1 0 24104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1030_
timestamp 1649977179
transform -1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1031_
timestamp 1649977179
transform -1 0 13524 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1032_
timestamp 1649977179
transform -1 0 12788 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1033_
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1034_
timestamp 1649977179
transform 1 0 10672 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1035_
timestamp 1649977179
transform -1 0 12788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1036_
timestamp 1649977179
transform 1 0 13156 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1037_
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1038_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1649977179
transform -1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1040_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1041_
timestamp 1649977179
transform -1 0 11040 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1042_
timestamp 1649977179
transform -1 0 4416 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1043_
timestamp 1649977179
transform 1 0 4784 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1044_
timestamp 1649977179
transform 1 0 5520 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1045_
timestamp 1649977179
transform -1 0 5888 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1046_
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1047_
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1048_
timestamp 1649977179
transform -1 0 12972 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1049_
timestamp 1649977179
transform 1 0 12328 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1050_
timestamp 1649977179
transform 1 0 12696 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1051_
timestamp 1649977179
transform -1 0 4876 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o311a_1  _1052_
timestamp 1649977179
transform 1 0 10120 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1053_
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1054_
timestamp 1649977179
transform -1 0 17112 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1055_
timestamp 1649977179
transform -1 0 15088 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1056_
timestamp 1649977179
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1057_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1058_
timestamp 1649977179
transform 1 0 14168 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1649977179
transform -1 0 15272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1060_
timestamp 1649977179
transform 1 0 14076 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1061_
timestamp 1649977179
transform 1 0 14168 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1062_
timestamp 1649977179
transform -1 0 14444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _1063_
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1064_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 1649977179
transform -1 0 15456 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1066_
timestamp 1649977179
transform 1 0 14536 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1067_
timestamp 1649977179
transform -1 0 16192 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1068_
timestamp 1649977179
transform -1 0 16192 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1069_
timestamp 1649977179
transform -1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1070_
timestamp 1649977179
transform 1 0 14812 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1071_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1072_
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1073_
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1074_
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1075_
timestamp 1649977179
transform 1 0 26496 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1076_
timestamp 1649977179
transform -1 0 15364 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1077_
timestamp 1649977179
transform -1 0 14996 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1078_
timestamp 1649977179
transform -1 0 9660 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1079_
timestamp 1649977179
transform -1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1080_
timestamp 1649977179
transform 1 0 20148 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1081_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1082_
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1083_
timestamp 1649977179
transform -1 0 15916 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1084_
timestamp 1649977179
transform 1 0 16652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1085_
timestamp 1649977179
transform -1 0 17572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1649977179
transform -1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1087_
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1088_
timestamp 1649977179
transform -1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1089_
timestamp 1649977179
transform -1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1090_
timestamp 1649977179
transform -1 0 15180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1091_
timestamp 1649977179
transform 1 0 15456 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1092_
timestamp 1649977179
transform -1 0 17940 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1649977179
transform -1 0 19228 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _1094_
timestamp 1649977179
transform -1 0 18768 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1095_
timestamp 1649977179
transform -1 0 20148 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1096_
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1097_
timestamp 1649977179
transform 1 0 15272 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1098_
timestamp 1649977179
transform -1 0 16744 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1099_
timestamp 1649977179
transform -1 0 25760 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1100_
timestamp 1649977179
transform 1 0 25668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1101_
timestamp 1649977179
transform 1 0 25944 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1102_
timestamp 1649977179
transform 1 0 25208 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1103_
timestamp 1649977179
transform -1 0 17940 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1104_
timestamp 1649977179
transform 1 0 16928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1105_
timestamp 1649977179
transform -1 0 17848 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1649977179
transform 1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1107_
timestamp 1649977179
transform -1 0 16928 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1649977179
transform -1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1109_
timestamp 1649977179
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1110_
timestamp 1649977179
transform -1 0 23920 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1111_
timestamp 1649977179
transform 1 0 22632 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1112_
timestamp 1649977179
transform -1 0 20976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1113_
timestamp 1649977179
transform -1 0 21068 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1114_
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1115_
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1116_
timestamp 1649977179
transform -1 0 22356 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1117_
timestamp 1649977179
transform 1 0 20424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1118_
timestamp 1649977179
transform -1 0 22264 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1119_
timestamp 1649977179
transform 1 0 20976 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1120_
timestamp 1649977179
transform -1 0 23736 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1121_
timestamp 1649977179
transform -1 0 25576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1122_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24840 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1123_
timestamp 1649977179
transform 1 0 24932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1124_
timestamp 1649977179
transform -1 0 24196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1125_
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1126_
timestamp 1649977179
transform 1 0 22724 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1127_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1128_
timestamp 1649977179
transform -1 0 23736 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1129_
timestamp 1649977179
transform -1 0 22540 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1130_
timestamp 1649977179
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1131_
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1132_
timestamp 1649977179
transform 1 0 21896 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1133_
timestamp 1649977179
transform -1 0 22908 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _1134_
timestamp 1649977179
transform -1 0 22540 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_4  _1135_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__xnor2_1  _1136_
timestamp 1649977179
transform 1 0 1748 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1137_
timestamp 1649977179
transform -1 0 2576 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1138_
timestamp 1649977179
transform -1 0 2392 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1139_
timestamp 1649977179
transform 1 0 5796 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1140_
timestamp 1649977179
transform 1 0 7544 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1141_
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1142_
timestamp 1649977179
transform -1 0 9568 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1143_
timestamp 1649977179
transform -1 0 6992 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1144_
timestamp 1649977179
transform -1 0 2392 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1145_
timestamp 1649977179
transform -1 0 2392 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1146_
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1147_
timestamp 1649977179
transform -1 0 2392 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1148_
timestamp 1649977179
transform 1 0 1932 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1149_
timestamp 1649977179
transform 1 0 2024 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1150_
timestamp 1649977179
transform 1 0 2208 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _1151_
timestamp 1649977179
transform -1 0 19412 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1152_
timestamp 1649977179
transform -1 0 13248 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1153_
timestamp 1649977179
transform -1 0 20148 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1154_
timestamp 1649977179
transform 1 0 19872 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1155_
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1156_
timestamp 1649977179
transform 1 0 24932 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1157_
timestamp 1649977179
transform 1 0 24472 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1158_
timestamp 1649977179
transform 1 0 23184 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1159_
timestamp 1649977179
transform 1 0 19596 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1160_
timestamp 1649977179
transform -1 0 21160 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1161_
timestamp 1649977179
transform -1 0 21804 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1162_
timestamp 1649977179
transform 1 0 20976 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1163_
timestamp 1649977179
transform 1 0 20976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1164_
timestamp 1649977179
transform 1 0 20056 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1649977179
transform 1 0 2116 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1166_
timestamp 1649977179
transform -1 0 3404 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1167_
timestamp 1649977179
transform -1 0 9476 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1168_
timestamp 1649977179
transform -1 0 7268 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1169_
timestamp 1649977179
transform -1 0 6624 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1170_
timestamp 1649977179
transform -1 0 2944 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _1171_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1932 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1172_
timestamp 1649977179
transform 1 0 24104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1173_
timestamp 1649977179
transform 1 0 22908 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1174_
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _1175_
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1176_
timestamp 1649977179
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1649977179
transform 1 0 18124 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1649977179
transform 1 0 1472 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1649977179
transform -1 0 28796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1649977179
transform 1 0 2024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1649977179
transform -1 0 28796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1649977179
transform -1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1649977179
transform 1 0 2668 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1649977179
transform -1 0 28796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1649977179
transform -1 0 28796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input12
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 28520 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input14
timestamp 1649977179
transform 1 0 1748 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1649977179
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input16
timestamp 1649977179
transform 1 0 15548 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 1472 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform -1 0 28796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1649977179
transform -1 0 28796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1649977179
transform 1 0 24564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1649977179
transform -1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform -1 0 28796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform -1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1649977179
transform -1 0 28796 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1649977179
transform 1 0 21988 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input30
timestamp 1649977179
transform 1 0 7176 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input31
timestamp 1649977179
transform 1 0 14076 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input32
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input35
timestamp 1649977179
transform 1 0 1748 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1649977179
transform 1 0 20056 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input37
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform 1 0 27692 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform -1 0 10764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform 1 0 28428 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1649977179
transform 1 0 27692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1649977179
transform 1 0 11684 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1649977179
transform 1 0 28428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1649977179
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform 1 0 28428 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform -1 0 5612 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform 1 0 9108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform -1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform 1 0 28428 0 -1 14144
box -38 -48 406 592
<< labels >>
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 i_carry
port 0 nsew signal input
flabel metal2 s 18050 31965 18106 32765 0 FreeSans 224 90 0 0 i_l[0]
port 1 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 i_l[10]
port 2 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 i_l[11]
port 3 nsew signal input
flabel metal3 s 29821 9528 30621 9648 0 FreeSans 480 0 0 0 i_l[12]
port 4 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 i_l[13]
port 5 nsew signal input
flabel metal3 s 29821 7488 30621 7608 0 FreeSans 480 0 0 0 i_l[14]
port 6 nsew signal input
flabel metal3 s 29821 25848 30621 25968 0 FreeSans 480 0 0 0 i_l[15]
port 7 nsew signal input
flabel metal2 s 2594 31965 2650 32765 0 FreeSans 224 90 0 0 i_l[1]
port 8 nsew signal input
flabel metal3 s 29821 5448 30621 5568 0 FreeSans 480 0 0 0 i_l[2]
port 9 nsew signal input
flabel metal3 s 29821 21088 30621 21208 0 FreeSans 480 0 0 0 i_l[3]
port 10 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 i_l[4]
port 11 nsew signal input
flabel metal3 s 29821 19048 30621 19168 0 FreeSans 480 0 0 0 i_l[5]
port 12 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 i_l[6]
port 13 nsew signal input
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 i_l[7]
port 14 nsew signal input
flabel metal2 s 15474 31965 15530 32765 0 FreeSans 224 90 0 0 i_l[8]
port 15 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 i_l[9]
port 16 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 i_mode[0]
port 17 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 i_mode[1]
port 18 nsew signal input
flabel metal3 s 29821 27888 30621 28008 0 FreeSans 480 0 0 0 i_mode[2]
port 19 nsew signal input
flabel metal3 s 29821 16328 30621 16448 0 FreeSans 480 0 0 0 i_mode[3]
port 20 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 i_r[0]
port 21 nsew signal input
flabel metal2 s 24490 31965 24546 32765 0 FreeSans 224 90 0 0 i_r[10]
port 22 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 i_r[11]
port 23 nsew signal input
flabel metal3 s 29821 688 30621 808 0 FreeSans 480 0 0 0 i_r[12]
port 24 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 i_r[13]
port 25 nsew signal input
flabel metal3 s 29821 2728 30621 2848 0 FreeSans 480 0 0 0 i_r[14]
port 26 nsew signal input
flabel metal2 s 30286 31965 30342 32765 0 FreeSans 224 90 0 0 i_r[15]
port 27 nsew signal input
flabel metal2 s 21914 31965 21970 32765 0 FreeSans 224 90 0 0 i_r[1]
port 28 nsew signal input
flabel metal2 s 7102 31965 7158 32765 0 FreeSans 224 90 0 0 i_r[2]
port 29 nsew signal input
flabel metal2 s 13542 31965 13598 32765 0 FreeSans 224 90 0 0 i_r[3]
port 30 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 i_r[4]
port 31 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 i_r[5]
port 32 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 i_r[6]
port 33 nsew signal input
flabel metal2 s 662 31965 718 32765 0 FreeSans 224 90 0 0 i_r[7]
port 34 nsew signal input
flabel metal2 s 19982 31965 20038 32765 0 FreeSans 224 90 0 0 i_r[8]
port 35 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 i_r[9]
port 36 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 o_flags[0]
port 37 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 o_flags[1]
port 38 nsew signal tristate
flabel metal3 s 29821 29928 30621 30048 0 FreeSans 480 0 0 0 o_flags[2]
port 39 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 o_flags[3]
port 40 nsew signal tristate
flabel metal3 s 29821 23128 30621 23248 0 FreeSans 480 0 0 0 o_flags[4]
port 41 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 o_out[0]
port 42 nsew signal tristate
flabel metal2 s 11610 31965 11666 32765 0 FreeSans 224 90 0 0 o_out[10]
port 43 nsew signal tristate
flabel metal3 s 29821 12248 30621 12368 0 FreeSans 480 0 0 0 o_out[11]
port 44 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 o_out[12]
port 45 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 o_out[13]
port 46 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 o_out[14]
port 47 nsew signal tristate
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 o_out[15]
port 48 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 o_out[1]
port 49 nsew signal tristate
flabel metal2 s 28354 31965 28410 32765 0 FreeSans 224 90 0 0 o_out[2]
port 50 nsew signal tristate
flabel metal2 s 26422 31965 26478 32765 0 FreeSans 224 90 0 0 o_out[3]
port 51 nsew signal tristate
flabel metal2 s 5170 31965 5226 32765 0 FreeSans 224 90 0 0 o_out[4]
port 52 nsew signal tristate
flabel metal2 s 9034 31965 9090 32765 0 FreeSans 224 90 0 0 o_out[5]
port 53 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 o_out[6]
port 54 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 o_out[7]
port 55 nsew signal tristate
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 o_out[8]
port 56 nsew signal tristate
flabel metal3 s 29821 14288 30621 14408 0 FreeSans 480 0 0 0 o_out[9]
port 57 nsew signal tristate
flabel metal4 s 4486 2128 4806 30512 0 FreeSans 1920 90 0 0 vccd1
port 58 nsew power bidirectional
flabel metal4 s 11570 2128 11890 30512 0 FreeSans 1920 90 0 0 vccd1
port 58 nsew power bidirectional
flabel metal4 s 18654 2128 18974 30512 0 FreeSans 1920 90 0 0 vccd1
port 58 nsew power bidirectional
flabel metal4 s 25738 2128 26058 30512 0 FreeSans 1920 90 0 0 vccd1
port 58 nsew power bidirectional
flabel metal4 s 8028 2128 8348 30512 0 FreeSans 1920 90 0 0 vssd1
port 59 nsew ground bidirectional
flabel metal4 s 15112 2128 15432 30512 0 FreeSans 1920 90 0 0 vssd1
port 59 nsew ground bidirectional
flabel metal4 s 22196 2128 22516 30512 0 FreeSans 1920 90 0 0 vssd1
port 59 nsew ground bidirectional
flabel metal4 s 29280 2128 29600 30512 0 FreeSans 1920 90 0 0 vssd1
port 59 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30621 32765
<< end >>
