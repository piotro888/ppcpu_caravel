VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core1
  CLASS BLOCK ;
  FOREIGN core1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 1000.000 ;
  PIN dbg_pc[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 996.000 54.320 1000.000 ;
    END
  END dbg_pc[0]
  PIN dbg_pc[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 318.080 996.000 318.640 1000.000 ;
    END
  END dbg_pc[10]
  PIN dbg_pc[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 996.000 341.040 1000.000 ;
    END
  END dbg_pc[11]
  PIN dbg_pc[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 996.000 363.440 1000.000 ;
    END
  END dbg_pc[12]
  PIN dbg_pc[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 385.280 996.000 385.840 1000.000 ;
    END
  END dbg_pc[13]
  PIN dbg_pc[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 407.680 996.000 408.240 1000.000 ;
    END
  END dbg_pc[14]
  PIN dbg_pc[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 996.000 430.640 1000.000 ;
    END
  END dbg_pc[15]
  PIN dbg_pc[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 996.000 83.440 1000.000 ;
    END
  END dbg_pc[1]
  PIN dbg_pc[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 996.000 112.560 1000.000 ;
    END
  END dbg_pc[2]
  PIN dbg_pc[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 996.000 139.440 1000.000 ;
    END
  END dbg_pc[3]
  PIN dbg_pc[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 996.000 166.320 1000.000 ;
    END
  END dbg_pc[4]
  PIN dbg_pc[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 996.000 193.200 1000.000 ;
    END
  END dbg_pc[5]
  PIN dbg_pc[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 996.000 220.080 1000.000 ;
    END
  END dbg_pc[6]
  PIN dbg_pc[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 996.000 246.960 1000.000 ;
    END
  END dbg_pc[7]
  PIN dbg_pc[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 996.000 273.840 1000.000 ;
    END
  END dbg_pc[8]
  PIN dbg_pc[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 996.000 296.240 1000.000 ;
    END
  END dbg_pc[9]
  PIN dbg_r0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 996.000 56.560 1000.000 ;
    END
  END dbg_r0[0]
  PIN dbg_r0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 996.000 320.880 1000.000 ;
    END
  END dbg_r0[10]
  PIN dbg_r0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 996.000 343.280 1000.000 ;
    END
  END dbg_r0[11]
  PIN dbg_r0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 996.000 365.680 1000.000 ;
    END
  END dbg_r0[12]
  PIN dbg_r0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 996.000 388.080 1000.000 ;
    END
  END dbg_r0[13]
  PIN dbg_r0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 996.000 410.480 1000.000 ;
    END
  END dbg_r0[14]
  PIN dbg_r0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 996.000 432.880 1000.000 ;
    END
  END dbg_r0[15]
  PIN dbg_r0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 996.000 85.680 1000.000 ;
    END
  END dbg_r0[1]
  PIN dbg_r0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 996.000 114.800 1000.000 ;
    END
  END dbg_r0[2]
  PIN dbg_r0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 996.000 141.680 1000.000 ;
    END
  END dbg_r0[3]
  PIN dbg_r0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 996.000 168.560 1000.000 ;
    END
  END dbg_r0[4]
  PIN dbg_r0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 996.000 195.440 1000.000 ;
    END
  END dbg_r0[5]
  PIN dbg_r0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 996.000 222.320 1000.000 ;
    END
  END dbg_r0[6]
  PIN dbg_r0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 996.000 249.200 1000.000 ;
    END
  END dbg_r0[7]
  PIN dbg_r0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 996.000 276.080 1000.000 ;
    END
  END dbg_r0[8]
  PIN dbg_r0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 996.000 298.480 1000.000 ;
    END
  END dbg_r0[9]
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 996.000 14.000 1000.000 ;
    END
  END i_clk
  PIN i_core_int_sreg[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 996.000 58.800 1000.000 ;
    END
  END i_core_int_sreg[0]
  PIN i_core_int_sreg[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 996.000 323.120 1000.000 ;
    END
  END i_core_int_sreg[10]
  PIN i_core_int_sreg[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 344.960 996.000 345.520 1000.000 ;
    END
  END i_core_int_sreg[11]
  PIN i_core_int_sreg[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 996.000 367.920 1000.000 ;
    END
  END i_core_int_sreg[12]
  PIN i_core_int_sreg[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 996.000 390.320 1000.000 ;
    END
  END i_core_int_sreg[13]
  PIN i_core_int_sreg[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 412.160 996.000 412.720 1000.000 ;
    END
  END i_core_int_sreg[14]
  PIN i_core_int_sreg[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 996.000 435.120 1000.000 ;
    END
  END i_core_int_sreg[15]
  PIN i_core_int_sreg[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 996.000 87.920 1000.000 ;
    END
  END i_core_int_sreg[1]
  PIN i_core_int_sreg[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 996.000 117.040 1000.000 ;
    END
  END i_core_int_sreg[2]
  PIN i_core_int_sreg[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 996.000 143.920 1000.000 ;
    END
  END i_core_int_sreg[3]
  PIN i_core_int_sreg[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 996.000 170.800 1000.000 ;
    END
  END i_core_int_sreg[4]
  PIN i_core_int_sreg[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 996.000 197.680 1000.000 ;
    END
  END i_core_int_sreg[5]
  PIN i_core_int_sreg[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 996.000 224.560 1000.000 ;
    END
  END i_core_int_sreg[6]
  PIN i_core_int_sreg[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 250.880 996.000 251.440 1000.000 ;
    END
  END i_core_int_sreg[7]
  PIN i_core_int_sreg[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 996.000 278.320 1000.000 ;
    END
  END i_core_int_sreg[8]
  PIN i_core_int_sreg[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 300.160 996.000 300.720 1000.000 ;
    END
  END i_core_int_sreg[9]
  PIN i_disable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 996.000 16.240 1000.000 ;
    END
  END i_disable
  PIN i_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 17.920 996.000 18.480 1000.000 ;
    END
  END i_irq
  PIN i_mc_core_int
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 996.000 20.720 1000.000 ;
    END
  END i_mc_core_int
  PIN i_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 996.000 22.960 1000.000 ;
    END
  END i_mem_ack
  PIN i_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 996.000 61.040 1000.000 ;
    END
  END i_mem_data[0]
  PIN i_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 996.000 325.360 1000.000 ;
    END
  END i_mem_data[10]
  PIN i_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 996.000 347.760 1000.000 ;
    END
  END i_mem_data[11]
  PIN i_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 996.000 370.160 1000.000 ;
    END
  END i_mem_data[12]
  PIN i_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 996.000 392.560 1000.000 ;
    END
  END i_mem_data[13]
  PIN i_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 996.000 414.960 1000.000 ;
    END
  END i_mem_data[14]
  PIN i_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 996.000 437.360 1000.000 ;
    END
  END i_mem_data[15]
  PIN i_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 996.000 90.160 1000.000 ;
    END
  END i_mem_data[1]
  PIN i_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 996.000 119.280 1000.000 ;
    END
  END i_mem_data[2]
  PIN i_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 996.000 146.160 1000.000 ;
    END
  END i_mem_data[3]
  PIN i_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 996.000 173.040 1000.000 ;
    END
  END i_mem_data[4]
  PIN i_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 996.000 199.920 1000.000 ;
    END
  END i_mem_data[5]
  PIN i_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 996.000 226.800 1000.000 ;
    END
  END i_mem_data[6]
  PIN i_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 996.000 253.680 1000.000 ;
    END
  END i_mem_data[7]
  PIN i_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 996.000 280.560 1000.000 ;
    END
  END i_mem_data[8]
  PIN i_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 996.000 302.960 1000.000 ;
    END
  END i_mem_data[9]
  PIN i_mem_exception
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 996.000 25.200 1000.000 ;
    END
  END i_mem_exception
  PIN i_req_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 996.000 63.280 1000.000 ;
    END
  END i_req_data[0]
  PIN i_req_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 327.040 996.000 327.600 1000.000 ;
    END
  END i_req_data[10]
  PIN i_req_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 996.000 350.000 1000.000 ;
    END
  END i_req_data[11]
  PIN i_req_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 371.840 996.000 372.400 1000.000 ;
    END
  END i_req_data[12]
  PIN i_req_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 996.000 394.800 1000.000 ;
    END
  END i_req_data[13]
  PIN i_req_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 996.000 417.200 1000.000 ;
    END
  END i_req_data[14]
  PIN i_req_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.040 996.000 439.600 1000.000 ;
    END
  END i_req_data[15]
  PIN i_req_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 452.480 996.000 453.040 1000.000 ;
    END
  END i_req_data[16]
  PIN i_req_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 996.000 455.280 1000.000 ;
    END
  END i_req_data[17]
  PIN i_req_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 996.000 457.520 1000.000 ;
    END
  END i_req_data[18]
  PIN i_req_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 996.000 459.760 1000.000 ;
    END
  END i_req_data[19]
  PIN i_req_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 996.000 92.400 1000.000 ;
    END
  END i_req_data[1]
  PIN i_req_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 996.000 462.000 1000.000 ;
    END
  END i_req_data[20]
  PIN i_req_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 996.000 464.240 1000.000 ;
    END
  END i_req_data[21]
  PIN i_req_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 465.920 996.000 466.480 1000.000 ;
    END
  END i_req_data[22]
  PIN i_req_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 996.000 468.720 1000.000 ;
    END
  END i_req_data[23]
  PIN i_req_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 996.000 470.960 1000.000 ;
    END
  END i_req_data[24]
  PIN i_req_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 472.640 996.000 473.200 1000.000 ;
    END
  END i_req_data[25]
  PIN i_req_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 474.880 996.000 475.440 1000.000 ;
    END
  END i_req_data[26]
  PIN i_req_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 996.000 477.680 1000.000 ;
    END
  END i_req_data[27]
  PIN i_req_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 479.360 996.000 479.920 1000.000 ;
    END
  END i_req_data[28]
  PIN i_req_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 996.000 482.160 1000.000 ;
    END
  END i_req_data[29]
  PIN i_req_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 996.000 121.520 1000.000 ;
    END
  END i_req_data[2]
  PIN i_req_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 996.000 484.400 1000.000 ;
    END
  END i_req_data[30]
  PIN i_req_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 486.080 996.000 486.640 1000.000 ;
    END
  END i_req_data[31]
  PIN i_req_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 996.000 148.400 1000.000 ;
    END
  END i_req_data[3]
  PIN i_req_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 996.000 175.280 1000.000 ;
    END
  END i_req_data[4]
  PIN i_req_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 996.000 202.160 1000.000 ;
    END
  END i_req_data[5]
  PIN i_req_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 996.000 229.040 1000.000 ;
    END
  END i_req_data[6]
  PIN i_req_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 996.000 255.920 1000.000 ;
    END
  END i_req_data[7]
  PIN i_req_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 996.000 282.800 1000.000 ;
    END
  END i_req_data[8]
  PIN i_req_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 304.640 996.000 305.200 1000.000 ;
    END
  END i_req_data[9]
  PIN i_req_data_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 996.000 27.440 1000.000 ;
    END
  END i_req_data_valid
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 996.000 29.680 1000.000 ;
    END
  END i_rst
  PIN o_c_data_page
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 996.000 31.920 1000.000 ;
    END
  END o_c_data_page
  PIN o_c_instr_long
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 996.000 34.160 1000.000 ;
    END
  END o_c_instr_long
  PIN o_c_instr_page
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 996.000 36.400 1000.000 ;
    END
  END o_c_instr_page
  PIN o_icache_flush
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 996.000 38.640 1000.000 ;
    END
  END o_icache_flush
  PIN o_instr_long_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 996.000 65.520 1000.000 ;
    END
  END o_instr_long_addr[0]
  PIN o_instr_long_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 996.000 94.640 1000.000 ;
    END
  END o_instr_long_addr[1]
  PIN o_instr_long_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 996.000 123.760 1000.000 ;
    END
  END o_instr_long_addr[2]
  PIN o_instr_long_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 996.000 150.640 1000.000 ;
    END
  END o_instr_long_addr[3]
  PIN o_instr_long_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 996.000 177.520 1000.000 ;
    END
  END o_instr_long_addr[4]
  PIN o_instr_long_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 996.000 204.400 1000.000 ;
    END
  END o_instr_long_addr[5]
  PIN o_instr_long_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 996.000 231.280 1000.000 ;
    END
  END o_instr_long_addr[6]
  PIN o_instr_long_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 996.000 258.160 1000.000 ;
    END
  END o_instr_long_addr[7]
  PIN o_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 996.000 67.760 1000.000 ;
    END
  END o_mem_addr[0]
  PIN o_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 996.000 329.840 1000.000 ;
    END
  END o_mem_addr[10]
  PIN o_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 996.000 352.240 1000.000 ;
    END
  END o_mem_addr[11]
  PIN o_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 996.000 374.640 1000.000 ;
    END
  END o_mem_addr[12]
  PIN o_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 996.000 397.040 1000.000 ;
    END
  END o_mem_addr[13]
  PIN o_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 996.000 419.440 1000.000 ;
    END
  END o_mem_addr[14]
  PIN o_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 996.000 441.840 1000.000 ;
    END
  END o_mem_addr[15]
  PIN o_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 996.000 96.880 1000.000 ;
    END
  END o_mem_addr[1]
  PIN o_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 996.000 126.000 1000.000 ;
    END
  END o_mem_addr[2]
  PIN o_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 996.000 152.880 1000.000 ;
    END
  END o_mem_addr[3]
  PIN o_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 996.000 179.760 1000.000 ;
    END
  END o_mem_addr[4]
  PIN o_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 996.000 206.640 1000.000 ;
    END
  END o_mem_addr[5]
  PIN o_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 232.960 996.000 233.520 1000.000 ;
    END
  END o_mem_addr[6]
  PIN o_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 996.000 260.400 1000.000 ;
    END
  END o_mem_addr[7]
  PIN o_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 996.000 285.040 1000.000 ;
    END
  END o_mem_addr[8]
  PIN o_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 996.000 307.440 1000.000 ;
    END
  END o_mem_addr[9]
  PIN o_mem_addr_high[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 996.000 70.000 1000.000 ;
    END
  END o_mem_addr_high[0]
  PIN o_mem_addr_high[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 996.000 99.120 1000.000 ;
    END
  END o_mem_addr_high[1]
  PIN o_mem_addr_high[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 996.000 128.240 1000.000 ;
    END
  END o_mem_addr_high[2]
  PIN o_mem_addr_high[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 996.000 155.120 1000.000 ;
    END
  END o_mem_addr_high[3]
  PIN o_mem_addr_high[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 996.000 182.000 1000.000 ;
    END
  END o_mem_addr_high[4]
  PIN o_mem_addr_high[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 996.000 208.880 1000.000 ;
    END
  END o_mem_addr_high[5]
  PIN o_mem_addr_high[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 996.000 235.760 1000.000 ;
    END
  END o_mem_addr_high[6]
  PIN o_mem_addr_high[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 996.000 262.640 1000.000 ;
    END
  END o_mem_addr_high[7]
  PIN o_mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 996.000 72.240 1000.000 ;
    END
  END o_mem_data[0]
  PIN o_mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 331.520 996.000 332.080 1000.000 ;
    END
  END o_mem_data[10]
  PIN o_mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 996.000 354.480 1000.000 ;
    END
  END o_mem_data[11]
  PIN o_mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 996.000 376.880 1000.000 ;
    END
  END o_mem_data[12]
  PIN o_mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 996.000 399.280 1000.000 ;
    END
  END o_mem_data[13]
  PIN o_mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 996.000 421.680 1000.000 ;
    END
  END o_mem_data[14]
  PIN o_mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 996.000 444.080 1000.000 ;
    END
  END o_mem_data[15]
  PIN o_mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 996.000 101.360 1000.000 ;
    END
  END o_mem_data[1]
  PIN o_mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 996.000 130.480 1000.000 ;
    END
  END o_mem_data[2]
  PIN o_mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 996.000 157.360 1000.000 ;
    END
  END o_mem_data[3]
  PIN o_mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 996.000 184.240 1000.000 ;
    END
  END o_mem_data[4]
  PIN o_mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 996.000 211.120 1000.000 ;
    END
  END o_mem_data[5]
  PIN o_mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 996.000 238.000 1000.000 ;
    END
  END o_mem_data[6]
  PIN o_mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 264.320 996.000 264.880 1000.000 ;
    END
  END o_mem_data[7]
  PIN o_mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 996.000 287.280 1000.000 ;
    END
  END o_mem_data[8]
  PIN o_mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 996.000 309.680 1000.000 ;
    END
  END o_mem_data[9]
  PIN o_mem_long
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 996.000 40.880 1000.000 ;
    END
  END o_mem_long
  PIN o_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 996.000 43.120 1000.000 ;
    END
  END o_mem_req
  PIN o_mem_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 996.000 74.480 1000.000 ;
    END
  END o_mem_sel[0]
  PIN o_mem_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 996.000 103.600 1000.000 ;
    END
  END o_mem_sel[1]
  PIN o_mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 996.000 45.360 1000.000 ;
    END
  END o_mem_we
  PIN o_req_active
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 996.000 47.600 1000.000 ;
    END
  END o_req_active
  PIN o_req_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 996.000 76.720 1000.000 ;
    END
  END o_req_addr[0]
  PIN o_req_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 996.000 334.320 1000.000 ;
    END
  END o_req_addr[10]
  PIN o_req_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 996.000 356.720 1000.000 ;
    END
  END o_req_addr[11]
  PIN o_req_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 996.000 379.120 1000.000 ;
    END
  END o_req_addr[12]
  PIN o_req_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 996.000 401.520 1000.000 ;
    END
  END o_req_addr[13]
  PIN o_req_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 996.000 423.920 1000.000 ;
    END
  END o_req_addr[14]
  PIN o_req_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 996.000 446.320 1000.000 ;
    END
  END o_req_addr[15]
  PIN o_req_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 996.000 105.840 1000.000 ;
    END
  END o_req_addr[1]
  PIN o_req_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 996.000 132.720 1000.000 ;
    END
  END o_req_addr[2]
  PIN o_req_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 996.000 159.600 1000.000 ;
    END
  END o_req_addr[3]
  PIN o_req_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 996.000 186.480 1000.000 ;
    END
  END o_req_addr[4]
  PIN o_req_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 996.000 213.360 1000.000 ;
    END
  END o_req_addr[5]
  PIN o_req_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 996.000 240.240 1000.000 ;
    END
  END o_req_addr[6]
  PIN o_req_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 996.000 267.120 1000.000 ;
    END
  END o_req_addr[7]
  PIN o_req_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 996.000 289.520 1000.000 ;
    END
  END o_req_addr[8]
  PIN o_req_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 996.000 311.920 1000.000 ;
    END
  END o_req_addr[9]
  PIN o_req_ppl_submit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 996.000 49.840 1000.000 ;
    END
  END o_req_ppl_submit
  PIN sr_bus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 996.000 78.960 1000.000 ;
    END
  END sr_bus_addr[0]
  PIN sr_bus_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 996.000 336.560 1000.000 ;
    END
  END sr_bus_addr[10]
  PIN sr_bus_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 358.400 996.000 358.960 1000.000 ;
    END
  END sr_bus_addr[11]
  PIN sr_bus_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 996.000 381.360 1000.000 ;
    END
  END sr_bus_addr[12]
  PIN sr_bus_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 996.000 403.760 1000.000 ;
    END
  END sr_bus_addr[13]
  PIN sr_bus_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 425.600 996.000 426.160 1000.000 ;
    END
  END sr_bus_addr[14]
  PIN sr_bus_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 996.000 448.560 1000.000 ;
    END
  END sr_bus_addr[15]
  PIN sr_bus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 996.000 108.080 1000.000 ;
    END
  END sr_bus_addr[1]
  PIN sr_bus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 996.000 134.960 1000.000 ;
    END
  END sr_bus_addr[2]
  PIN sr_bus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 996.000 161.840 1000.000 ;
    END
  END sr_bus_addr[3]
  PIN sr_bus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 996.000 188.720 1000.000 ;
    END
  END sr_bus_addr[4]
  PIN sr_bus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 996.000 215.600 1000.000 ;
    END
  END sr_bus_addr[5]
  PIN sr_bus_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 996.000 242.480 1000.000 ;
    END
  END sr_bus_addr[6]
  PIN sr_bus_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 996.000 269.360 1000.000 ;
    END
  END sr_bus_addr[7]
  PIN sr_bus_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 996.000 291.760 1000.000 ;
    END
  END sr_bus_addr[8]
  PIN sr_bus_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 996.000 314.160 1000.000 ;
    END
  END sr_bus_addr[9]
  PIN sr_bus_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 996.000 81.200 1000.000 ;
    END
  END sr_bus_data_o[0]
  PIN sr_bus_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 996.000 338.800 1000.000 ;
    END
  END sr_bus_data_o[10]
  PIN sr_bus_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 996.000 361.200 1000.000 ;
    END
  END sr_bus_data_o[11]
  PIN sr_bus_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 996.000 383.600 1000.000 ;
    END
  END sr_bus_data_o[12]
  PIN sr_bus_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 996.000 406.000 1000.000 ;
    END
  END sr_bus_data_o[13]
  PIN sr_bus_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 427.840 996.000 428.400 1000.000 ;
    END
  END sr_bus_data_o[14]
  PIN sr_bus_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 996.000 450.800 1000.000 ;
    END
  END sr_bus_data_o[15]
  PIN sr_bus_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 996.000 110.320 1000.000 ;
    END
  END sr_bus_data_o[1]
  PIN sr_bus_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 996.000 137.200 1000.000 ;
    END
  END sr_bus_data_o[2]
  PIN sr_bus_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 996.000 164.080 1000.000 ;
    END
  END sr_bus_data_o[3]
  PIN sr_bus_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 996.000 190.960 1000.000 ;
    END
  END sr_bus_data_o[4]
  PIN sr_bus_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 996.000 217.840 1000.000 ;
    END
  END sr_bus_data_o[5]
  PIN sr_bus_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 996.000 244.720 1000.000 ;
    END
  END sr_bus_data_o[6]
  PIN sr_bus_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 996.000 271.600 1000.000 ;
    END
  END sr_bus_data_o[7]
  PIN sr_bus_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 996.000 294.000 1000.000 ;
    END
  END sr_bus_data_o[8]
  PIN sr_bus_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 996.000 316.400 1000.000 ;
    END
  END sr_bus_data_o[9]
  PIN sr_bus_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 996.000 52.080 1000.000 ;
    END
  END sr_bus_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 984.220 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 984.220 ;
    END
  END vssd1
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 492.800 987.130 ;
      LAYER Metal2 ;
        RECT 4.620 995.700 13.140 996.000 ;
        RECT 14.300 995.700 15.380 996.000 ;
        RECT 16.540 995.700 17.620 996.000 ;
        RECT 18.780 995.700 19.860 996.000 ;
        RECT 21.020 995.700 22.100 996.000 ;
        RECT 23.260 995.700 24.340 996.000 ;
        RECT 25.500 995.700 26.580 996.000 ;
        RECT 27.740 995.700 28.820 996.000 ;
        RECT 29.980 995.700 31.060 996.000 ;
        RECT 32.220 995.700 33.300 996.000 ;
        RECT 34.460 995.700 35.540 996.000 ;
        RECT 36.700 995.700 37.780 996.000 ;
        RECT 38.940 995.700 40.020 996.000 ;
        RECT 41.180 995.700 42.260 996.000 ;
        RECT 43.420 995.700 44.500 996.000 ;
        RECT 45.660 995.700 46.740 996.000 ;
        RECT 47.900 995.700 48.980 996.000 ;
        RECT 50.140 995.700 51.220 996.000 ;
        RECT 52.380 995.700 53.460 996.000 ;
        RECT 54.620 995.700 55.700 996.000 ;
        RECT 56.860 995.700 57.940 996.000 ;
        RECT 59.100 995.700 60.180 996.000 ;
        RECT 61.340 995.700 62.420 996.000 ;
        RECT 63.580 995.700 64.660 996.000 ;
        RECT 65.820 995.700 66.900 996.000 ;
        RECT 68.060 995.700 69.140 996.000 ;
        RECT 70.300 995.700 71.380 996.000 ;
        RECT 72.540 995.700 73.620 996.000 ;
        RECT 74.780 995.700 75.860 996.000 ;
        RECT 77.020 995.700 78.100 996.000 ;
        RECT 79.260 995.700 80.340 996.000 ;
        RECT 81.500 995.700 82.580 996.000 ;
        RECT 83.740 995.700 84.820 996.000 ;
        RECT 85.980 995.700 87.060 996.000 ;
        RECT 88.220 995.700 89.300 996.000 ;
        RECT 90.460 995.700 91.540 996.000 ;
        RECT 92.700 995.700 93.780 996.000 ;
        RECT 94.940 995.700 96.020 996.000 ;
        RECT 97.180 995.700 98.260 996.000 ;
        RECT 99.420 995.700 100.500 996.000 ;
        RECT 101.660 995.700 102.740 996.000 ;
        RECT 103.900 995.700 104.980 996.000 ;
        RECT 106.140 995.700 107.220 996.000 ;
        RECT 108.380 995.700 109.460 996.000 ;
        RECT 110.620 995.700 111.700 996.000 ;
        RECT 112.860 995.700 113.940 996.000 ;
        RECT 115.100 995.700 116.180 996.000 ;
        RECT 117.340 995.700 118.420 996.000 ;
        RECT 119.580 995.700 120.660 996.000 ;
        RECT 121.820 995.700 122.900 996.000 ;
        RECT 124.060 995.700 125.140 996.000 ;
        RECT 126.300 995.700 127.380 996.000 ;
        RECT 128.540 995.700 129.620 996.000 ;
        RECT 130.780 995.700 131.860 996.000 ;
        RECT 133.020 995.700 134.100 996.000 ;
        RECT 135.260 995.700 136.340 996.000 ;
        RECT 137.500 995.700 138.580 996.000 ;
        RECT 139.740 995.700 140.820 996.000 ;
        RECT 141.980 995.700 143.060 996.000 ;
        RECT 144.220 995.700 145.300 996.000 ;
        RECT 146.460 995.700 147.540 996.000 ;
        RECT 148.700 995.700 149.780 996.000 ;
        RECT 150.940 995.700 152.020 996.000 ;
        RECT 153.180 995.700 154.260 996.000 ;
        RECT 155.420 995.700 156.500 996.000 ;
        RECT 157.660 995.700 158.740 996.000 ;
        RECT 159.900 995.700 160.980 996.000 ;
        RECT 162.140 995.700 163.220 996.000 ;
        RECT 164.380 995.700 165.460 996.000 ;
        RECT 166.620 995.700 167.700 996.000 ;
        RECT 168.860 995.700 169.940 996.000 ;
        RECT 171.100 995.700 172.180 996.000 ;
        RECT 173.340 995.700 174.420 996.000 ;
        RECT 175.580 995.700 176.660 996.000 ;
        RECT 177.820 995.700 178.900 996.000 ;
        RECT 180.060 995.700 181.140 996.000 ;
        RECT 182.300 995.700 183.380 996.000 ;
        RECT 184.540 995.700 185.620 996.000 ;
        RECT 186.780 995.700 187.860 996.000 ;
        RECT 189.020 995.700 190.100 996.000 ;
        RECT 191.260 995.700 192.340 996.000 ;
        RECT 193.500 995.700 194.580 996.000 ;
        RECT 195.740 995.700 196.820 996.000 ;
        RECT 197.980 995.700 199.060 996.000 ;
        RECT 200.220 995.700 201.300 996.000 ;
        RECT 202.460 995.700 203.540 996.000 ;
        RECT 204.700 995.700 205.780 996.000 ;
        RECT 206.940 995.700 208.020 996.000 ;
        RECT 209.180 995.700 210.260 996.000 ;
        RECT 211.420 995.700 212.500 996.000 ;
        RECT 213.660 995.700 214.740 996.000 ;
        RECT 215.900 995.700 216.980 996.000 ;
        RECT 218.140 995.700 219.220 996.000 ;
        RECT 220.380 995.700 221.460 996.000 ;
        RECT 222.620 995.700 223.700 996.000 ;
        RECT 224.860 995.700 225.940 996.000 ;
        RECT 227.100 995.700 228.180 996.000 ;
        RECT 229.340 995.700 230.420 996.000 ;
        RECT 231.580 995.700 232.660 996.000 ;
        RECT 233.820 995.700 234.900 996.000 ;
        RECT 236.060 995.700 237.140 996.000 ;
        RECT 238.300 995.700 239.380 996.000 ;
        RECT 240.540 995.700 241.620 996.000 ;
        RECT 242.780 995.700 243.860 996.000 ;
        RECT 245.020 995.700 246.100 996.000 ;
        RECT 247.260 995.700 248.340 996.000 ;
        RECT 249.500 995.700 250.580 996.000 ;
        RECT 251.740 995.700 252.820 996.000 ;
        RECT 253.980 995.700 255.060 996.000 ;
        RECT 256.220 995.700 257.300 996.000 ;
        RECT 258.460 995.700 259.540 996.000 ;
        RECT 260.700 995.700 261.780 996.000 ;
        RECT 262.940 995.700 264.020 996.000 ;
        RECT 265.180 995.700 266.260 996.000 ;
        RECT 267.420 995.700 268.500 996.000 ;
        RECT 269.660 995.700 270.740 996.000 ;
        RECT 271.900 995.700 272.980 996.000 ;
        RECT 274.140 995.700 275.220 996.000 ;
        RECT 276.380 995.700 277.460 996.000 ;
        RECT 278.620 995.700 279.700 996.000 ;
        RECT 280.860 995.700 281.940 996.000 ;
        RECT 283.100 995.700 284.180 996.000 ;
        RECT 285.340 995.700 286.420 996.000 ;
        RECT 287.580 995.700 288.660 996.000 ;
        RECT 289.820 995.700 290.900 996.000 ;
        RECT 292.060 995.700 293.140 996.000 ;
        RECT 294.300 995.700 295.380 996.000 ;
        RECT 296.540 995.700 297.620 996.000 ;
        RECT 298.780 995.700 299.860 996.000 ;
        RECT 301.020 995.700 302.100 996.000 ;
        RECT 303.260 995.700 304.340 996.000 ;
        RECT 305.500 995.700 306.580 996.000 ;
        RECT 307.740 995.700 308.820 996.000 ;
        RECT 309.980 995.700 311.060 996.000 ;
        RECT 312.220 995.700 313.300 996.000 ;
        RECT 314.460 995.700 315.540 996.000 ;
        RECT 316.700 995.700 317.780 996.000 ;
        RECT 318.940 995.700 320.020 996.000 ;
        RECT 321.180 995.700 322.260 996.000 ;
        RECT 323.420 995.700 324.500 996.000 ;
        RECT 325.660 995.700 326.740 996.000 ;
        RECT 327.900 995.700 328.980 996.000 ;
        RECT 330.140 995.700 331.220 996.000 ;
        RECT 332.380 995.700 333.460 996.000 ;
        RECT 334.620 995.700 335.700 996.000 ;
        RECT 336.860 995.700 337.940 996.000 ;
        RECT 339.100 995.700 340.180 996.000 ;
        RECT 341.340 995.700 342.420 996.000 ;
        RECT 343.580 995.700 344.660 996.000 ;
        RECT 345.820 995.700 346.900 996.000 ;
        RECT 348.060 995.700 349.140 996.000 ;
        RECT 350.300 995.700 351.380 996.000 ;
        RECT 352.540 995.700 353.620 996.000 ;
        RECT 354.780 995.700 355.860 996.000 ;
        RECT 357.020 995.700 358.100 996.000 ;
        RECT 359.260 995.700 360.340 996.000 ;
        RECT 361.500 995.700 362.580 996.000 ;
        RECT 363.740 995.700 364.820 996.000 ;
        RECT 365.980 995.700 367.060 996.000 ;
        RECT 368.220 995.700 369.300 996.000 ;
        RECT 370.460 995.700 371.540 996.000 ;
        RECT 372.700 995.700 373.780 996.000 ;
        RECT 374.940 995.700 376.020 996.000 ;
        RECT 377.180 995.700 378.260 996.000 ;
        RECT 379.420 995.700 380.500 996.000 ;
        RECT 381.660 995.700 382.740 996.000 ;
        RECT 383.900 995.700 384.980 996.000 ;
        RECT 386.140 995.700 387.220 996.000 ;
        RECT 388.380 995.700 389.460 996.000 ;
        RECT 390.620 995.700 391.700 996.000 ;
        RECT 392.860 995.700 393.940 996.000 ;
        RECT 395.100 995.700 396.180 996.000 ;
        RECT 397.340 995.700 398.420 996.000 ;
        RECT 399.580 995.700 400.660 996.000 ;
        RECT 401.820 995.700 402.900 996.000 ;
        RECT 404.060 995.700 405.140 996.000 ;
        RECT 406.300 995.700 407.380 996.000 ;
        RECT 408.540 995.700 409.620 996.000 ;
        RECT 410.780 995.700 411.860 996.000 ;
        RECT 413.020 995.700 414.100 996.000 ;
        RECT 415.260 995.700 416.340 996.000 ;
        RECT 417.500 995.700 418.580 996.000 ;
        RECT 419.740 995.700 420.820 996.000 ;
        RECT 421.980 995.700 423.060 996.000 ;
        RECT 424.220 995.700 425.300 996.000 ;
        RECT 426.460 995.700 427.540 996.000 ;
        RECT 428.700 995.700 429.780 996.000 ;
        RECT 430.940 995.700 432.020 996.000 ;
        RECT 433.180 995.700 434.260 996.000 ;
        RECT 435.420 995.700 436.500 996.000 ;
        RECT 437.660 995.700 438.740 996.000 ;
        RECT 439.900 995.700 440.980 996.000 ;
        RECT 442.140 995.700 443.220 996.000 ;
        RECT 444.380 995.700 445.460 996.000 ;
        RECT 446.620 995.700 447.700 996.000 ;
        RECT 448.860 995.700 449.940 996.000 ;
        RECT 451.100 995.700 452.180 996.000 ;
        RECT 453.340 995.700 454.420 996.000 ;
        RECT 455.580 995.700 456.660 996.000 ;
        RECT 457.820 995.700 458.900 996.000 ;
        RECT 460.060 995.700 461.140 996.000 ;
        RECT 462.300 995.700 463.380 996.000 ;
        RECT 464.540 995.700 465.620 996.000 ;
        RECT 466.780 995.700 467.860 996.000 ;
        RECT 469.020 995.700 470.100 996.000 ;
        RECT 471.260 995.700 472.340 996.000 ;
        RECT 473.500 995.700 474.580 996.000 ;
        RECT 475.740 995.700 476.820 996.000 ;
        RECT 477.980 995.700 479.060 996.000 ;
        RECT 480.220 995.700 481.300 996.000 ;
        RECT 482.460 995.700 483.540 996.000 ;
        RECT 484.700 995.700 485.780 996.000 ;
        RECT 486.940 995.700 492.100 996.000 ;
        RECT 4.620 15.490 492.100 995.700 ;
      LAYER Metal3 ;
        RECT 4.570 15.540 492.150 985.460 ;
      LAYER Metal4 ;
        RECT 24.220 30.330 98.740 981.590 ;
        RECT 100.940 30.330 175.540 981.590 ;
        RECT 177.740 30.330 252.340 981.590 ;
        RECT 254.540 30.330 329.140 981.590 ;
        RECT 331.340 30.330 405.940 981.590 ;
        RECT 408.140 30.330 482.740 981.590 ;
        RECT 484.940 30.330 487.060 981.590 ;
  END
END core1
END LIBRARY

