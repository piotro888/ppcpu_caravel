module int_ram (i_clk,
    i_we,
    vccd1,
    vssd1,
    i_addr,
    i_data,
    o_data);
 input i_clk;
 input i_we;
 input vccd1;
 input vssd1;
 input [5:0] i_addr;
 input [15:0] i_data;
 output [15:0] o_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire clknet_0_i_clk;
 wire clknet_3_0_0_i_clk;
 wire clknet_3_1_0_i_clk;
 wire clknet_3_2_0_i_clk;
 wire clknet_3_3_0_i_clk;
 wire clknet_3_4_0_i_clk;
 wire clknet_3_5_0_i_clk;
 wire clknet_3_6_0_i_clk;
 wire clknet_3_7_0_i_clk;
 wire clknet_4_0__leaf_i_clk;
 wire clknet_4_10__leaf_i_clk;
 wire clknet_4_11__leaf_i_clk;
 wire clknet_4_12__leaf_i_clk;
 wire clknet_4_13__leaf_i_clk;
 wire clknet_4_14__leaf_i_clk;
 wire clknet_4_15__leaf_i_clk;
 wire clknet_4_1__leaf_i_clk;
 wire clknet_4_2__leaf_i_clk;
 wire clknet_4_3__leaf_i_clk;
 wire clknet_4_4__leaf_i_clk;
 wire clknet_4_5__leaf_i_clk;
 wire clknet_4_6__leaf_i_clk;
 wire clknet_4_7__leaf_i_clk;
 wire clknet_4_8__leaf_i_clk;
 wire clknet_4_9__leaf_i_clk;
 wire clknet_leaf_0_i_clk;
 wire clknet_leaf_100_i_clk;
 wire clknet_leaf_101_i_clk;
 wire clknet_leaf_102_i_clk;
 wire clknet_leaf_103_i_clk;
 wire clknet_leaf_104_i_clk;
 wire clknet_leaf_105_i_clk;
 wire clknet_leaf_106_i_clk;
 wire clknet_leaf_107_i_clk;
 wire clknet_leaf_108_i_clk;
 wire clknet_leaf_109_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_110_i_clk;
 wire clknet_leaf_111_i_clk;
 wire clknet_leaf_112_i_clk;
 wire clknet_leaf_113_i_clk;
 wire clknet_leaf_114_i_clk;
 wire clknet_leaf_115_i_clk;
 wire clknet_leaf_116_i_clk;
 wire clknet_leaf_117_i_clk;
 wire clknet_leaf_118_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_52_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_62_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_65_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_67_i_clk;
 wire clknet_leaf_68_i_clk;
 wire clknet_leaf_69_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_70_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_72_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_75_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_79_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_80_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_82_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_86_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_90_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_94_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_leaf_96_i_clk;
 wire clknet_leaf_97_i_clk;
 wire clknet_leaf_98_i_clk;
 wire clknet_leaf_99_i_clk;
 wire clknet_leaf_9_i_clk;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[16][0] ;
 wire \mem[16][10] ;
 wire \mem[16][11] ;
 wire \mem[16][12] ;
 wire \mem[16][13] ;
 wire \mem[16][14] ;
 wire \mem[16][15] ;
 wire \mem[16][1] ;
 wire \mem[16][2] ;
 wire \mem[16][3] ;
 wire \mem[16][4] ;
 wire \mem[16][5] ;
 wire \mem[16][6] ;
 wire \mem[16][7] ;
 wire \mem[16][8] ;
 wire \mem[16][9] ;
 wire \mem[17][0] ;
 wire \mem[17][10] ;
 wire \mem[17][11] ;
 wire \mem[17][12] ;
 wire \mem[17][13] ;
 wire \mem[17][14] ;
 wire \mem[17][15] ;
 wire \mem[17][1] ;
 wire \mem[17][2] ;
 wire \mem[17][3] ;
 wire \mem[17][4] ;
 wire \mem[17][5] ;
 wire \mem[17][6] ;
 wire \mem[17][7] ;
 wire \mem[17][8] ;
 wire \mem[17][9] ;
 wire \mem[18][0] ;
 wire \mem[18][10] ;
 wire \mem[18][11] ;
 wire \mem[18][12] ;
 wire \mem[18][13] ;
 wire \mem[18][14] ;
 wire \mem[18][15] ;
 wire \mem[18][1] ;
 wire \mem[18][2] ;
 wire \mem[18][3] ;
 wire \mem[18][4] ;
 wire \mem[18][5] ;
 wire \mem[18][6] ;
 wire \mem[18][7] ;
 wire \mem[18][8] ;
 wire \mem[18][9] ;
 wire \mem[19][0] ;
 wire \mem[19][10] ;
 wire \mem[19][11] ;
 wire \mem[19][12] ;
 wire \mem[19][13] ;
 wire \mem[19][14] ;
 wire \mem[19][15] ;
 wire \mem[19][1] ;
 wire \mem[19][2] ;
 wire \mem[19][3] ;
 wire \mem[19][4] ;
 wire \mem[19][5] ;
 wire \mem[19][6] ;
 wire \mem[19][7] ;
 wire \mem[19][8] ;
 wire \mem[19][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[20][0] ;
 wire \mem[20][10] ;
 wire \mem[20][11] ;
 wire \mem[20][12] ;
 wire \mem[20][13] ;
 wire \mem[20][14] ;
 wire \mem[20][15] ;
 wire \mem[20][1] ;
 wire \mem[20][2] ;
 wire \mem[20][3] ;
 wire \mem[20][4] ;
 wire \mem[20][5] ;
 wire \mem[20][6] ;
 wire \mem[20][7] ;
 wire \mem[20][8] ;
 wire \mem[20][9] ;
 wire \mem[21][0] ;
 wire \mem[21][10] ;
 wire \mem[21][11] ;
 wire \mem[21][12] ;
 wire \mem[21][13] ;
 wire \mem[21][14] ;
 wire \mem[21][15] ;
 wire \mem[21][1] ;
 wire \mem[21][2] ;
 wire \mem[21][3] ;
 wire \mem[21][4] ;
 wire \mem[21][5] ;
 wire \mem[21][6] ;
 wire \mem[21][7] ;
 wire \mem[21][8] ;
 wire \mem[21][9] ;
 wire \mem[22][0] ;
 wire \mem[22][10] ;
 wire \mem[22][11] ;
 wire \mem[22][12] ;
 wire \mem[22][13] ;
 wire \mem[22][14] ;
 wire \mem[22][15] ;
 wire \mem[22][1] ;
 wire \mem[22][2] ;
 wire \mem[22][3] ;
 wire \mem[22][4] ;
 wire \mem[22][5] ;
 wire \mem[22][6] ;
 wire \mem[22][7] ;
 wire \mem[22][8] ;
 wire \mem[22][9] ;
 wire \mem[23][0] ;
 wire \mem[23][10] ;
 wire \mem[23][11] ;
 wire \mem[23][12] ;
 wire \mem[23][13] ;
 wire \mem[23][14] ;
 wire \mem[23][15] ;
 wire \mem[23][1] ;
 wire \mem[23][2] ;
 wire \mem[23][3] ;
 wire \mem[23][4] ;
 wire \mem[23][5] ;
 wire \mem[23][6] ;
 wire \mem[23][7] ;
 wire \mem[23][8] ;
 wire \mem[23][9] ;
 wire \mem[24][0] ;
 wire \mem[24][10] ;
 wire \mem[24][11] ;
 wire \mem[24][12] ;
 wire \mem[24][13] ;
 wire \mem[24][14] ;
 wire \mem[24][15] ;
 wire \mem[24][1] ;
 wire \mem[24][2] ;
 wire \mem[24][3] ;
 wire \mem[24][4] ;
 wire \mem[24][5] ;
 wire \mem[24][6] ;
 wire \mem[24][7] ;
 wire \mem[24][8] ;
 wire \mem[24][9] ;
 wire \mem[25][0] ;
 wire \mem[25][10] ;
 wire \mem[25][11] ;
 wire \mem[25][12] ;
 wire \mem[25][13] ;
 wire \mem[25][14] ;
 wire \mem[25][15] ;
 wire \mem[25][1] ;
 wire \mem[25][2] ;
 wire \mem[25][3] ;
 wire \mem[25][4] ;
 wire \mem[25][5] ;
 wire \mem[25][6] ;
 wire \mem[25][7] ;
 wire \mem[25][8] ;
 wire \mem[25][9] ;
 wire \mem[26][0] ;
 wire \mem[26][10] ;
 wire \mem[26][11] ;
 wire \mem[26][12] ;
 wire \mem[26][13] ;
 wire \mem[26][14] ;
 wire \mem[26][15] ;
 wire \mem[26][1] ;
 wire \mem[26][2] ;
 wire \mem[26][3] ;
 wire \mem[26][4] ;
 wire \mem[26][5] ;
 wire \mem[26][6] ;
 wire \mem[26][7] ;
 wire \mem[26][8] ;
 wire \mem[26][9] ;
 wire \mem[27][0] ;
 wire \mem[27][10] ;
 wire \mem[27][11] ;
 wire \mem[27][12] ;
 wire \mem[27][13] ;
 wire \mem[27][14] ;
 wire \mem[27][15] ;
 wire \mem[27][1] ;
 wire \mem[27][2] ;
 wire \mem[27][3] ;
 wire \mem[27][4] ;
 wire \mem[27][5] ;
 wire \mem[27][6] ;
 wire \mem[27][7] ;
 wire \mem[27][8] ;
 wire \mem[27][9] ;
 wire \mem[28][0] ;
 wire \mem[28][10] ;
 wire \mem[28][11] ;
 wire \mem[28][12] ;
 wire \mem[28][13] ;
 wire \mem[28][14] ;
 wire \mem[28][15] ;
 wire \mem[28][1] ;
 wire \mem[28][2] ;
 wire \mem[28][3] ;
 wire \mem[28][4] ;
 wire \mem[28][5] ;
 wire \mem[28][6] ;
 wire \mem[28][7] ;
 wire \mem[28][8] ;
 wire \mem[28][9] ;
 wire \mem[29][0] ;
 wire \mem[29][10] ;
 wire \mem[29][11] ;
 wire \mem[29][12] ;
 wire \mem[29][13] ;
 wire \mem[29][14] ;
 wire \mem[29][15] ;
 wire \mem[29][1] ;
 wire \mem[29][2] ;
 wire \mem[29][3] ;
 wire \mem[29][4] ;
 wire \mem[29][5] ;
 wire \mem[29][6] ;
 wire \mem[29][7] ;
 wire \mem[29][8] ;
 wire \mem[29][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[30][0] ;
 wire \mem[30][10] ;
 wire \mem[30][11] ;
 wire \mem[30][12] ;
 wire \mem[30][13] ;
 wire \mem[30][14] ;
 wire \mem[30][15] ;
 wire \mem[30][1] ;
 wire \mem[30][2] ;
 wire \mem[30][3] ;
 wire \mem[30][4] ;
 wire \mem[30][5] ;
 wire \mem[30][6] ;
 wire \mem[30][7] ;
 wire \mem[30][8] ;
 wire \mem[30][9] ;
 wire \mem[31][0] ;
 wire \mem[31][10] ;
 wire \mem[31][11] ;
 wire \mem[31][12] ;
 wire \mem[31][13] ;
 wire \mem[31][14] ;
 wire \mem[31][15] ;
 wire \mem[31][1] ;
 wire \mem[31][2] ;
 wire \mem[31][3] ;
 wire \mem[31][4] ;
 wire \mem[31][5] ;
 wire \mem[31][6] ;
 wire \mem[31][7] ;
 wire \mem[31][8] ;
 wire \mem[31][9] ;
 wire \mem[32][0] ;
 wire \mem[32][10] ;
 wire \mem[32][11] ;
 wire \mem[32][12] ;
 wire \mem[32][13] ;
 wire \mem[32][14] ;
 wire \mem[32][15] ;
 wire \mem[32][1] ;
 wire \mem[32][2] ;
 wire \mem[32][3] ;
 wire \mem[32][4] ;
 wire \mem[32][5] ;
 wire \mem[32][6] ;
 wire \mem[32][7] ;
 wire \mem[32][8] ;
 wire \mem[32][9] ;
 wire \mem[33][0] ;
 wire \mem[33][10] ;
 wire \mem[33][11] ;
 wire \mem[33][12] ;
 wire \mem[33][13] ;
 wire \mem[33][14] ;
 wire \mem[33][15] ;
 wire \mem[33][1] ;
 wire \mem[33][2] ;
 wire \mem[33][3] ;
 wire \mem[33][4] ;
 wire \mem[33][5] ;
 wire \mem[33][6] ;
 wire \mem[33][7] ;
 wire \mem[33][8] ;
 wire \mem[33][9] ;
 wire \mem[34][0] ;
 wire \mem[34][10] ;
 wire \mem[34][11] ;
 wire \mem[34][12] ;
 wire \mem[34][13] ;
 wire \mem[34][14] ;
 wire \mem[34][15] ;
 wire \mem[34][1] ;
 wire \mem[34][2] ;
 wire \mem[34][3] ;
 wire \mem[34][4] ;
 wire \mem[34][5] ;
 wire \mem[34][6] ;
 wire \mem[34][7] ;
 wire \mem[34][8] ;
 wire \mem[34][9] ;
 wire \mem[35][0] ;
 wire \mem[35][10] ;
 wire \mem[35][11] ;
 wire \mem[35][12] ;
 wire \mem[35][13] ;
 wire \mem[35][14] ;
 wire \mem[35][15] ;
 wire \mem[35][1] ;
 wire \mem[35][2] ;
 wire \mem[35][3] ;
 wire \mem[35][4] ;
 wire \mem[35][5] ;
 wire \mem[35][6] ;
 wire \mem[35][7] ;
 wire \mem[35][8] ;
 wire \mem[35][9] ;
 wire \mem[36][0] ;
 wire \mem[36][10] ;
 wire \mem[36][11] ;
 wire \mem[36][12] ;
 wire \mem[36][13] ;
 wire \mem[36][14] ;
 wire \mem[36][15] ;
 wire \mem[36][1] ;
 wire \mem[36][2] ;
 wire \mem[36][3] ;
 wire \mem[36][4] ;
 wire \mem[36][5] ;
 wire \mem[36][6] ;
 wire \mem[36][7] ;
 wire \mem[36][8] ;
 wire \mem[36][9] ;
 wire \mem[37][0] ;
 wire \mem[37][10] ;
 wire \mem[37][11] ;
 wire \mem[37][12] ;
 wire \mem[37][13] ;
 wire \mem[37][14] ;
 wire \mem[37][15] ;
 wire \mem[37][1] ;
 wire \mem[37][2] ;
 wire \mem[37][3] ;
 wire \mem[37][4] ;
 wire \mem[37][5] ;
 wire \mem[37][6] ;
 wire \mem[37][7] ;
 wire \mem[37][8] ;
 wire \mem[37][9] ;
 wire \mem[38][0] ;
 wire \mem[38][10] ;
 wire \mem[38][11] ;
 wire \mem[38][12] ;
 wire \mem[38][13] ;
 wire \mem[38][14] ;
 wire \mem[38][15] ;
 wire \mem[38][1] ;
 wire \mem[38][2] ;
 wire \mem[38][3] ;
 wire \mem[38][4] ;
 wire \mem[38][5] ;
 wire \mem[38][6] ;
 wire \mem[38][7] ;
 wire \mem[38][8] ;
 wire \mem[38][9] ;
 wire \mem[39][0] ;
 wire \mem[39][10] ;
 wire \mem[39][11] ;
 wire \mem[39][12] ;
 wire \mem[39][13] ;
 wire \mem[39][14] ;
 wire \mem[39][15] ;
 wire \mem[39][1] ;
 wire \mem[39][2] ;
 wire \mem[39][3] ;
 wire \mem[39][4] ;
 wire \mem[39][5] ;
 wire \mem[39][6] ;
 wire \mem[39][7] ;
 wire \mem[39][8] ;
 wire \mem[39][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[40][0] ;
 wire \mem[40][10] ;
 wire \mem[40][11] ;
 wire \mem[40][12] ;
 wire \mem[40][13] ;
 wire \mem[40][14] ;
 wire \mem[40][15] ;
 wire \mem[40][1] ;
 wire \mem[40][2] ;
 wire \mem[40][3] ;
 wire \mem[40][4] ;
 wire \mem[40][5] ;
 wire \mem[40][6] ;
 wire \mem[40][7] ;
 wire \mem[40][8] ;
 wire \mem[40][9] ;
 wire \mem[41][0] ;
 wire \mem[41][10] ;
 wire \mem[41][11] ;
 wire \mem[41][12] ;
 wire \mem[41][13] ;
 wire \mem[41][14] ;
 wire \mem[41][15] ;
 wire \mem[41][1] ;
 wire \mem[41][2] ;
 wire \mem[41][3] ;
 wire \mem[41][4] ;
 wire \mem[41][5] ;
 wire \mem[41][6] ;
 wire \mem[41][7] ;
 wire \mem[41][8] ;
 wire \mem[41][9] ;
 wire \mem[42][0] ;
 wire \mem[42][10] ;
 wire \mem[42][11] ;
 wire \mem[42][12] ;
 wire \mem[42][13] ;
 wire \mem[42][14] ;
 wire \mem[42][15] ;
 wire \mem[42][1] ;
 wire \mem[42][2] ;
 wire \mem[42][3] ;
 wire \mem[42][4] ;
 wire \mem[42][5] ;
 wire \mem[42][6] ;
 wire \mem[42][7] ;
 wire \mem[42][8] ;
 wire \mem[42][9] ;
 wire \mem[43][0] ;
 wire \mem[43][10] ;
 wire \mem[43][11] ;
 wire \mem[43][12] ;
 wire \mem[43][13] ;
 wire \mem[43][14] ;
 wire \mem[43][15] ;
 wire \mem[43][1] ;
 wire \mem[43][2] ;
 wire \mem[43][3] ;
 wire \mem[43][4] ;
 wire \mem[43][5] ;
 wire \mem[43][6] ;
 wire \mem[43][7] ;
 wire \mem[43][8] ;
 wire \mem[43][9] ;
 wire \mem[44][0] ;
 wire \mem[44][10] ;
 wire \mem[44][11] ;
 wire \mem[44][12] ;
 wire \mem[44][13] ;
 wire \mem[44][14] ;
 wire \mem[44][15] ;
 wire \mem[44][1] ;
 wire \mem[44][2] ;
 wire \mem[44][3] ;
 wire \mem[44][4] ;
 wire \mem[44][5] ;
 wire \mem[44][6] ;
 wire \mem[44][7] ;
 wire \mem[44][8] ;
 wire \mem[44][9] ;
 wire \mem[45][0] ;
 wire \mem[45][10] ;
 wire \mem[45][11] ;
 wire \mem[45][12] ;
 wire \mem[45][13] ;
 wire \mem[45][14] ;
 wire \mem[45][15] ;
 wire \mem[45][1] ;
 wire \mem[45][2] ;
 wire \mem[45][3] ;
 wire \mem[45][4] ;
 wire \mem[45][5] ;
 wire \mem[45][6] ;
 wire \mem[45][7] ;
 wire \mem[45][8] ;
 wire \mem[45][9] ;
 wire \mem[46][0] ;
 wire \mem[46][10] ;
 wire \mem[46][11] ;
 wire \mem[46][12] ;
 wire \mem[46][13] ;
 wire \mem[46][14] ;
 wire \mem[46][15] ;
 wire \mem[46][1] ;
 wire \mem[46][2] ;
 wire \mem[46][3] ;
 wire \mem[46][4] ;
 wire \mem[46][5] ;
 wire \mem[46][6] ;
 wire \mem[46][7] ;
 wire \mem[46][8] ;
 wire \mem[46][9] ;
 wire \mem[47][0] ;
 wire \mem[47][10] ;
 wire \mem[47][11] ;
 wire \mem[47][12] ;
 wire \mem[47][13] ;
 wire \mem[47][14] ;
 wire \mem[47][15] ;
 wire \mem[47][1] ;
 wire \mem[47][2] ;
 wire \mem[47][3] ;
 wire \mem[47][4] ;
 wire \mem[47][5] ;
 wire \mem[47][6] ;
 wire \mem[47][7] ;
 wire \mem[47][8] ;
 wire \mem[47][9] ;
 wire \mem[48][0] ;
 wire \mem[48][10] ;
 wire \mem[48][11] ;
 wire \mem[48][12] ;
 wire \mem[48][13] ;
 wire \mem[48][14] ;
 wire \mem[48][15] ;
 wire \mem[48][1] ;
 wire \mem[48][2] ;
 wire \mem[48][3] ;
 wire \mem[48][4] ;
 wire \mem[48][5] ;
 wire \mem[48][6] ;
 wire \mem[48][7] ;
 wire \mem[48][8] ;
 wire \mem[48][9] ;
 wire \mem[49][0] ;
 wire \mem[49][10] ;
 wire \mem[49][11] ;
 wire \mem[49][12] ;
 wire \mem[49][13] ;
 wire \mem[49][14] ;
 wire \mem[49][15] ;
 wire \mem[49][1] ;
 wire \mem[49][2] ;
 wire \mem[49][3] ;
 wire \mem[49][4] ;
 wire \mem[49][5] ;
 wire \mem[49][6] ;
 wire \mem[49][7] ;
 wire \mem[49][8] ;
 wire \mem[49][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[50][0] ;
 wire \mem[50][10] ;
 wire \mem[50][11] ;
 wire \mem[50][12] ;
 wire \mem[50][13] ;
 wire \mem[50][14] ;
 wire \mem[50][15] ;
 wire \mem[50][1] ;
 wire \mem[50][2] ;
 wire \mem[50][3] ;
 wire \mem[50][4] ;
 wire \mem[50][5] ;
 wire \mem[50][6] ;
 wire \mem[50][7] ;
 wire \mem[50][8] ;
 wire \mem[50][9] ;
 wire \mem[51][0] ;
 wire \mem[51][10] ;
 wire \mem[51][11] ;
 wire \mem[51][12] ;
 wire \mem[51][13] ;
 wire \mem[51][14] ;
 wire \mem[51][15] ;
 wire \mem[51][1] ;
 wire \mem[51][2] ;
 wire \mem[51][3] ;
 wire \mem[51][4] ;
 wire \mem[51][5] ;
 wire \mem[51][6] ;
 wire \mem[51][7] ;
 wire \mem[51][8] ;
 wire \mem[51][9] ;
 wire \mem[52][0] ;
 wire \mem[52][10] ;
 wire \mem[52][11] ;
 wire \mem[52][12] ;
 wire \mem[52][13] ;
 wire \mem[52][14] ;
 wire \mem[52][15] ;
 wire \mem[52][1] ;
 wire \mem[52][2] ;
 wire \mem[52][3] ;
 wire \mem[52][4] ;
 wire \mem[52][5] ;
 wire \mem[52][6] ;
 wire \mem[52][7] ;
 wire \mem[52][8] ;
 wire \mem[52][9] ;
 wire \mem[53][0] ;
 wire \mem[53][10] ;
 wire \mem[53][11] ;
 wire \mem[53][12] ;
 wire \mem[53][13] ;
 wire \mem[53][14] ;
 wire \mem[53][15] ;
 wire \mem[53][1] ;
 wire \mem[53][2] ;
 wire \mem[53][3] ;
 wire \mem[53][4] ;
 wire \mem[53][5] ;
 wire \mem[53][6] ;
 wire \mem[53][7] ;
 wire \mem[53][8] ;
 wire \mem[53][9] ;
 wire \mem[54][0] ;
 wire \mem[54][10] ;
 wire \mem[54][11] ;
 wire \mem[54][12] ;
 wire \mem[54][13] ;
 wire \mem[54][14] ;
 wire \mem[54][15] ;
 wire \mem[54][1] ;
 wire \mem[54][2] ;
 wire \mem[54][3] ;
 wire \mem[54][4] ;
 wire \mem[54][5] ;
 wire \mem[54][6] ;
 wire \mem[54][7] ;
 wire \mem[54][8] ;
 wire \mem[54][9] ;
 wire \mem[55][0] ;
 wire \mem[55][10] ;
 wire \mem[55][11] ;
 wire \mem[55][12] ;
 wire \mem[55][13] ;
 wire \mem[55][14] ;
 wire \mem[55][15] ;
 wire \mem[55][1] ;
 wire \mem[55][2] ;
 wire \mem[55][3] ;
 wire \mem[55][4] ;
 wire \mem[55][5] ;
 wire \mem[55][6] ;
 wire \mem[55][7] ;
 wire \mem[55][8] ;
 wire \mem[55][9] ;
 wire \mem[56][0] ;
 wire \mem[56][10] ;
 wire \mem[56][11] ;
 wire \mem[56][12] ;
 wire \mem[56][13] ;
 wire \mem[56][14] ;
 wire \mem[56][15] ;
 wire \mem[56][1] ;
 wire \mem[56][2] ;
 wire \mem[56][3] ;
 wire \mem[56][4] ;
 wire \mem[56][5] ;
 wire \mem[56][6] ;
 wire \mem[56][7] ;
 wire \mem[56][8] ;
 wire \mem[56][9] ;
 wire \mem[57][0] ;
 wire \mem[57][10] ;
 wire \mem[57][11] ;
 wire \mem[57][12] ;
 wire \mem[57][13] ;
 wire \mem[57][14] ;
 wire \mem[57][15] ;
 wire \mem[57][1] ;
 wire \mem[57][2] ;
 wire \mem[57][3] ;
 wire \mem[57][4] ;
 wire \mem[57][5] ;
 wire \mem[57][6] ;
 wire \mem[57][7] ;
 wire \mem[57][8] ;
 wire \mem[57][9] ;
 wire \mem[58][0] ;
 wire \mem[58][10] ;
 wire \mem[58][11] ;
 wire \mem[58][12] ;
 wire \mem[58][13] ;
 wire \mem[58][14] ;
 wire \mem[58][15] ;
 wire \mem[58][1] ;
 wire \mem[58][2] ;
 wire \mem[58][3] ;
 wire \mem[58][4] ;
 wire \mem[58][5] ;
 wire \mem[58][6] ;
 wire \mem[58][7] ;
 wire \mem[58][8] ;
 wire \mem[58][9] ;
 wire \mem[59][0] ;
 wire \mem[59][10] ;
 wire \mem[59][11] ;
 wire \mem[59][12] ;
 wire \mem[59][13] ;
 wire \mem[59][14] ;
 wire \mem[59][15] ;
 wire \mem[59][1] ;
 wire \mem[59][2] ;
 wire \mem[59][3] ;
 wire \mem[59][4] ;
 wire \mem[59][5] ;
 wire \mem[59][6] ;
 wire \mem[59][7] ;
 wire \mem[59][8] ;
 wire \mem[59][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[60][0] ;
 wire \mem[60][10] ;
 wire \mem[60][11] ;
 wire \mem[60][12] ;
 wire \mem[60][13] ;
 wire \mem[60][14] ;
 wire \mem[60][15] ;
 wire \mem[60][1] ;
 wire \mem[60][2] ;
 wire \mem[60][3] ;
 wire \mem[60][4] ;
 wire \mem[60][5] ;
 wire \mem[60][6] ;
 wire \mem[60][7] ;
 wire \mem[60][8] ;
 wire \mem[60][9] ;
 wire \mem[61][0] ;
 wire \mem[61][10] ;
 wire \mem[61][11] ;
 wire \mem[61][12] ;
 wire \mem[61][13] ;
 wire \mem[61][14] ;
 wire \mem[61][15] ;
 wire \mem[61][1] ;
 wire \mem[61][2] ;
 wire \mem[61][3] ;
 wire \mem[61][4] ;
 wire \mem[61][5] ;
 wire \mem[61][6] ;
 wire \mem[61][7] ;
 wire \mem[61][8] ;
 wire \mem[61][9] ;
 wire \mem[62][0] ;
 wire \mem[62][10] ;
 wire \mem[62][11] ;
 wire \mem[62][12] ;
 wire \mem[62][13] ;
 wire \mem[62][14] ;
 wire \mem[62][15] ;
 wire \mem[62][1] ;
 wire \mem[62][2] ;
 wire \mem[62][3] ;
 wire \mem[62][4] ;
 wire \mem[62][5] ;
 wire \mem[62][6] ;
 wire \mem[62][7] ;
 wire \mem[62][8] ;
 wire \mem[62][9] ;
 wire \mem[63][0] ;
 wire \mem[63][10] ;
 wire \mem[63][11] ;
 wire \mem[63][12] ;
 wire \mem[63][13] ;
 wire \mem[63][14] ;
 wire \mem[63][15] ;
 wire \mem[63][1] ;
 wire \mem[63][2] ;
 wire \mem[63][3] ;
 wire \mem[63][4] ;
 wire \mem[63][5] ;
 wire \mem[63][6] ;
 wire \mem[63][7] ;
 wire \mem[63][8] ;
 wire \mem[63][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_00007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(_00009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_888 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1066 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_899 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1086 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_744 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_878 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1005 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1024 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1041 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_423 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_420 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_965 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_987 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1004 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1016 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_806 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_880 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_421 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_71 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_910 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1066 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_641 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1093 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_446 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_880 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_526 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_956 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1076 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_464 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_528 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_665 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_621 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_91 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1035 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_587 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_601 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_423 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_71 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_841 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_918 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_90 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1015 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1062 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1035 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1058 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_771 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1099 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_54 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_64 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_78 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_790 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_895 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_530 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_895 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_975 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_565 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1001 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1076 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_30 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_413 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_549 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_802 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_14 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_388 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_618 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_78 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_880 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_91 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_351 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_544 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_587 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_630 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_94 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_455 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_46 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_62 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_78 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_423 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_701 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1020 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_575 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_657 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_967 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1036 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_673 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_717 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_925 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_501 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_71 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_835 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_994 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_20 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_608 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_932 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1006 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1050 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_411 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_774 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_86 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_897 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_899 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_972 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_48 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_525 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_56 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_668 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_878 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_959 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_573 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1059 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_39 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_51 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_806 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_92 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_940 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_996 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_532 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_571 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_587 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_79 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_910 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1096 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_385 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_6 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_67 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_671 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_821 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_950 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_26 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_423 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_510 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_533 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_712 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1016 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1020 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1086 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_412 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_42 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_525 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_566 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_598 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_600 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_68 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_763 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_895 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_897 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1010 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1331 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_229 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_465 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_490 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1070 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1355 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_43 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_432 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_47 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_485 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_57 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_721 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_81 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_854 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_897 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_899 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1031 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_74 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_925 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1037 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_12 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_21 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_29 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_33 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_43 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_52 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_700 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_866 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_895 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_10 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1072 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_22 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_327 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_430 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_434 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_44 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_60 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_736 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_957 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1210 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_428 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_463 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_564 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_851 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_995 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1018 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1020 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1034 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1042 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1077 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_216 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_336 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_338 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_590 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_689 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_792 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_794 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_824 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_481 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_55 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_552 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_59 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_611 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_993 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1028 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1044 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1371 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_623 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_643 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_659 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_715 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_723 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_736 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_796 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_953 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1051 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1060 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1075 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1083 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_509 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_536 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_617 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_728 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_779 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_841 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_870 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_892 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_923 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_999 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1088 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1228 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1264 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_389 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_439 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_49 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_645 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_752 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_788 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_990 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1018 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1020 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1091 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_149 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_287 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_301 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_609 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_766 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_805 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_837 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_962 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1054 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1072 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_323 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_350 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_513 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_541 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_638 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_660 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_678 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_82 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_826 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_90 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_980 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1026 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1030 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1097 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_162 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_479 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_487 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_577 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_743 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_79 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_798 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_814 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_83 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_919 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_969 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_309 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_345 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_45 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_466 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_497 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_567 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_637 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_653 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_755 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_83 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_901 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_905 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_911 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1035 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1098 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_261 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_373 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_38 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_40 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_408 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_534 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_582 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_622 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_668 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_676 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_692 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_758 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_863 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_895 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1053 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1183 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1322 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_357 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_370 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_41 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_450 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_560 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_647 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_753 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_773 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_856 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_913 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_97 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_989 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_991 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1072 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1079 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1103 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_588 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_596 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_636 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_642 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_697 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_776 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_778 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_809 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_813 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_829 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_833 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_844 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_931 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_945 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_965 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1061 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1069 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1080 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1218 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1364 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_254 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_353 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_391 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_405 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_423 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_425 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_563 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_613 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_713 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_731 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_983 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1295 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_241 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_414 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_456 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_460 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_468 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_484 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_50 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_58 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_735 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_787 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_817 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_881 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_891 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_902 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_943 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1007 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1152 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1159 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1253 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1280 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_148 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_324 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_361 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_383 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_409 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_469 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_477 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_521 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_585 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_655 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_683 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_685 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_812 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_860 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_897 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_929 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1035 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1180 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1211 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_359 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_378 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_480 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_554 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_606 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_649 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_651 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_686 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_722 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_785 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_808 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_810 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_828 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_850 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_907 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_935 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_939 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_963 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1072 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1078 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1181 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_121 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_341 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_365 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_462 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_515 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_529 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_569 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_583 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_767 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_77 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_797 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_845 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_853 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_89 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_922 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_983 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_985 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1068 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1076 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_126 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1293 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_169 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_263 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_339 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_355 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_363 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_440 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_461 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_537 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_553 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_557 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_589 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_593 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_604 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_639 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_652 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_775 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_800 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_804 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_827 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_834 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_857 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_868 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_872 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_903 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_926 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_928 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_937 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_958 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1040 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1072 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1130 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1134 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1334 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_249 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_265 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_319 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_426 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_436 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_445 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_447 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_489 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_507 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_540 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_581 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_625 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_693 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_739 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_76 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_760 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_819 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_906 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1023 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1029 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1063 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1071 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1240 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1276 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1284 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_307 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_333 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_418 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_448 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_452 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_454 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_475 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_490 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_508 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_53 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_531 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_542 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_548 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_578 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_607 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_61 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_65 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_650 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_658 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_684 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_690 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_704 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_729 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_845 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_893 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_897 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_921 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_934 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_96 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_986 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_997 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1225 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_292 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_312 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_374 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_382 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_386 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_388 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_402 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_499 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_503 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_505 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_646 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_662 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_670 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_734 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_742 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_746 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_748 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_757 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_765 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_772 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_780 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_839 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_849 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_865 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_876 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_884 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_974 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_978 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_992 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1000 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1008 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1012 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_102 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1073 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1123 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1127 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1151 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1157 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1161 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1163 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1186 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1221 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_125 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_230 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_252 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_354 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_384 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_420 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_451 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_504 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_517 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_535 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_631 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_661 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_679 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_706 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_727 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_85 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_87 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_877 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_889 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_896 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_933 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_970 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_98 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1014 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1057 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1113 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1117 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1203 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1232 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1268 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1332 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_272 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_300 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_335 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_344 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_375 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_415 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_424 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_438 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_442 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_516 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_556 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_579 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_602 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_615 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_698 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_732 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_88 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_927 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_95 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_984 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_99 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1003 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1074 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1094 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1213 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1273 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1289 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1306 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1346 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1398 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_165 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_167 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_256 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_285 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_355 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_381 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_403 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_429 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_433 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_457 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_514 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_633 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_635 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_708 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_71 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_726 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_733 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_737 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_754 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_770 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_782 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_786 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_822 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_830 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_840 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_874 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_885 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_887 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_955 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_971 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1002 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1018 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1038 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1046 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1081 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1281 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1315 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1394 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_193 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_200 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_204 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_288 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_296 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_390 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_476 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_591 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_595 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_610 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_616 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_624 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_628 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_664 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_680 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_688 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_694 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_749 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_769 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_816 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_842 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_909 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_917 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_924 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_965 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1009 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1025 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1033 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1039 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1041 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1055 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1064 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1072 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1076 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1116 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1153 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1219 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1369 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_291 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_302 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_392 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_431 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_470 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_518 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_522 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_572 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_584 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_592 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_605 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_612 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_654 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_656 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_677 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_695 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_703 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_705 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_793 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_820 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_858 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_862 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_864 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_952 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_960 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_964 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_966 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1011 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1013 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1089 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_110 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1115 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1146 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1154 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1237 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1259 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1267 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1310 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1316 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1337 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_173 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_217 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_233 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_311 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_343 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_380 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_396 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_400 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_417 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_419 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_422 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_453 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_506 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_538 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_550 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_570 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_574 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_626 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_640 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_764 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_768 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_801 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_838 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_871 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_875 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_912 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_914 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_973 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1032 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1052 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1084 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1132 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_114 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1170 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_118 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1185 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1189 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1222 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1236 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1248 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_129 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1304 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_133 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1340 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1397 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1399 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_168 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_184 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_188 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_226 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_234 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_238 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_277 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_348 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_356 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_377 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_393 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_407 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_427 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_435 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_437 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_443 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_459 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_467 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_474 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_500 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_502 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_511 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_519 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_558 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_620 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_634 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_687 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_696 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_707 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_709 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_719 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_762 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_781 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_783 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_789 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_795 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_811 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_825 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_847 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_855 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_859 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_861 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_867 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_875 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_883 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_968 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_976 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1022 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1056 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1090 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1158 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1192 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_120 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1255 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1257 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1260 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_131 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1328 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1367 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_206 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_269 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_271 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_274 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_290 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_308 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_342 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_358 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_36 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_366 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_376 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_410 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_444 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_478 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_486 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_488 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_494 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_546 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_614 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_648 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_682 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_716 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_725 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_741 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_745 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_750 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_784 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_818 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_852 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_886 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_894 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_908 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_916 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_920 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_936 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_947 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_951 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_954 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_988 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1017 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1021 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1048 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1087 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_109 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1147 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1175 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1194 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1224 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1227 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_124 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1245 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1275 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1297 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_135 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1401 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_143 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_145 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_190 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_199 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_251 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_266 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_313 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_387 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_395 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_404 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_406 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_441 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_449 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_491 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_493 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_523 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_527 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_547 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_555 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_568 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_576 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_580 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_586 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_597 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_599 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_672 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_674 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_681 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_718 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_720 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_75 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_756 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_791 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_799 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_803 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_807 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_823 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_832 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_848 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_869 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_873 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_882 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_898 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_900 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_930 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_938 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_942 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_944 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_981 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_985 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_100 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1019 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1027 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1043 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1047 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1049 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_106 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1065 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1067 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1082 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1095 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1111 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1119 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_112 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1122 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1138 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1140 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1178 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1182 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1239 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1258 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1262 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_128 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1299 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_156 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_198 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_207 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_223 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_235 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_270 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_278 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_303 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_320 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_347 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_349 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_352 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_360 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_362 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_368 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_372 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_379 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_458 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_471 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_473 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_482 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_492 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_496 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_498 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_512 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_520 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_524 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_539 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_543 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_545 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_551 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_559 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_562 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_594 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_603 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_619 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_627 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_629 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_632 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_644 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_663 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_667 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_669 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_675 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_691 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_699 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_702 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_710 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_714 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_724 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_730 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_738 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_740 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_747 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_751 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_759 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_761 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_777 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_80 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_815 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_831 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_84 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_879 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_890 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_93 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_941 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_949 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_961 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_977 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_979 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_982 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_998 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_81 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_91 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_92 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_93 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_94 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_95 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_96 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_97 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_98 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_99 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_100 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_82 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_102 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_103 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_104 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_106 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_107 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_109 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_110 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_83 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_111 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_112 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_113 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_114 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_115 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_116 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_117 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_118 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_119 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_120 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_84 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_121 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_122 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_123 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_124 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_125 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_126 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_127 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_128 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_129 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_130 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_85 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_133 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_134 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_135 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_136 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_138 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_140 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_86 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_143 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_145 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_146 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_147 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_148 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_149 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_150 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_87 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_151 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_152 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_153 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_154 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_155 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_156 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_157 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_158 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_159 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_160 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_88 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_161 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_89 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_90 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_162 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_163 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_164 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_165 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_166 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_167 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_168 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_169 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_170 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_171 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_173 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_174 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_175 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_177 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_178 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_180 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_181 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_182 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_183 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_184 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_185 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_186 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_187 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_188 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_189 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_190 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_191 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_193 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_194 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_195 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_196 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_197 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_198 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_199 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_200 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_201 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_202 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_383 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_384 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_386 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_387 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_388 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_390 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_391 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_393 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_394 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_395 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_396 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_397 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_398 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_399 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_400 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_401 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_402 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_403 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_404 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_406 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_407 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_409 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_410 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_411 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_415 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_418 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_420 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_421 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_422 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_423 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_424 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_425 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_426 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_427 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_428 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_429 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_430 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_431 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_432 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_433 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_434 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_435 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_436 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_437 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_438 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_439 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_440 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_441 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_442 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_443 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_444 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_445 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_446 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_447 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_448 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_449 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_450 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_451 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_452 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_453 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_454 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_455 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_456 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_457 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_458 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_459 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_460 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_461 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_462 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_463 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_464 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_465 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_466 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_467 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_468 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_469 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_470 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_471 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_472 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_473 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_474 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_475 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_476 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_477 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_478 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_479 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_480 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_481 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_482 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_483 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_484 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_485 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_486 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_487 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_488 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_489 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_490 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_491 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_492 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_493 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_494 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_495 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_496 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_497 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_498 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_499 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_500 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_501 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_502 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_503 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_504 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_505 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_506 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_507 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_508 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_509 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_510 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_511 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_512 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_513 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_514 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_515 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_516 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_517 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_518 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_519 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_520 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_521 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_522 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_523 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_524 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_525 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_526 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_527 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_528 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_529 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_530 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_531 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_532 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_533 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_534 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_535 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_536 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_537 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_538 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_539 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_540 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_541 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_542 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_543 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_544 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_545 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_546 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_547 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_548 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_549 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_550 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_551 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_552 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_553 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_554 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_555 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_556 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_557 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_558 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_559 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_560 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_561 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_562 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_563 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_564 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_565 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_566 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_567 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_568 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_569 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_570 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_571 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_572 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_573 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_574 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_575 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_576 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_577 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_578 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_579 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_580 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_581 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_582 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_203 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_204 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_205 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_206 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_207 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_210 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_211 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_213 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_214 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_216 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_217 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_218 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_219 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_220 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_221 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_222 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_583 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_584 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_585 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_586 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_587 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_588 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_589 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_590 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_591 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_592 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_593 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_594 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_595 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_596 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_597 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_598 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_599 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_600 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_601 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_602 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_603 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_604 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_605 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_606 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_607 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_608 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_609 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_610 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_611 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_612 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_613 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_614 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_615 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_616 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_617 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_618 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_619 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_620 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_621 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_622 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_623 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_624 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_625 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_626 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_627 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_628 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_629 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_630 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_631 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_632 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_633 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_634 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_635 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_636 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_637 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_638 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_639 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_640 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_641 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_642 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_643 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_644 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_645 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_646 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_647 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_648 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_649 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_650 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_651 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_652 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_653 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_654 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_655 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_656 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_657 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_658 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_659 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_660 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_661 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_662 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_663 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_664 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_665 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_666 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_667 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_668 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_669 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_670 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_671 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_672 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_673 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_674 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_675 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_676 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_677 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_678 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_679 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_680 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_681 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_682 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_683 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_684 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_685 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_686 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_687 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_688 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_689 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_690 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_691 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_692 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_693 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_694 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_695 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_696 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_697 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_698 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_699 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_700 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_701 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_702 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_703 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_704 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_705 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_706 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_707 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_708 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_709 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_710 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_711 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_712 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_713 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_714 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_715 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_716 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_717 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_718 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_719 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_720 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_721 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_722 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_723 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_724 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_725 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_726 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_727 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_728 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_729 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_730 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_731 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_732 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_733 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_734 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_735 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_736 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_737 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_738 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_739 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_740 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_741 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_742 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_743 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_744 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_745 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_746 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_747 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_748 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_749 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_750 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_751 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_752 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_753 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_754 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_755 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_756 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_757 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_758 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_759 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_760 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_761 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_762 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_763 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_764 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_765 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_766 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_767 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_768 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_769 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_770 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_771 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_772 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_773 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_774 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_775 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_776 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_777 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_778 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_779 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_780 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_781 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_782 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_223 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_224 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_225 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_226 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_227 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_228 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_229 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_230 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_231 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_232 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_233 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_234 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_235 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_236 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_237 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_238 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_239 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_240 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_241 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_242 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_783 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_784 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_785 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_786 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_787 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_788 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_789 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_790 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_791 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_792 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_793 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_794 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_795 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_796 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_797 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_798 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_799 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_800 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_801 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_802 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_803 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_804 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_805 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_806 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_807 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_808 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_809 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_810 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_811 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_812 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_813 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_814 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_815 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_816 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_817 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_818 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_819 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_820 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_821 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_822 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_823 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_824 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_825 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_826 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_827 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_828 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_829 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_830 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_831 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_832 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_833 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_834 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_835 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_836 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_837 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_838 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_839 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_840 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_841 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_842 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_843 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_844 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_845 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_846 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_847 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_848 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_849 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_850 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_851 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_852 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_853 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_854 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_855 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_856 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_857 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_858 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_859 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_860 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_861 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_862 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_863 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_864 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_865 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_866 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_867 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_868 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_869 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_870 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_871 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_872 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_873 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_874 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_875 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_876 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_877 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_878 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_879 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_880 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_881 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_882 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_883 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_884 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_885 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_886 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_887 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_888 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_889 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_890 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_891 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_892 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_893 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_894 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_895 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_896 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_897 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_898 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_899 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_900 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_901 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_902 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_903 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_904 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_905 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_906 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_907 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_908 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_909 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_910 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_911 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_912 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_913 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_914 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_915 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_916 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_917 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_918 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_919 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_920 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_921 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_922 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_923 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_924 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_925 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_926 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_927 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_928 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_929 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_930 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_931 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_932 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_933 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_934 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_935 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_936 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_937 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_938 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_939 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_940 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_941 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_942 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_943 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_944 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_945 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_946 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_947 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_948 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_949 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_950 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_951 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_952 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_953 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_954 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_955 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_956 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_957 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_958 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_959 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_960 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_961 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_962 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_963 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_964 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_965 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_966 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_967 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_968 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_969 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_970 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_971 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_972 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_973 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_974 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_975 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_976 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_977 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_978 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_979 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_980 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_981 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_982 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_244 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_245 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_246 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_248 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_249 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_251 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_252 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_253 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_254 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_255 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_256 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_257 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_258 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_259 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_260 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_261 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_262 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1000 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1001 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1002 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_983 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_984 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_985 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_986 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_987 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_988 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_989 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_990 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_991 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_992 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_993 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_994 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_995 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_996 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_997 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_998 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_999 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1003 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1004 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1005 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1006 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1007 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1008 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1009 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1010 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1011 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1012 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1013 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1014 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1015 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1016 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1017 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1018 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1019 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1020 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1021 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1022 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1023 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1024 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1025 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1026 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1027 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1028 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1029 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1030 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1031 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1032 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1033 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1034 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1035 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1036 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1037 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1038 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1039 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1040 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1041 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1042 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1043 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1044 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1045 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1046 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1047 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1048 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1049 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1050 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1051 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1052 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1053 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1054 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1055 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1056 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1057 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1058 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1059 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1060 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1061 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1062 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1063 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1064 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1065 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1066 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1067 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1068 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1069 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1070 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1071 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1072 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1073 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1074 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1075 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1076 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1077 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1078 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1079 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1080 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1081 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1082 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1083 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1084 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1085 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1086 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1087 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1088 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1089 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1090 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1091 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1092 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1093 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1094 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1095 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1096 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1097 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1098 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1099 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1100 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1102 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1103 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1104 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1106 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1107 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1109 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1110 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1111 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1112 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1113 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1114 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1115 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1116 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1117 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1118 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1119 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1120 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1121 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1122 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1123 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1124 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1125 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1126 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1127 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1128 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1129 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1130 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1133 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1134 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1135 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1136 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1138 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1140 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1143 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1145 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1146 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1147 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1148 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1149 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1150 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1151 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1152 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1153 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1154 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1155 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1156 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1157 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1158 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1159 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1160 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1161 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1162 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1163 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1164 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1165 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1166 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1167 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1168 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1169 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1170 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1171 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1173 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1174 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1175 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1177 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1178 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1180 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1181 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1182 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_263 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_264 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_265 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_266 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_267 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_268 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_269 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_270 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_271 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_272 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_273 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_274 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_275 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_276 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_277 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_278 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_280 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_281 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_282 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1183 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1184 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1185 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1186 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1187 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1188 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1189 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1190 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1191 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1193 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1194 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1195 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1196 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1197 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1198 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1199 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1200 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1201 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1202 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1203 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1204 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1205 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1206 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1207 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1210 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1211 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1213 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1214 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1216 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1217 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1218 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1219 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1220 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1221 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1222 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1223 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1224 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1225 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1226 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1227 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1228 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1229 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1230 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1231 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1232 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1233 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1234 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1235 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1236 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1237 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1238 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1239 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1240 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1241 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1242 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1244 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1245 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1246 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1248 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1249 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1251 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1252 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1253 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1254 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1255 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1256 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1257 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1258 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1259 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1260 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1261 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1262 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1263 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1264 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1265 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1266 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1267 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1268 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1269 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1270 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1271 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1272 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1273 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1274 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1275 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1276 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1277 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1278 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1280 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1281 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1282 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1284 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1285 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1287 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1288 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1289 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1290 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1291 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1292 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1293 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1294 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1295 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1296 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1297 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1298 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1299 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1300 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1301 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1302 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1303 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1304 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1305 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1306 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1307 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1308 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1309 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1310 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1311 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1312 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1313 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1315 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1316 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1317 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1319 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1320 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1322 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1323 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1324 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1325 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1326 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1327 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1328 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1329 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1330 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1331 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1332 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1333 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1334 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1335 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1336 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1337 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1338 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1339 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1340 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1341 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1342 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1343 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1344 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1345 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1346 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1347 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1348 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1349 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1351 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1353 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1355 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1356 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1358 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1359 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1360 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1361 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1362 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1363 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1364 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1365 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1366 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1367 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1368 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1369 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1370 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1371 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1372 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1373 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1374 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1375 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1376 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1377 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1378 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1379 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1380 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1381 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1382 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_284 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_285 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_287 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_288 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_289 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_290 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_291 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_292 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_293 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_294 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_295 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_296 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_297 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_298 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_299 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_300 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_301 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_302 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1383 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1384 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1386 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1387 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1388 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1390 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1391 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1393 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1394 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1395 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1396 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1397 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1398 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1399 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1400 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1401 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1402 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1403 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1404 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1406 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1407 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1409 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1410 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1411 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1415 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1418 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1420 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1421 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1422 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1423 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1424 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1425 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1426 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1427 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1428 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1429 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1430 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1431 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1432 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1433 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1434 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1435 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1436 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1437 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1438 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1439 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1440 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1441 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1442 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1443 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1444 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1445 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1446 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1447 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1448 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1449 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1450 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1451 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1452 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1453 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1454 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1455 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1456 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1457 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1458 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1459 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1460 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1461 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1462 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1463 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1464 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1465 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1466 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1467 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1468 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1469 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1470 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1471 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1472 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1473 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1474 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1475 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1476 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1477 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1478 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1479 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1480 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1481 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1482 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1483 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1484 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1485 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1486 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1487 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1488 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1489 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1490 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1491 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1492 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1493 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1494 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1495 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1496 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1497 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1498 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1499 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1500 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1501 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1502 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1503 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1504 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1505 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1506 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1507 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1508 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1509 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1510 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1511 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1512 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1513 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1514 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1515 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1516 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1517 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1518 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1519 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1520 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1521 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1522 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1523 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1524 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1525 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1526 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1527 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1528 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1529 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1530 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1531 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1532 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1533 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1534 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1535 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1536 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1537 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1538 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1539 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1540 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1541 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1542 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1543 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1544 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1545 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1546 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1547 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1548 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1549 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1550 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1551 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1552 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1553 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1554 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1555 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1556 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1557 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1558 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1559 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1560 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1561 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1562 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1563 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1564 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1565 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1566 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1567 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1568 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1569 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1570 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1571 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1572 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1573 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1574 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1575 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1576 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1577 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1578 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1579 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1580 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1581 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1582 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_303 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_304 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_305 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_306 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_307 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_308 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_309 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_310 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_311 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_312 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_313 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_315 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_316 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_317 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_319 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_320 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_322 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1583 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1584 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1585 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1586 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1587 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1588 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1589 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1590 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1591 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1592 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1593 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1594 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1595 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1596 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1597 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1598 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1599 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1600 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1601 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1602 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1603 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1604 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1605 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1606 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1607 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1608 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1609 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1610 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1611 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1612 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1613 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1614 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1615 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1616 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1617 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1618 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1619 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1620 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1621 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1622 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1623 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1624 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1625 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1626 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1627 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1628 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1629 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1630 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1631 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1632 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1633 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1634 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1635 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1636 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1637 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1638 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1639 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1640 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1641 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1642 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1643 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1644 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1645 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1646 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1647 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1648 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1649 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1650 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1651 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1652 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1653 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1654 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1655 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1656 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1657 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1658 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1659 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1660 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1661 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1662 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1663 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1664 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1665 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1666 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1667 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1668 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1669 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1670 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1671 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1672 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1673 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1674 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1675 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1676 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1677 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1678 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1679 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1680 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1681 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1682 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1683 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1684 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1685 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1686 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1687 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1688 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1689 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1690 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1691 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1692 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1693 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1694 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1695 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1696 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1697 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1698 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1699 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1700 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1701 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1702 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1703 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1704 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1705 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1706 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1707 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1708 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1709 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1710 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1711 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1712 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1713 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1714 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1715 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1716 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1717 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1718 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1719 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1720 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1721 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1722 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1723 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1724 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1725 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1726 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1727 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1728 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1729 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1730 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1731 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1732 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1733 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1734 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1735 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1736 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1737 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1738 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1739 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1740 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1741 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1742 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1743 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1744 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1745 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1746 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1747 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1748 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1749 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1750 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1751 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1752 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1753 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1754 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1755 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1756 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1757 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1758 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1759 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1760 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1761 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1762 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1763 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1764 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1765 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1766 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1767 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1768 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1769 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1770 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1771 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1772 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1773 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1774 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1775 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1776 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1777 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1778 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1779 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1780 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1781 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1782 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_323 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_324 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_325 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_326 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_327 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_328 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_329 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_330 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_331 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_332 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_333 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_334 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_335 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_336 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_337 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_338 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_339 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_340 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_341 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_342 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1783 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1784 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1785 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1786 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1787 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1788 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1789 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1790 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1791 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1792 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1793 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1794 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1795 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1796 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1797 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1798 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1799 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1800 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1801 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1802 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1803 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1804 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1805 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1806 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1807 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1808 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1809 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1810 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1811 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1812 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1813 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1814 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1815 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1816 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1817 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1818 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1819 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1820 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1821 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1822 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1823 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_343 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_344 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_345 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_346 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_347 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_348 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_349 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_351 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_353 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_355 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_356 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_358 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_359 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_360 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_361 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_362 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_363 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_364 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_365 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_366 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_367 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_368 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_369 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_370 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_371 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_372 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_373 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_374 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_375 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_376 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_377 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_378 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_379 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_380 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_381 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_382 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04854_ (.A1(_04153_),
    .A2(_04133_),
    .B(_04154_),
    .ZN(_00508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _04855_ (.I(_03489_),
    .Z(_04155_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04856_ (.A1(_04143_),
    .A2(\mem[33][10] ),
    .ZN(_04156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04857_ (.A1(_04155_),
    .A2(_04134_),
    .B(_04156_),
    .ZN(_00509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _04858_ (.I(_03492_),
    .Z(_04157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04859_ (.A1(_04143_),
    .A2(\mem[33][11] ),
    .ZN(_04158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04860_ (.A1(_04157_),
    .A2(_04134_),
    .B(_04158_),
    .ZN(_00510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _04861_ (.I(_03495_),
    .Z(_04159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04862_ (.A1(_04143_),
    .A2(\mem[33][12] ),
    .ZN(_04160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04863_ (.A1(_04159_),
    .A2(_04134_),
    .B(_04160_),
    .ZN(_00511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04864_ (.A1(_04143_),
    .A2(\mem[33][13] ),
    .ZN(_04161_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04865_ (.A1(_04125_),
    .A2(_04134_),
    .B(_04161_),
    .ZN(_00512_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04866_ (.A1(_04132_),
    .A2(\mem[33][14] ),
    .ZN(_04162_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04867_ (.A1(_04127_),
    .A2(_04134_),
    .B(_04162_),
    .ZN(_00513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04868_ (.A1(_04132_),
    .A2(\mem[33][15] ),
    .ZN(_04163_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04869_ (.A1(_04129_),
    .A2(_04134_),
    .B(_04163_),
    .ZN(_00514_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _04870_ (.A1(_03631_),
    .A2(_03440_),
    .ZN(_04164_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _04871_ (.A1(_04164_),
    .A2(_01127_),
    .ZN(_04165_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04872_ (.I(_04165_),
    .Z(_04166_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04873_ (.I(_04165_),
    .Z(_04167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04874_ (.A1(_04167_),
    .A2(\mem[34][0] ),
    .ZN(_04168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04875_ (.A1(_04131_),
    .A2(_04166_),
    .B(_04168_),
    .ZN(_00515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04876_ (.A1(_04167_),
    .A2(\mem[34][1] ),
    .ZN(_04169_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04877_ (.A1(_04136_),
    .A2(_04166_),
    .B(_04169_),
    .ZN(_00516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04878_ (.A1(_04167_),
    .A2(\mem[34][2] ),
    .ZN(_04170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04879_ (.A1(_04138_),
    .A2(_04166_),
    .B(_04170_),
    .ZN(_00517_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04880_ (.A1(_04167_),
    .A2(\mem[34][3] ),
    .ZN(_04171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04881_ (.A1(_04140_),
    .A2(_04166_),
    .B(_04171_),
    .ZN(_00518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04882_ (.I(_04165_),
    .Z(_04172_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04883_ (.A1(_04172_),
    .A2(\mem[34][4] ),
    .ZN(_04173_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04884_ (.A1(_04142_),
    .A2(_04166_),
    .B(_04173_),
    .ZN(_00519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04885_ (.A1(_04172_),
    .A2(\mem[34][5] ),
    .ZN(_04174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04886_ (.A1(_04145_),
    .A2(_04166_),
    .B(_04174_),
    .ZN(_00520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04887_ (.A1(_04172_),
    .A2(\mem[34][6] ),
    .ZN(_04175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04888_ (.A1(_04147_),
    .A2(_04166_),
    .B(_04175_),
    .ZN(_00521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04889_ (.A1(_04172_),
    .A2(\mem[34][7] ),
    .ZN(_04176_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04890_ (.A1(_04149_),
    .A2(_04166_),
    .B(_04176_),
    .ZN(_00522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04891_ (.A1(_04172_),
    .A2(\mem[34][8] ),
    .ZN(_04177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04892_ (.A1(_04151_),
    .A2(_04166_),
    .B(_04177_),
    .ZN(_00523_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04893_ (.A1(_04172_),
    .A2(\mem[34][9] ),
    .ZN(_04178_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04894_ (.A1(_04153_),
    .A2(_04166_),
    .B(_04178_),
    .ZN(_00524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04895_ (.A1(_04172_),
    .A2(\mem[34][10] ),
    .ZN(_04179_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04896_ (.A1(_04155_),
    .A2(_04167_),
    .B(_04179_),
    .ZN(_00525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04897_ (.A1(_04172_),
    .A2(\mem[34][11] ),
    .ZN(_04180_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04898_ (.A1(_04157_),
    .A2(_04167_),
    .B(_04180_),
    .ZN(_00526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04899_ (.A1(_04172_),
    .A2(\mem[34][12] ),
    .ZN(_04181_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04900_ (.A1(_04159_),
    .A2(_04167_),
    .B(_04181_),
    .ZN(_00527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04901_ (.A1(_04172_),
    .A2(\mem[34][13] ),
    .ZN(_04182_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04902_ (.A1(_04125_),
    .A2(_04167_),
    .B(_04182_),
    .ZN(_00528_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04903_ (.A1(_04165_),
    .A2(\mem[34][14] ),
    .ZN(_04183_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04904_ (.A1(_04127_),
    .A2(_04167_),
    .B(_04183_),
    .ZN(_00529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04905_ (.A1(_04165_),
    .A2(\mem[34][15] ),
    .ZN(_04184_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04906_ (.A1(_04129_),
    .A2(_04167_),
    .B(_04184_),
    .ZN(_00530_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _04907_ (.A1(_03543_),
    .A2(net76),
    .ZN(_04185_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04908_ (.I(_04185_),
    .Z(_04186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04909_ (.I(_04185_),
    .Z(_04187_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04910_ (.A1(_04187_),
    .A2(\mem[35][0] ),
    .ZN(_04188_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04911_ (.A1(_04131_),
    .A2(_04186_),
    .B(_04188_),
    .ZN(_00531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04912_ (.A1(_04187_),
    .A2(\mem[35][1] ),
    .ZN(_04189_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04913_ (.A1(_04136_),
    .A2(_04186_),
    .B(_04189_),
    .ZN(_00532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04914_ (.A1(_04187_),
    .A2(\mem[35][2] ),
    .ZN(_04190_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04915_ (.A1(_04138_),
    .A2(_04186_),
    .B(_04190_),
    .ZN(_00533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04916_ (.A1(_04187_),
    .A2(\mem[35][3] ),
    .ZN(_04191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04917_ (.A1(_04140_),
    .A2(_04186_),
    .B(_04191_),
    .ZN(_00534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04918_ (.I(_04185_),
    .Z(_04192_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04919_ (.A1(_04192_),
    .A2(\mem[35][4] ),
    .ZN(_04193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04920_ (.A1(_04142_),
    .A2(_04186_),
    .B(_04193_),
    .ZN(_00535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04921_ (.A1(_04192_),
    .A2(\mem[35][5] ),
    .ZN(_04194_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04922_ (.A1(_04145_),
    .A2(_04186_),
    .B(_04194_),
    .ZN(_00536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04923_ (.A1(_04192_),
    .A2(\mem[35][6] ),
    .ZN(_04195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04924_ (.A1(_04147_),
    .A2(_04186_),
    .B(_04195_),
    .ZN(_00537_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04925_ (.A1(_04192_),
    .A2(\mem[35][7] ),
    .ZN(_04196_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04926_ (.A1(_04149_),
    .A2(_04186_),
    .B(_04196_),
    .ZN(_00538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04927_ (.A1(_04192_),
    .A2(\mem[35][8] ),
    .ZN(_04197_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04928_ (.A1(_04151_),
    .A2(_04186_),
    .B(_04197_),
    .ZN(_00539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04929_ (.A1(_04192_),
    .A2(\mem[35][9] ),
    .ZN(_04198_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04930_ (.A1(_04153_),
    .A2(_04186_),
    .B(_04198_),
    .ZN(_00540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04931_ (.A1(_04192_),
    .A2(\mem[35][10] ),
    .ZN(_04199_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04932_ (.A1(_04155_),
    .A2(_04187_),
    .B(_04199_),
    .ZN(_00541_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04933_ (.A1(_04192_),
    .A2(\mem[35][11] ),
    .ZN(_04200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04934_ (.A1(_04157_),
    .A2(_04187_),
    .B(_04200_),
    .ZN(_00542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04935_ (.A1(_04192_),
    .A2(\mem[35][12] ),
    .ZN(_04201_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04936_ (.A1(_04159_),
    .A2(_04187_),
    .B(_04201_),
    .ZN(_00543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04937_ (.A1(_04192_),
    .A2(\mem[35][13] ),
    .ZN(_04202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04938_ (.A1(_04125_),
    .A2(_04187_),
    .B(_04202_),
    .ZN(_00544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04939_ (.A1(_04185_),
    .A2(\mem[35][14] ),
    .ZN(_04203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04940_ (.A1(_04127_),
    .A2(_04187_),
    .B(_04203_),
    .ZN(_00545_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04941_ (.A1(_04185_),
    .A2(\mem[35][15] ),
    .ZN(_04204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04942_ (.A1(_04129_),
    .A2(_04187_),
    .B(_04204_),
    .ZN(_00546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _04943_ (.A1(net132),
    .A2(net91),
    .Z(_04205_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _04944_ (.A1(_04205_),
    .A2(net76),
    .ZN(_04206_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04945_ (.I(_04206_),
    .Z(_04207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04946_ (.I(_04206_),
    .Z(_04208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04947_ (.A1(_04208_),
    .A2(\mem[36][0] ),
    .ZN(_04209_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04948_ (.A1(_04131_),
    .A2(_04207_),
    .B(_04209_),
    .ZN(_00547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04949_ (.A1(_04208_),
    .A2(\mem[36][1] ),
    .ZN(_04210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04950_ (.A1(_04136_),
    .A2(_04207_),
    .B(_04210_),
    .ZN(_00548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04951_ (.A1(_04208_),
    .A2(\mem[36][2] ),
    .ZN(_04211_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04952_ (.A1(_04138_),
    .A2(_04207_),
    .B(_04211_),
    .ZN(_00549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04953_ (.A1(_04208_),
    .A2(\mem[36][3] ),
    .ZN(_04212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04954_ (.A1(_04140_),
    .A2(_04207_),
    .B(_04212_),
    .ZN(_00550_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04955_ (.I(_04206_),
    .Z(_04213_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04956_ (.A1(_04213_),
    .A2(\mem[36][4] ),
    .ZN(_04214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04957_ (.A1(_04142_),
    .A2(_04207_),
    .B(_04214_),
    .ZN(_00551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04958_ (.A1(_04213_),
    .A2(\mem[36][5] ),
    .ZN(_04215_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04959_ (.A1(_04145_),
    .A2(_04207_),
    .B(_04215_),
    .ZN(_00552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04960_ (.A1(_04213_),
    .A2(\mem[36][6] ),
    .ZN(_04216_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04961_ (.A1(_04147_),
    .A2(_04207_),
    .B(_04216_),
    .ZN(_00553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04962_ (.A1(_04213_),
    .A2(\mem[36][7] ),
    .ZN(_04217_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04963_ (.A1(_04149_),
    .A2(_04207_),
    .B(_04217_),
    .ZN(_00554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04964_ (.A1(_04213_),
    .A2(\mem[36][8] ),
    .ZN(_04218_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04965_ (.A1(_04151_),
    .A2(_04207_),
    .B(_04218_),
    .ZN(_00555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04966_ (.A1(_04213_),
    .A2(\mem[36][9] ),
    .ZN(_04219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04967_ (.A1(_04153_),
    .A2(_04207_),
    .B(_04219_),
    .ZN(_00556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04968_ (.A1(_04213_),
    .A2(\mem[36][10] ),
    .ZN(_04220_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04969_ (.A1(_04155_),
    .A2(_04208_),
    .B(_04220_),
    .ZN(_00557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04970_ (.A1(_04213_),
    .A2(\mem[36][11] ),
    .ZN(_04221_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04971_ (.A1(_04157_),
    .A2(_04208_),
    .B(_04221_),
    .ZN(_00558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04972_ (.A1(_04213_),
    .A2(\mem[36][12] ),
    .ZN(_04222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04973_ (.A1(_04159_),
    .A2(_04208_),
    .B(_04222_),
    .ZN(_00559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04974_ (.A1(_04213_),
    .A2(\mem[36][13] ),
    .ZN(_04223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04975_ (.A1(_04125_),
    .A2(_04208_),
    .B(_04223_),
    .ZN(_00560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04976_ (.A1(_04206_),
    .A2(\mem[36][14] ),
    .ZN(_04224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04977_ (.A1(_04127_),
    .A2(_04208_),
    .B(_04224_),
    .ZN(_00561_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04978_ (.A1(_04206_),
    .A2(\mem[36][15] ),
    .ZN(_04225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04979_ (.A1(_04129_),
    .A2(_04208_),
    .B(_04225_),
    .ZN(_00562_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _04980_ (.A1(_03565_),
    .A2(_03440_),
    .ZN(_04226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _04981_ (.A1(_04226_),
    .A2(net76),
    .ZN(_04227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04982_ (.I(_04227_),
    .Z(_04228_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04983_ (.I(_04227_),
    .Z(_04229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04984_ (.A1(_04229_),
    .A2(\mem[37][0] ),
    .ZN(_04230_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04985_ (.A1(_04131_),
    .A2(_04228_),
    .B(_04230_),
    .ZN(_00563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04986_ (.A1(_04229_),
    .A2(\mem[37][1] ),
    .ZN(_04231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04987_ (.A1(_04136_),
    .A2(_04228_),
    .B(_04231_),
    .ZN(_00564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04988_ (.A1(_04229_),
    .A2(\mem[37][2] ),
    .ZN(_04232_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04989_ (.A1(_04138_),
    .A2(_04228_),
    .B(_04232_),
    .ZN(_00565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04990_ (.A1(_04229_),
    .A2(\mem[37][3] ),
    .ZN(_04233_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04991_ (.A1(_04140_),
    .A2(_04228_),
    .B(_04233_),
    .ZN(_00566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _04992_ (.I(_04227_),
    .Z(_04234_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04993_ (.A1(_04234_),
    .A2(\mem[37][4] ),
    .ZN(_04235_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04994_ (.A1(_04142_),
    .A2(_04228_),
    .B(_04235_),
    .ZN(_00567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04995_ (.A1(_04234_),
    .A2(\mem[37][5] ),
    .ZN(_04236_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04996_ (.A1(_04145_),
    .A2(_04228_),
    .B(_04236_),
    .ZN(_00568_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04997_ (.A1(_04234_),
    .A2(\mem[37][6] ),
    .ZN(_04237_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04998_ (.A1(_04147_),
    .A2(_04228_),
    .B(_04237_),
    .ZN(_00569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04999_ (.A1(_04234_),
    .A2(\mem[37][7] ),
    .ZN(_04238_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05000_ (.A1(_04149_),
    .A2(_04228_),
    .B(_04238_),
    .ZN(_00570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05001_ (.A1(_04234_),
    .A2(\mem[37][8] ),
    .ZN(_04239_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05002_ (.A1(_04151_),
    .A2(_04228_),
    .B(_04239_),
    .ZN(_00571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05003_ (.A1(_04234_),
    .A2(\mem[37][9] ),
    .ZN(_04240_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05004_ (.A1(_04153_),
    .A2(_04228_),
    .B(_04240_),
    .ZN(_00572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05005_ (.A1(_04234_),
    .A2(\mem[37][10] ),
    .ZN(_04241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05006_ (.A1(_04155_),
    .A2(_04229_),
    .B(_04241_),
    .ZN(_00573_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05007_ (.A1(_04234_),
    .A2(\mem[37][11] ),
    .ZN(_04242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05008_ (.A1(_04157_),
    .A2(_04229_),
    .B(_04242_),
    .ZN(_00574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05009_ (.A1(_04234_),
    .A2(\mem[37][12] ),
    .ZN(_04243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05010_ (.A1(_04159_),
    .A2(_04229_),
    .B(_04243_),
    .ZN(_00575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05011_ (.A1(_04234_),
    .A2(\mem[37][13] ),
    .ZN(_04244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05012_ (.A1(_04125_),
    .A2(_04229_),
    .B(_04244_),
    .ZN(_00576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05013_ (.A1(_04227_),
    .A2(\mem[37][14] ),
    .ZN(_04245_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05014_ (.A1(_04127_),
    .A2(_04229_),
    .B(_04245_),
    .ZN(_00577_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05015_ (.A1(_04227_),
    .A2(\mem[37][15] ),
    .ZN(_04246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05016_ (.A1(_04129_),
    .A2(_04229_),
    .B(_04246_),
    .ZN(_00578_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05017_ (.A1(net59),
    .A2(_01121_),
    .A3(_03440_),
    .ZN(_04247_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05018_ (.A1(_04247_),
    .A2(net76),
    .ZN(_04248_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05019_ (.I(_04248_),
    .Z(_04249_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05020_ (.I(_04248_),
    .Z(_04250_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05021_ (.A1(_04250_),
    .A2(\mem[38][0] ),
    .ZN(_04251_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05022_ (.A1(_04131_),
    .A2(_04249_),
    .B(_04251_),
    .ZN(_00579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05023_ (.A1(_04250_),
    .A2(\mem[38][1] ),
    .ZN(_04252_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05024_ (.A1(_04136_),
    .A2(_04249_),
    .B(_04252_),
    .ZN(_00580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05025_ (.A1(_04250_),
    .A2(\mem[38][2] ),
    .ZN(_04253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05026_ (.A1(_04138_),
    .A2(_04249_),
    .B(_04253_),
    .ZN(_00581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05027_ (.A1(_04250_),
    .A2(\mem[38][3] ),
    .ZN(_04254_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05028_ (.A1(_04140_),
    .A2(_04249_),
    .B(_04254_),
    .ZN(_00582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05029_ (.I(_04248_),
    .Z(_04255_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05030_ (.A1(_04255_),
    .A2(\mem[38][4] ),
    .ZN(_04256_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05031_ (.A1(_04142_),
    .A2(_04249_),
    .B(_04256_),
    .ZN(_00583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05032_ (.A1(_04255_),
    .A2(\mem[38][5] ),
    .ZN(_04257_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05033_ (.A1(_04145_),
    .A2(_04249_),
    .B(_04257_),
    .ZN(_00584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05034_ (.A1(_04255_),
    .A2(\mem[38][6] ),
    .ZN(_04258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05035_ (.A1(_04147_),
    .A2(_04249_),
    .B(_04258_),
    .ZN(_00585_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05036_ (.A1(_04255_),
    .A2(\mem[38][7] ),
    .ZN(_04259_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05037_ (.A1(_04149_),
    .A2(_04249_),
    .B(_04259_),
    .ZN(_00586_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05038_ (.A1(_04255_),
    .A2(\mem[38][8] ),
    .ZN(_04260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05039_ (.A1(_04151_),
    .A2(_04249_),
    .B(_04260_),
    .ZN(_00587_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05040_ (.A1(_04255_),
    .A2(\mem[38][9] ),
    .ZN(_04261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05041_ (.A1(_04153_),
    .A2(_04249_),
    .B(_04261_),
    .ZN(_00588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05042_ (.A1(_04255_),
    .A2(\mem[38][10] ),
    .ZN(_04262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05043_ (.A1(_04155_),
    .A2(_04250_),
    .B(_04262_),
    .ZN(_00589_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05044_ (.A1(_04255_),
    .A2(\mem[38][11] ),
    .ZN(_04263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05045_ (.A1(_04157_),
    .A2(_04250_),
    .B(_04263_),
    .ZN(_00590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05046_ (.A1(_04255_),
    .A2(\mem[38][12] ),
    .ZN(_04264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05047_ (.A1(_04159_),
    .A2(_04250_),
    .B(_04264_),
    .ZN(_00591_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05048_ (.A1(_04255_),
    .A2(\mem[38][13] ),
    .ZN(_04265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05049_ (.A1(_04125_),
    .A2(_04250_),
    .B(_04265_),
    .ZN(_00592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05050_ (.A1(_04248_),
    .A2(\mem[38][14] ),
    .ZN(_04266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05051_ (.A1(_04127_),
    .A2(_04250_),
    .B(_04266_),
    .ZN(_00593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05052_ (.A1(_04248_),
    .A2(\mem[38][15] ),
    .ZN(_04267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05053_ (.A1(_04129_),
    .A2(_04250_),
    .B(_04267_),
    .ZN(_00594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05054_ (.A1(_03522_),
    .A2(_03456_),
    .ZN(_04268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05055_ (.I(_04268_),
    .Z(_04269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05056_ (.I(_04268_),
    .Z(_04270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05057_ (.A1(_04270_),
    .A2(\mem[3][0] ),
    .ZN(_04271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05058_ (.A1(_04131_),
    .A2(_04269_),
    .B(_04271_),
    .ZN(_00595_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05059_ (.A1(_04270_),
    .A2(\mem[3][1] ),
    .ZN(_04272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05060_ (.A1(_04136_),
    .A2(_04269_),
    .B(_04272_),
    .ZN(_00596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05061_ (.A1(_04270_),
    .A2(\mem[3][2] ),
    .ZN(_04273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05062_ (.A1(_04138_),
    .A2(_04269_),
    .B(_04273_),
    .ZN(_00597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05063_ (.A1(_04270_),
    .A2(\mem[3][3] ),
    .ZN(_04274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05064_ (.A1(_04140_),
    .A2(_04269_),
    .B(_04274_),
    .ZN(_00598_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05065_ (.I(_04268_),
    .Z(_04275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05066_ (.A1(_04275_),
    .A2(\mem[3][4] ),
    .ZN(_04276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05067_ (.A1(_04142_),
    .A2(_04269_),
    .B(_04276_),
    .ZN(_00599_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05068_ (.A1(_04275_),
    .A2(\mem[3][5] ),
    .ZN(_04277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05069_ (.A1(_04145_),
    .A2(_04269_),
    .B(_04277_),
    .ZN(_00600_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05070_ (.A1(_04275_),
    .A2(\mem[3][6] ),
    .ZN(_04278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05071_ (.A1(_04147_),
    .A2(_04269_),
    .B(_04278_),
    .ZN(_00601_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05072_ (.A1(_04275_),
    .A2(\mem[3][7] ),
    .ZN(_04279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05073_ (.A1(_04149_),
    .A2(_04269_),
    .B(_04279_),
    .ZN(_00602_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05074_ (.A1(_04275_),
    .A2(\mem[3][8] ),
    .ZN(_04280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05075_ (.A1(_04151_),
    .A2(_04269_),
    .B(_04280_),
    .ZN(_00603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05076_ (.A1(_04275_),
    .A2(\mem[3][9] ),
    .ZN(_04281_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05077_ (.A1(_04153_),
    .A2(_04269_),
    .B(_04281_),
    .ZN(_00604_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05078_ (.A1(_04275_),
    .A2(\mem[3][10] ),
    .ZN(_04282_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05079_ (.A1(_04155_),
    .A2(_04270_),
    .B(_04282_),
    .ZN(_00605_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05080_ (.A1(_04275_),
    .A2(\mem[3][11] ),
    .ZN(_04283_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05081_ (.A1(_04157_),
    .A2(_04270_),
    .B(_04283_),
    .ZN(_00606_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05082_ (.A1(_04275_),
    .A2(\mem[3][12] ),
    .ZN(_04284_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05083_ (.A1(_04159_),
    .A2(_04270_),
    .B(_04284_),
    .ZN(_00607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05084_ (.A1(_04275_),
    .A2(\mem[3][13] ),
    .ZN(_04285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05085_ (.A1(_04125_),
    .A2(_04270_),
    .B(_04285_),
    .ZN(_00608_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05086_ (.A1(_04268_),
    .A2(\mem[3][14] ),
    .ZN(_04286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05087_ (.A1(_04127_),
    .A2(_04270_),
    .B(_04286_),
    .ZN(_00609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05088_ (.A1(_04268_),
    .A2(\mem[3][15] ),
    .ZN(_04287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05089_ (.A1(_04129_),
    .A2(_04270_),
    .B(_04287_),
    .ZN(_00610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05090_ (.A1(_01149_),
    .A2(_03588_),
    .ZN(_04288_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05091_ (.I(_04288_),
    .Z(_04289_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05092_ (.I(_04288_),
    .Z(_04290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05093_ (.A1(_04290_),
    .A2(\mem[40][0] ),
    .ZN(_04291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05094_ (.A1(_04131_),
    .A2(_04289_),
    .B(_04291_),
    .ZN(_00611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05095_ (.A1(_04290_),
    .A2(\mem[40][1] ),
    .ZN(_04292_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05096_ (.A1(_04136_),
    .A2(_04289_),
    .B(_04292_),
    .ZN(_00612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05097_ (.A1(_04290_),
    .A2(\mem[40][2] ),
    .ZN(_04293_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05098_ (.A1(_04138_),
    .A2(_04289_),
    .B(_04293_),
    .ZN(_00613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05099_ (.A1(_04290_),
    .A2(\mem[40][3] ),
    .ZN(_04294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05100_ (.A1(_04140_),
    .A2(_04289_),
    .B(_04294_),
    .ZN(_00614_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05101_ (.I(_04288_),
    .Z(_04295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05102_ (.A1(_04295_),
    .A2(\mem[40][4] ),
    .ZN(_04296_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05103_ (.A1(_04142_),
    .A2(_04289_),
    .B(_04296_),
    .ZN(_00615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05104_ (.A1(_04295_),
    .A2(\mem[40][5] ),
    .ZN(_04297_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05105_ (.A1(_04145_),
    .A2(_04289_),
    .B(_04297_),
    .ZN(_00616_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05106_ (.A1(_04295_),
    .A2(\mem[40][6] ),
    .ZN(_04298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05107_ (.A1(_04147_),
    .A2(_04289_),
    .B(_04298_),
    .ZN(_00617_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05108_ (.A1(_04295_),
    .A2(\mem[40][7] ),
    .ZN(_04299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05109_ (.A1(_04149_),
    .A2(_04289_),
    .B(_04299_),
    .ZN(_00618_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05110_ (.A1(_04295_),
    .A2(\mem[40][8] ),
    .ZN(_04300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05111_ (.A1(_04151_),
    .A2(_04289_),
    .B(_04300_),
    .ZN(_00619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05112_ (.A1(_04295_),
    .A2(\mem[40][9] ),
    .ZN(_04301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05113_ (.A1(_04153_),
    .A2(_04289_),
    .B(_04301_),
    .ZN(_00620_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05114_ (.A1(_04295_),
    .A2(\mem[40][10] ),
    .ZN(_04302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05115_ (.A1(_04155_),
    .A2(_04290_),
    .B(_04302_),
    .ZN(_00621_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05116_ (.A1(_04295_),
    .A2(\mem[40][11] ),
    .ZN(_04303_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05117_ (.A1(_04157_),
    .A2(_04290_),
    .B(_04303_),
    .ZN(_00622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05118_ (.A1(_04295_),
    .A2(\mem[40][12] ),
    .ZN(_04304_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05119_ (.A1(_04159_),
    .A2(_04290_),
    .B(_04304_),
    .ZN(_00623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05120_ (.A1(_04295_),
    .A2(\mem[40][13] ),
    .ZN(_04305_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05121_ (.A1(_04125_),
    .A2(_04290_),
    .B(_04305_),
    .ZN(_00624_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05122_ (.A1(_04288_),
    .A2(\mem[40][14] ),
    .ZN(_04306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05123_ (.A1(_04127_),
    .A2(_04290_),
    .B(_04306_),
    .ZN(_00625_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05124_ (.A1(_04288_),
    .A2(\mem[40][15] ),
    .ZN(_04307_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05125_ (.A1(_04129_),
    .A2(_04290_),
    .B(_04307_),
    .ZN(_00626_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05126_ (.A1(_01149_),
    .A2(net93),
    .ZN(_04308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05127_ (.I(_04308_),
    .Z(_04309_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05128_ (.I(_04308_),
    .Z(_04310_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05129_ (.A1(_04310_),
    .A2(\mem[41][0] ),
    .ZN(_04311_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05130_ (.A1(_04131_),
    .A2(_04309_),
    .B(_04311_),
    .ZN(_00627_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05131_ (.A1(_04310_),
    .A2(\mem[41][1] ),
    .ZN(_04312_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05132_ (.A1(_04136_),
    .A2(_04309_),
    .B(_04312_),
    .ZN(_00628_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05133_ (.A1(_04310_),
    .A2(\mem[41][2] ),
    .ZN(_04313_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05134_ (.A1(_04138_),
    .A2(_04309_),
    .B(_04313_),
    .ZN(_00629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05135_ (.A1(_04310_),
    .A2(\mem[41][3] ),
    .ZN(_04314_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05136_ (.A1(_04140_),
    .A2(_04309_),
    .B(_04314_),
    .ZN(_00630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05137_ (.I(_04308_),
    .Z(_04315_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05138_ (.A1(_04315_),
    .A2(\mem[41][4] ),
    .ZN(_04316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05139_ (.A1(_04142_),
    .A2(_04309_),
    .B(_04316_),
    .ZN(_00631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05140_ (.A1(_04315_),
    .A2(\mem[41][5] ),
    .ZN(_04317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05141_ (.A1(_04145_),
    .A2(_04309_),
    .B(_04317_),
    .ZN(_00632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05142_ (.A1(_04315_),
    .A2(\mem[41][6] ),
    .ZN(_04318_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05143_ (.A1(_04147_),
    .A2(_04309_),
    .B(_04318_),
    .ZN(_00633_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05144_ (.A1(_04315_),
    .A2(\mem[41][7] ),
    .ZN(_04319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05145_ (.A1(_04149_),
    .A2(_04309_),
    .B(_04319_),
    .ZN(_00634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05146_ (.A1(_04315_),
    .A2(\mem[41][8] ),
    .ZN(_04320_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05147_ (.A1(_04151_),
    .A2(_04309_),
    .B(_04320_),
    .ZN(_00635_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05148_ (.A1(_04315_),
    .A2(\mem[41][9] ),
    .ZN(_04321_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05149_ (.A1(_04153_),
    .A2(_04309_),
    .B(_04321_),
    .ZN(_00636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05150_ (.A1(_04315_),
    .A2(\mem[41][10] ),
    .ZN(_04322_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05151_ (.A1(_04155_),
    .A2(_04310_),
    .B(_04322_),
    .ZN(_00637_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05152_ (.A1(_04315_),
    .A2(\mem[41][11] ),
    .ZN(_04323_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05153_ (.A1(_04157_),
    .A2(_04310_),
    .B(_04323_),
    .ZN(_00638_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05154_ (.A1(_04315_),
    .A2(\mem[41][12] ),
    .ZN(_04324_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05155_ (.A1(_04159_),
    .A2(_04310_),
    .B(_04324_),
    .ZN(_00639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05156_ (.A1(_04315_),
    .A2(\mem[41][13] ),
    .ZN(_04325_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05157_ (.A1(_04125_),
    .A2(_04310_),
    .B(_04325_),
    .ZN(_00640_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05158_ (.A1(_04308_),
    .A2(\mem[41][14] ),
    .ZN(_04326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05159_ (.A1(_04127_),
    .A2(_04310_),
    .B(_04326_),
    .ZN(_00641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05160_ (.A1(_04308_),
    .A2(\mem[41][15] ),
    .ZN(_04327_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05161_ (.A1(_04129_),
    .A2(_04310_),
    .B(_04327_),
    .ZN(_00642_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05162_ (.A1(_04164_),
    .A2(_01148_),
    .ZN(_04328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05163_ (.I(_04328_),
    .Z(_04329_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05164_ (.I(_04328_),
    .Z(_04330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05165_ (.A1(_04330_),
    .A2(\mem[42][0] ),
    .ZN(_04331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05166_ (.A1(_04131_),
    .A2(_04329_),
    .B(_04331_),
    .ZN(_00643_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05167_ (.A1(_04330_),
    .A2(\mem[42][1] ),
    .ZN(_04332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05168_ (.A1(_04136_),
    .A2(_04329_),
    .B(_04332_),
    .ZN(_00644_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05169_ (.A1(_04330_),
    .A2(\mem[42][2] ),
    .ZN(_04333_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05170_ (.A1(_04138_),
    .A2(_04329_),
    .B(_04333_),
    .ZN(_00645_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05171_ (.A1(_04330_),
    .A2(\mem[42][3] ),
    .ZN(_04334_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05172_ (.A1(_04140_),
    .A2(_04329_),
    .B(_04334_),
    .ZN(_00646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05173_ (.I(_04328_),
    .Z(_04335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05174_ (.A1(_04335_),
    .A2(\mem[42][4] ),
    .ZN(_04336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05175_ (.A1(_04142_),
    .A2(_04329_),
    .B(_04336_),
    .ZN(_00647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05176_ (.A1(_04335_),
    .A2(\mem[42][5] ),
    .ZN(_04337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05177_ (.A1(_04145_),
    .A2(_04329_),
    .B(_04337_),
    .ZN(_00648_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05178_ (.A1(_04335_),
    .A2(\mem[42][6] ),
    .ZN(_04338_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05179_ (.A1(_04147_),
    .A2(_04329_),
    .B(_04338_),
    .ZN(_00649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05180_ (.A1(_04335_),
    .A2(\mem[42][7] ),
    .ZN(_04339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05181_ (.A1(_04149_),
    .A2(_04329_),
    .B(_04339_),
    .ZN(_00650_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05182_ (.A1(_04335_),
    .A2(\mem[42][8] ),
    .ZN(_04340_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05183_ (.A1(_04151_),
    .A2(_04329_),
    .B(_04340_),
    .ZN(_00651_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05184_ (.A1(_04335_),
    .A2(\mem[42][9] ),
    .ZN(_04341_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05185_ (.A1(_04153_),
    .A2(_04329_),
    .B(_04341_),
    .ZN(_00652_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05186_ (.A1(_04335_),
    .A2(\mem[42][10] ),
    .ZN(_04342_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05187_ (.A1(_04155_),
    .A2(_04330_),
    .B(_04342_),
    .ZN(_00653_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05188_ (.A1(_04335_),
    .A2(\mem[42][11] ),
    .ZN(_04343_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05189_ (.A1(_04157_),
    .A2(_04330_),
    .B(_04343_),
    .ZN(_00654_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05190_ (.A1(_04335_),
    .A2(\mem[42][12] ),
    .ZN(_04344_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05191_ (.A1(_04159_),
    .A2(_04330_),
    .B(_04344_),
    .ZN(_00655_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05192_ (.I(_03438_),
    .Z(_04345_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05193_ (.A1(_04335_),
    .A2(\mem[42][13] ),
    .ZN(_04346_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05194_ (.A1(_04345_),
    .A2(_04330_),
    .B(_04346_),
    .ZN(_00656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05195_ (.I(_03446_),
    .Z(_04347_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05196_ (.A1(_04328_),
    .A2(\mem[42][14] ),
    .ZN(_04348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05197_ (.A1(_04347_),
    .A2(_04330_),
    .B(_04348_),
    .ZN(_00657_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05198_ (.I(_03449_),
    .Z(_04349_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05199_ (.A1(_04328_),
    .A2(\mem[42][15] ),
    .ZN(_04350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05200_ (.A1(_04349_),
    .A2(_04330_),
    .B(_04350_),
    .ZN(_00658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05201_ (.I(_03452_),
    .Z(_04351_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05202_ (.A1(_03543_),
    .A2(_01148_),
    .ZN(_04352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05203_ (.I(_04352_),
    .Z(_04353_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05204_ (.I(_04352_),
    .Z(_04354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05205_ (.A1(_04354_),
    .A2(\mem[43][0] ),
    .ZN(_04355_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05206_ (.A1(_04351_),
    .A2(_04353_),
    .B(_04355_),
    .ZN(_00659_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05207_ (.I(_03461_),
    .Z(_04356_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05208_ (.A1(_04354_),
    .A2(\mem[43][1] ),
    .ZN(_04357_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05209_ (.A1(_04356_),
    .A2(_04353_),
    .B(_04357_),
    .ZN(_00660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05210_ (.I(_03464_),
    .Z(_04358_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05211_ (.A1(_04354_),
    .A2(\mem[43][2] ),
    .ZN(_04359_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05212_ (.A1(_04358_),
    .A2(_04353_),
    .B(_04359_),
    .ZN(_00661_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05213_ (.I(_03467_),
    .Z(_04360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05214_ (.A1(_04354_),
    .A2(\mem[43][3] ),
    .ZN(_04361_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05215_ (.A1(_04360_),
    .A2(_04353_),
    .B(_04361_),
    .ZN(_00662_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05216_ (.I(_03470_),
    .Z(_04362_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05217_ (.I(_04352_),
    .Z(_04363_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05218_ (.A1(_04363_),
    .A2(\mem[43][4] ),
    .ZN(_04364_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05219_ (.A1(_04362_),
    .A2(_04353_),
    .B(_04364_),
    .ZN(_00663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05220_ (.I(_03474_),
    .Z(_04365_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05221_ (.A1(_04363_),
    .A2(\mem[43][5] ),
    .ZN(_04366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05222_ (.A1(_04365_),
    .A2(_04353_),
    .B(_04366_),
    .ZN(_00664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05223_ (.I(_03477_),
    .Z(_04367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05224_ (.A1(_04363_),
    .A2(\mem[43][6] ),
    .ZN(_04368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05225_ (.A1(_04367_),
    .A2(_04353_),
    .B(_04368_),
    .ZN(_00665_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05226_ (.I(_03480_),
    .Z(_04369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05227_ (.A1(_04363_),
    .A2(\mem[43][7] ),
    .ZN(_04370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05228_ (.A1(_04369_),
    .A2(_04353_),
    .B(_04370_),
    .ZN(_00666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05229_ (.I(_03483_),
    .Z(_04371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05230_ (.A1(_04363_),
    .A2(\mem[43][8] ),
    .ZN(_04372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05231_ (.A1(_04371_),
    .A2(_04353_),
    .B(_04372_),
    .ZN(_00667_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05232_ (.I(_03486_),
    .Z(_04373_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05233_ (.A1(_04363_),
    .A2(\mem[43][9] ),
    .ZN(_04374_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05234_ (.A1(_04373_),
    .A2(_04353_),
    .B(_04374_),
    .ZN(_00668_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05235_ (.I(_03489_),
    .Z(_04375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05236_ (.A1(_04363_),
    .A2(\mem[43][10] ),
    .ZN(_04376_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05237_ (.A1(_04375_),
    .A2(_04354_),
    .B(_04376_),
    .ZN(_00669_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05238_ (.I(_03492_),
    .Z(_04377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05239_ (.A1(_04363_),
    .A2(\mem[43][11] ),
    .ZN(_04378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05240_ (.A1(_04377_),
    .A2(_04354_),
    .B(_04378_),
    .ZN(_00670_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05241_ (.I(_03495_),
    .Z(_04379_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05242_ (.A1(_04363_),
    .A2(\mem[43][12] ),
    .ZN(_04380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05243_ (.A1(_04379_),
    .A2(_04354_),
    .B(_04380_),
    .ZN(_00671_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05244_ (.A1(_04363_),
    .A2(\mem[43][13] ),
    .ZN(_04381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05245_ (.A1(_04345_),
    .A2(_04354_),
    .B(_04381_),
    .ZN(_00672_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05246_ (.A1(_04352_),
    .A2(\mem[43][14] ),
    .ZN(_04382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05247_ (.A1(_04347_),
    .A2(_04354_),
    .B(_04382_),
    .ZN(_00673_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05248_ (.A1(_04352_),
    .A2(\mem[43][15] ),
    .ZN(_04383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05249_ (.A1(_04349_),
    .A2(_04354_),
    .B(_04383_),
    .ZN(_00674_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05250_ (.A1(_04205_),
    .A2(_01148_),
    .ZN(_04384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05251_ (.I(_04384_),
    .Z(_04385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05252_ (.I(_04384_),
    .Z(_04386_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05253_ (.A1(_04386_),
    .A2(\mem[44][0] ),
    .ZN(_04387_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05254_ (.A1(_04351_),
    .A2(_04385_),
    .B(_04387_),
    .ZN(_00675_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05255_ (.A1(_04386_),
    .A2(\mem[44][1] ),
    .ZN(_04388_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05256_ (.A1(_04356_),
    .A2(_04385_),
    .B(_04388_),
    .ZN(_00676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05257_ (.A1(_04386_),
    .A2(\mem[44][2] ),
    .ZN(_04389_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05258_ (.A1(_04358_),
    .A2(_04385_),
    .B(_04389_),
    .ZN(_00677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05259_ (.A1(_04386_),
    .A2(\mem[44][3] ),
    .ZN(_04390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05260_ (.A1(_04360_),
    .A2(_04385_),
    .B(_04390_),
    .ZN(_00678_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05261_ (.I(_04384_),
    .Z(_04391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05262_ (.A1(_04391_),
    .A2(\mem[44][4] ),
    .ZN(_04392_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05263_ (.A1(_04362_),
    .A2(_04385_),
    .B(_04392_),
    .ZN(_00679_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05264_ (.A1(_04391_),
    .A2(\mem[44][5] ),
    .ZN(_04393_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05265_ (.A1(_04365_),
    .A2(_04385_),
    .B(_04393_),
    .ZN(_00680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05266_ (.A1(_04391_),
    .A2(\mem[44][6] ),
    .ZN(_04394_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05267_ (.A1(_04367_),
    .A2(_04385_),
    .B(_04394_),
    .ZN(_00681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05268_ (.A1(_04391_),
    .A2(\mem[44][7] ),
    .ZN(_04395_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05269_ (.A1(_04369_),
    .A2(_04385_),
    .B(_04395_),
    .ZN(_00682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05270_ (.A1(_04391_),
    .A2(\mem[44][8] ),
    .ZN(_04396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05271_ (.A1(_04371_),
    .A2(_04385_),
    .B(_04396_),
    .ZN(_00683_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05272_ (.A1(_04391_),
    .A2(\mem[44][9] ),
    .ZN(_04397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05273_ (.A1(_04373_),
    .A2(_04385_),
    .B(_04397_),
    .ZN(_00684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05274_ (.A1(_04391_),
    .A2(\mem[44][10] ),
    .ZN(_04398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05275_ (.A1(_04375_),
    .A2(_04386_),
    .B(_04398_),
    .ZN(_00685_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05276_ (.A1(_04391_),
    .A2(\mem[44][11] ),
    .ZN(_04399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05277_ (.A1(_04377_),
    .A2(_04386_),
    .B(_04399_),
    .ZN(_00686_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05278_ (.A1(_04391_),
    .A2(\mem[44][12] ),
    .ZN(_04400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05279_ (.A1(_04379_),
    .A2(_04386_),
    .B(_04400_),
    .ZN(_00687_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05280_ (.A1(_04391_),
    .A2(\mem[44][13] ),
    .ZN(_04401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05281_ (.A1(_04345_),
    .A2(_04386_),
    .B(_04401_),
    .ZN(_00688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05282_ (.A1(_04384_),
    .A2(\mem[44][14] ),
    .ZN(_04402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05283_ (.A1(_04347_),
    .A2(_04386_),
    .B(_04402_),
    .ZN(_00689_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05284_ (.A1(_04384_),
    .A2(\mem[44][15] ),
    .ZN(_04403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05285_ (.A1(_04349_),
    .A2(_04386_),
    .B(_04403_),
    .ZN(_00690_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05286_ (.A1(_04226_),
    .A2(_01148_),
    .ZN(_04404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05287_ (.I(_04404_),
    .Z(_04405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05288_ (.I(_04404_),
    .Z(_04406_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05289_ (.A1(_04406_),
    .A2(\mem[45][0] ),
    .ZN(_04407_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05290_ (.A1(_04351_),
    .A2(_04405_),
    .B(_04407_),
    .ZN(_00691_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05291_ (.A1(_04406_),
    .A2(\mem[45][1] ),
    .ZN(_04408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05292_ (.A1(_04356_),
    .A2(_04405_),
    .B(_04408_),
    .ZN(_00692_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05293_ (.A1(_04406_),
    .A2(\mem[45][2] ),
    .ZN(_04409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05294_ (.A1(_04358_),
    .A2(_04405_),
    .B(_04409_),
    .ZN(_00693_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05295_ (.A1(_04406_),
    .A2(\mem[45][3] ),
    .ZN(_04410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05296_ (.A1(_04360_),
    .A2(_04405_),
    .B(_04410_),
    .ZN(_00694_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05297_ (.I(_04404_),
    .Z(_04411_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05298_ (.A1(_04411_),
    .A2(\mem[45][4] ),
    .ZN(_04412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05299_ (.A1(_04362_),
    .A2(_04405_),
    .B(_04412_),
    .ZN(_00695_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05300_ (.A1(_04411_),
    .A2(\mem[45][5] ),
    .ZN(_04413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05301_ (.A1(_04365_),
    .A2(_04405_),
    .B(_04413_),
    .ZN(_00696_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05302_ (.A1(_04411_),
    .A2(\mem[45][6] ),
    .ZN(_04414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05303_ (.A1(_04367_),
    .A2(_04405_),
    .B(_04414_),
    .ZN(_00697_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05304_ (.A1(_04411_),
    .A2(\mem[45][7] ),
    .ZN(_04415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05305_ (.A1(_04369_),
    .A2(_04405_),
    .B(_04415_),
    .ZN(_00698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05306_ (.A1(_04411_),
    .A2(\mem[45][8] ),
    .ZN(_04416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05307_ (.A1(_04371_),
    .A2(_04405_),
    .B(_04416_),
    .ZN(_00699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05308_ (.A1(_04411_),
    .A2(\mem[45][9] ),
    .ZN(_04417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05309_ (.A1(_04373_),
    .A2(_04405_),
    .B(_04417_),
    .ZN(_00700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05310_ (.A1(_04411_),
    .A2(\mem[45][10] ),
    .ZN(_04418_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05311_ (.A1(_04375_),
    .A2(_04406_),
    .B(_04418_),
    .ZN(_00701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05312_ (.A1(_04411_),
    .A2(\mem[45][11] ),
    .ZN(_04419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05313_ (.A1(_04377_),
    .A2(_04406_),
    .B(_04419_),
    .ZN(_00702_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05314_ (.A1(_04411_),
    .A2(\mem[45][12] ),
    .ZN(_04420_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05315_ (.A1(_04379_),
    .A2(_04406_),
    .B(_04420_),
    .ZN(_00703_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05316_ (.A1(_04411_),
    .A2(\mem[45][13] ),
    .ZN(_04421_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05317_ (.A1(_04345_),
    .A2(_04406_),
    .B(_04421_),
    .ZN(_00704_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05318_ (.A1(_04404_),
    .A2(\mem[45][14] ),
    .ZN(_04422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05319_ (.A1(_04347_),
    .A2(_04406_),
    .B(_04422_),
    .ZN(_00705_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05320_ (.A1(_04404_),
    .A2(\mem[45][15] ),
    .ZN(_04423_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05321_ (.A1(_04349_),
    .A2(_04406_),
    .B(_04423_),
    .ZN(_00706_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05322_ (.A1(_01149_),
    .A2(_04247_),
    .ZN(_04424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05323_ (.I(_04424_),
    .Z(_04425_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05324_ (.I(_04424_),
    .Z(_04426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05325_ (.A1(_04426_),
    .A2(\mem[46][0] ),
    .ZN(_04427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05326_ (.A1(_04351_),
    .A2(_04425_),
    .B(_04427_),
    .ZN(_00707_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05327_ (.A1(_04426_),
    .A2(\mem[46][1] ),
    .ZN(_04428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05328_ (.A1(_04356_),
    .A2(_04425_),
    .B(_04428_),
    .ZN(_00708_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05329_ (.A1(_04426_),
    .A2(\mem[46][2] ),
    .ZN(_04429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05330_ (.A1(_04358_),
    .A2(_04425_),
    .B(_04429_),
    .ZN(_00709_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05331_ (.A1(_04426_),
    .A2(\mem[46][3] ),
    .ZN(_04430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05332_ (.A1(_04360_),
    .A2(_04425_),
    .B(_04430_),
    .ZN(_00710_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05333_ (.I(_04424_),
    .Z(_04431_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05334_ (.A1(_04431_),
    .A2(\mem[46][4] ),
    .ZN(_04432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05335_ (.A1(_04362_),
    .A2(_04425_),
    .B(_04432_),
    .ZN(_00711_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05336_ (.A1(_04431_),
    .A2(\mem[46][5] ),
    .ZN(_04433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05337_ (.A1(_04365_),
    .A2(_04425_),
    .B(_04433_),
    .ZN(_00712_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05338_ (.A1(_04431_),
    .A2(\mem[46][6] ),
    .ZN(_04434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05339_ (.A1(_04367_),
    .A2(_04425_),
    .B(_04434_),
    .ZN(_00713_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05340_ (.A1(_04431_),
    .A2(\mem[46][7] ),
    .ZN(_04435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05341_ (.A1(_04369_),
    .A2(_04425_),
    .B(_04435_),
    .ZN(_00714_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05342_ (.A1(_04431_),
    .A2(\mem[46][8] ),
    .ZN(_04436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05343_ (.A1(_04371_),
    .A2(_04425_),
    .B(_04436_),
    .ZN(_00715_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05344_ (.A1(_04431_),
    .A2(\mem[46][9] ),
    .ZN(_04437_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05345_ (.A1(_04373_),
    .A2(_04425_),
    .B(_04437_),
    .ZN(_00716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05346_ (.A1(_04431_),
    .A2(\mem[46][10] ),
    .ZN(_04438_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05347_ (.A1(_04375_),
    .A2(_04426_),
    .B(_04438_),
    .ZN(_00717_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05348_ (.A1(_04431_),
    .A2(\mem[46][11] ),
    .ZN(_04439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05349_ (.A1(_04377_),
    .A2(_04426_),
    .B(_04439_),
    .ZN(_00718_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05350_ (.A1(_04431_),
    .A2(\mem[46][12] ),
    .ZN(_04440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05351_ (.A1(_04379_),
    .A2(_04426_),
    .B(_04440_),
    .ZN(_00719_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05352_ (.A1(_04431_),
    .A2(\mem[46][13] ),
    .ZN(_04441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05353_ (.A1(_04345_),
    .A2(_04426_),
    .B(_04441_),
    .ZN(_00720_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05354_ (.A1(_04424_),
    .A2(\mem[46][14] ),
    .ZN(_04442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05355_ (.A1(_04347_),
    .A2(_04426_),
    .B(_04442_),
    .ZN(_00721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05356_ (.A1(_04424_),
    .A2(\mem[46][15] ),
    .ZN(_04443_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05357_ (.A1(_04349_),
    .A2(_04426_),
    .B(_04443_),
    .ZN(_00722_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05358_ (.A1(_01148_),
    .A2(net60),
    .ZN(_04444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05359_ (.I(_04444_),
    .Z(_04445_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05360_ (.I(_04444_),
    .Z(_04446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05361_ (.A1(_04446_),
    .A2(\mem[47][0] ),
    .ZN(_04447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05362_ (.A1(_04351_),
    .A2(_04445_),
    .B(_04447_),
    .ZN(_00723_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05363_ (.A1(_04446_),
    .A2(\mem[47][1] ),
    .ZN(_04448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05364_ (.A1(_04356_),
    .A2(_04445_),
    .B(_04448_),
    .ZN(_00724_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05365_ (.A1(_04446_),
    .A2(\mem[47][2] ),
    .ZN(_04449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05366_ (.A1(_04358_),
    .A2(_04445_),
    .B(_04449_),
    .ZN(_00725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05367_ (.A1(_04446_),
    .A2(\mem[47][3] ),
    .ZN(_04450_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05368_ (.A1(_04360_),
    .A2(_04445_),
    .B(_04450_),
    .ZN(_00726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05369_ (.I(_04444_),
    .Z(_04451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05370_ (.A1(_04451_),
    .A2(\mem[47][4] ),
    .ZN(_04452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05371_ (.A1(_04362_),
    .A2(_04445_),
    .B(_04452_),
    .ZN(_00727_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05372_ (.A1(_04451_),
    .A2(\mem[47][5] ),
    .ZN(_04453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05373_ (.A1(_04365_),
    .A2(_04445_),
    .B(_04453_),
    .ZN(_00728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05374_ (.A1(_04451_),
    .A2(\mem[47][6] ),
    .ZN(_04454_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05375_ (.A1(_04367_),
    .A2(_04445_),
    .B(_04454_),
    .ZN(_00729_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05376_ (.A1(_04451_),
    .A2(\mem[47][7] ),
    .ZN(_04455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05377_ (.A1(_04369_),
    .A2(_04445_),
    .B(_04455_),
    .ZN(_00730_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05378_ (.A1(_04451_),
    .A2(\mem[47][8] ),
    .ZN(_04456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05379_ (.A1(_04371_),
    .A2(_04445_),
    .B(_04456_),
    .ZN(_00731_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05380_ (.A1(_04451_),
    .A2(\mem[47][9] ),
    .ZN(_04457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05381_ (.A1(_04373_),
    .A2(_04445_),
    .B(_04457_),
    .ZN(_00732_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05382_ (.A1(_04451_),
    .A2(\mem[47][10] ),
    .ZN(_04458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05383_ (.A1(_04375_),
    .A2(_04446_),
    .B(_04458_),
    .ZN(_00733_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05384_ (.A1(_04451_),
    .A2(\mem[47][11] ),
    .ZN(_04459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05385_ (.A1(_04377_),
    .A2(_04446_),
    .B(_04459_),
    .ZN(_00734_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05386_ (.A1(_04451_),
    .A2(\mem[47][12] ),
    .ZN(_04460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05387_ (.A1(_04379_),
    .A2(_04446_),
    .B(_04460_),
    .ZN(_00735_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05388_ (.A1(_04451_),
    .A2(\mem[47][13] ),
    .ZN(_04461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05389_ (.A1(_04345_),
    .A2(_04446_),
    .B(_04461_),
    .ZN(_00736_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05390_ (.A1(_04444_),
    .A2(\mem[47][14] ),
    .ZN(_04462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05391_ (.A1(_04347_),
    .A2(_04446_),
    .B(_04462_),
    .ZN(_00737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05392_ (.A1(_04444_),
    .A2(\mem[47][15] ),
    .ZN(_04463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05393_ (.A1(_04349_),
    .A2(_04446_),
    .B(_04463_),
    .ZN(_00738_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05394_ (.A1(_03588_),
    .A2(_01330_),
    .ZN(_04464_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05395_ (.I(_04464_),
    .Z(_04465_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05396_ (.I(_04464_),
    .Z(_04466_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05397_ (.A1(_04466_),
    .A2(\mem[48][0] ),
    .ZN(_04467_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05398_ (.A1(_04351_),
    .A2(_04465_),
    .B(_04467_),
    .ZN(_00739_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05399_ (.A1(_04466_),
    .A2(\mem[48][1] ),
    .ZN(_04468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05400_ (.A1(_04356_),
    .A2(_04465_),
    .B(_04468_),
    .ZN(_00740_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05401_ (.A1(_04466_),
    .A2(\mem[48][2] ),
    .ZN(_04469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05402_ (.A1(_04358_),
    .A2(_04465_),
    .B(_04469_),
    .ZN(_00741_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05403_ (.A1(_04466_),
    .A2(\mem[48][3] ),
    .ZN(_04470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05404_ (.A1(_04360_),
    .A2(_04465_),
    .B(_04470_),
    .ZN(_00742_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05405_ (.I(_04464_),
    .Z(_04471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05406_ (.A1(_04471_),
    .A2(\mem[48][4] ),
    .ZN(_04472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05407_ (.A1(_04362_),
    .A2(_04465_),
    .B(_04472_),
    .ZN(_00743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05408_ (.A1(_04471_),
    .A2(\mem[48][5] ),
    .ZN(_04473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05409_ (.A1(_04365_),
    .A2(_04465_),
    .B(_04473_),
    .ZN(_00744_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05410_ (.A1(_04471_),
    .A2(\mem[48][6] ),
    .ZN(_04474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05411_ (.A1(_04367_),
    .A2(_04465_),
    .B(_04474_),
    .ZN(_00745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05412_ (.A1(_04471_),
    .A2(\mem[48][7] ),
    .ZN(_04475_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05413_ (.A1(_04369_),
    .A2(_04465_),
    .B(_04475_),
    .ZN(_00746_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05414_ (.A1(_04471_),
    .A2(\mem[48][8] ),
    .ZN(_04476_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05415_ (.A1(_04371_),
    .A2(_04465_),
    .B(_04476_),
    .ZN(_00747_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05416_ (.A1(_04471_),
    .A2(\mem[48][9] ),
    .ZN(_04477_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05417_ (.A1(_04373_),
    .A2(_04465_),
    .B(_04477_),
    .ZN(_00748_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05418_ (.A1(_04471_),
    .A2(\mem[48][10] ),
    .ZN(_04478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05419_ (.A1(_04375_),
    .A2(_04466_),
    .B(_04478_),
    .ZN(_00749_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05420_ (.A1(_04471_),
    .A2(\mem[48][11] ),
    .ZN(_04479_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05421_ (.A1(_04377_),
    .A2(_04466_),
    .B(_04479_),
    .ZN(_00750_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05422_ (.A1(_04471_),
    .A2(\mem[48][12] ),
    .ZN(_04480_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05423_ (.A1(_04379_),
    .A2(_04466_),
    .B(_04480_),
    .ZN(_00751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05424_ (.A1(_04471_),
    .A2(\mem[48][13] ),
    .ZN(_04481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05425_ (.A1(_04345_),
    .A2(_04466_),
    .B(_04481_),
    .ZN(_00752_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05426_ (.A1(_04464_),
    .A2(\mem[48][14] ),
    .ZN(_04482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05427_ (.A1(_04347_),
    .A2(_04466_),
    .B(_04482_),
    .ZN(_00753_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05428_ (.A1(_04464_),
    .A2(\mem[48][15] ),
    .ZN(_04483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05429_ (.A1(_04349_),
    .A2(_04466_),
    .B(_04483_),
    .ZN(_00754_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05430_ (.A1(_03522_),
    .A2(net132),
    .ZN(_04484_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05431_ (.I(_04484_),
    .Z(_04485_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05432_ (.I(_04484_),
    .Z(_04486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05433_ (.A1(_04486_),
    .A2(\mem[4][0] ),
    .ZN(_04487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05434_ (.A1(_04351_),
    .A2(_04485_),
    .B(_04487_),
    .ZN(_00755_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05435_ (.A1(_04486_),
    .A2(\mem[4][1] ),
    .ZN(_04488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05436_ (.A1(_04356_),
    .A2(_04485_),
    .B(_04488_),
    .ZN(_00756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05437_ (.A1(_04486_),
    .A2(\mem[4][2] ),
    .ZN(_04489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05438_ (.A1(_04358_),
    .A2(_04485_),
    .B(_04489_),
    .ZN(_00757_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05439_ (.A1(_04486_),
    .A2(\mem[4][3] ),
    .ZN(_04490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05440_ (.A1(_04360_),
    .A2(_04485_),
    .B(_04490_),
    .ZN(_00758_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05441_ (.I(_04484_),
    .Z(_04491_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05442_ (.A1(_04491_),
    .A2(\mem[4][4] ),
    .ZN(_04492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05443_ (.A1(_04362_),
    .A2(_04485_),
    .B(_04492_),
    .ZN(_00759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05444_ (.A1(_04491_),
    .A2(\mem[4][5] ),
    .ZN(_04493_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05445_ (.A1(_04365_),
    .A2(_04485_),
    .B(_04493_),
    .ZN(_00760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05446_ (.A1(_04491_),
    .A2(\mem[4][6] ),
    .ZN(_04494_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05447_ (.A1(_04367_),
    .A2(_04485_),
    .B(_04494_),
    .ZN(_00761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05448_ (.A1(_04491_),
    .A2(\mem[4][7] ),
    .ZN(_04495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05449_ (.A1(_04369_),
    .A2(_04485_),
    .B(_04495_),
    .ZN(_00762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05450_ (.A1(_04491_),
    .A2(\mem[4][8] ),
    .ZN(_04496_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05451_ (.A1(_04371_),
    .A2(_04485_),
    .B(_04496_),
    .ZN(_00763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05452_ (.A1(_04491_),
    .A2(\mem[4][9] ),
    .ZN(_04497_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05453_ (.A1(_04373_),
    .A2(_04485_),
    .B(_04497_),
    .ZN(_00764_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05454_ (.A1(_04491_),
    .A2(\mem[4][10] ),
    .ZN(_04498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05455_ (.A1(_04375_),
    .A2(_04486_),
    .B(_04498_),
    .ZN(_00765_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05456_ (.A1(_04491_),
    .A2(\mem[4][11] ),
    .ZN(_04499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05457_ (.A1(_04377_),
    .A2(_04486_),
    .B(_04499_),
    .ZN(_00766_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05458_ (.A1(_04491_),
    .A2(\mem[4][12] ),
    .ZN(_04500_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05459_ (.A1(_04379_),
    .A2(_04486_),
    .B(_04500_),
    .ZN(_00767_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05460_ (.A1(_04491_),
    .A2(\mem[4][13] ),
    .ZN(_04501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05461_ (.A1(_04345_),
    .A2(_04486_),
    .B(_04501_),
    .ZN(_00768_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05462_ (.A1(_04484_),
    .A2(\mem[4][14] ),
    .ZN(_04502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05463_ (.A1(_04347_),
    .A2(_04486_),
    .B(_04502_),
    .ZN(_00769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05464_ (.A1(_04484_),
    .A2(\mem[4][15] ),
    .ZN(_04503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05465_ (.A1(_04349_),
    .A2(_04486_),
    .B(_04503_),
    .ZN(_00770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05466_ (.A1(_04164_),
    .A2(_01330_),
    .ZN(_04504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05467_ (.I(_04504_),
    .Z(_04505_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05468_ (.I(_04504_),
    .Z(_04506_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05469_ (.A1(_04506_),
    .A2(\mem[50][0] ),
    .ZN(_04507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05470_ (.A1(_04351_),
    .A2(_04505_),
    .B(_04507_),
    .ZN(_00771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05471_ (.A1(_04506_),
    .A2(\mem[50][1] ),
    .ZN(_04508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05472_ (.A1(_04356_),
    .A2(_04505_),
    .B(_04508_),
    .ZN(_00772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05473_ (.A1(_04506_),
    .A2(\mem[50][2] ),
    .ZN(_04509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05474_ (.A1(_04358_),
    .A2(_04505_),
    .B(_04509_),
    .ZN(_00773_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05475_ (.A1(_04506_),
    .A2(\mem[50][3] ),
    .ZN(_04510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05476_ (.A1(_04360_),
    .A2(_04505_),
    .B(_04510_),
    .ZN(_00774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05477_ (.I(_04504_),
    .Z(_04511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05478_ (.A1(_04511_),
    .A2(\mem[50][4] ),
    .ZN(_04512_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05479_ (.A1(_04362_),
    .A2(_04505_),
    .B(_04512_),
    .ZN(_00775_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05480_ (.A1(_04511_),
    .A2(\mem[50][5] ),
    .ZN(_04513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05481_ (.A1(_04365_),
    .A2(_04505_),
    .B(_04513_),
    .ZN(_00776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05482_ (.A1(_04511_),
    .A2(\mem[50][6] ),
    .ZN(_04514_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05483_ (.A1(_04367_),
    .A2(_04505_),
    .B(_04514_),
    .ZN(_00777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05484_ (.A1(_04511_),
    .A2(\mem[50][7] ),
    .ZN(_04515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05485_ (.A1(_04369_),
    .A2(_04505_),
    .B(_04515_),
    .ZN(_00778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05486_ (.A1(_04511_),
    .A2(\mem[50][8] ),
    .ZN(_04516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05487_ (.A1(_04371_),
    .A2(_04505_),
    .B(_04516_),
    .ZN(_00779_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05488_ (.A1(_04511_),
    .A2(\mem[50][9] ),
    .ZN(_04517_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05489_ (.A1(_04373_),
    .A2(_04505_),
    .B(_04517_),
    .ZN(_00780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05490_ (.A1(_04511_),
    .A2(\mem[50][10] ),
    .ZN(_04518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05491_ (.A1(_04375_),
    .A2(_04506_),
    .B(_04518_),
    .ZN(_00781_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05492_ (.A1(_04511_),
    .A2(\mem[50][11] ),
    .ZN(_04519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05493_ (.A1(_04377_),
    .A2(_04506_),
    .B(_04519_),
    .ZN(_00782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05494_ (.A1(_04511_),
    .A2(\mem[50][12] ),
    .ZN(_04520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05495_ (.A1(_04379_),
    .A2(_04506_),
    .B(_04520_),
    .ZN(_00783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05496_ (.A1(_04511_),
    .A2(\mem[50][13] ),
    .ZN(_04521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05497_ (.A1(_04345_),
    .A2(_04506_),
    .B(_04521_),
    .ZN(_00784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05498_ (.A1(_04504_),
    .A2(\mem[50][14] ),
    .ZN(_04522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05499_ (.A1(_04347_),
    .A2(_04506_),
    .B(_04522_),
    .ZN(_00785_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05500_ (.A1(_04504_),
    .A2(\mem[50][15] ),
    .ZN(_04523_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05501_ (.A1(_04349_),
    .A2(_04506_),
    .B(_04523_),
    .ZN(_00786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05502_ (.A1(_03543_),
    .A2(_01330_),
    .ZN(_04524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05503_ (.I(_04524_),
    .Z(_04525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05504_ (.I(_04524_),
    .Z(_04526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05505_ (.A1(_04526_),
    .A2(\mem[51][0] ),
    .ZN(_04527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05506_ (.A1(_04351_),
    .A2(_04525_),
    .B(_04527_),
    .ZN(_00787_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05507_ (.A1(_04526_),
    .A2(\mem[51][1] ),
    .ZN(_04528_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05508_ (.A1(_04356_),
    .A2(_04525_),
    .B(_04528_),
    .ZN(_00788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05509_ (.A1(_04526_),
    .A2(\mem[51][2] ),
    .ZN(_04529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05510_ (.A1(_04358_),
    .A2(_04525_),
    .B(_04529_),
    .ZN(_00789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05511_ (.A1(_04526_),
    .A2(\mem[51][3] ),
    .ZN(_04530_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05512_ (.A1(_04360_),
    .A2(_04525_),
    .B(_04530_),
    .ZN(_00790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05513_ (.I(_04524_),
    .Z(_04531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05514_ (.A1(_04531_),
    .A2(\mem[51][4] ),
    .ZN(_04532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05515_ (.A1(_04362_),
    .A2(_04525_),
    .B(_04532_),
    .ZN(_00791_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05516_ (.A1(_04531_),
    .A2(\mem[51][5] ),
    .ZN(_04533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05517_ (.A1(_04365_),
    .A2(_04525_),
    .B(_04533_),
    .ZN(_00792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05518_ (.A1(_04531_),
    .A2(\mem[51][6] ),
    .ZN(_04534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05519_ (.A1(_04367_),
    .A2(_04525_),
    .B(_04534_),
    .ZN(_00793_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05520_ (.A1(_04531_),
    .A2(\mem[51][7] ),
    .ZN(_04535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05521_ (.A1(_04369_),
    .A2(_04525_),
    .B(_04535_),
    .ZN(_00794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05522_ (.A1(_04531_),
    .A2(\mem[51][8] ),
    .ZN(_04536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05523_ (.A1(_04371_),
    .A2(_04525_),
    .B(_04536_),
    .ZN(_00795_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05524_ (.A1(_04531_),
    .A2(\mem[51][9] ),
    .ZN(_04537_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05525_ (.A1(_04373_),
    .A2(_04525_),
    .B(_04537_),
    .ZN(_00796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05526_ (.A1(_04531_),
    .A2(\mem[51][10] ),
    .ZN(_04538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05527_ (.A1(_04375_),
    .A2(_04526_),
    .B(_04538_),
    .ZN(_00797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05528_ (.A1(_04531_),
    .A2(\mem[51][11] ),
    .ZN(_04539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05529_ (.A1(_04377_),
    .A2(_04526_),
    .B(_04539_),
    .ZN(_00798_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05530_ (.A1(_04531_),
    .A2(\mem[51][12] ),
    .ZN(_04540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05531_ (.A1(_04379_),
    .A2(_04526_),
    .B(_04540_),
    .ZN(_00799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05532_ (.A1(_04531_),
    .A2(\mem[51][13] ),
    .ZN(_04541_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05533_ (.A1(_04345_),
    .A2(_04526_),
    .B(_04541_),
    .ZN(_00800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05534_ (.A1(_04524_),
    .A2(\mem[51][14] ),
    .ZN(_04542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05535_ (.A1(_04347_),
    .A2(_04526_),
    .B(_04542_),
    .ZN(_00801_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05536_ (.A1(_04524_),
    .A2(\mem[51][15] ),
    .ZN(_04543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05537_ (.A1(_04349_),
    .A2(_04526_),
    .B(_04543_),
    .ZN(_00802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05538_ (.A1(_04205_),
    .A2(_01330_),
    .ZN(_04544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05539_ (.I(_04544_),
    .Z(_04545_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05540_ (.I(_04544_),
    .Z(_04546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05541_ (.A1(_04546_),
    .A2(\mem[52][0] ),
    .ZN(_04547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05542_ (.A1(_04351_),
    .A2(_04545_),
    .B(_04547_),
    .ZN(_00803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05543_ (.A1(_04546_),
    .A2(\mem[52][1] ),
    .ZN(_04548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05544_ (.A1(_04356_),
    .A2(_04545_),
    .B(_04548_),
    .ZN(_00804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05545_ (.A1(_04546_),
    .A2(\mem[52][2] ),
    .ZN(_04549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05546_ (.A1(_04358_),
    .A2(_04545_),
    .B(_04549_),
    .ZN(_00805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05547_ (.A1(_04546_),
    .A2(\mem[52][3] ),
    .ZN(_04550_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05548_ (.A1(_04360_),
    .A2(_04545_),
    .B(_04550_),
    .ZN(_00806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05549_ (.I(_04544_),
    .Z(_04551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05550_ (.A1(_04551_),
    .A2(\mem[52][4] ),
    .ZN(_04552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05551_ (.A1(_04362_),
    .A2(_04545_),
    .B(_04552_),
    .ZN(_00807_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05552_ (.A1(_04551_),
    .A2(\mem[52][5] ),
    .ZN(_04553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05553_ (.A1(_04365_),
    .A2(_04545_),
    .B(_04553_),
    .ZN(_00808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05554_ (.A1(_04551_),
    .A2(\mem[52][6] ),
    .ZN(_04554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05555_ (.A1(_04367_),
    .A2(_04545_),
    .B(_04554_),
    .ZN(_00809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05556_ (.A1(_04551_),
    .A2(\mem[52][7] ),
    .ZN(_04555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05557_ (.A1(_04369_),
    .A2(_04545_),
    .B(_04555_),
    .ZN(_00810_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05558_ (.A1(_04551_),
    .A2(\mem[52][8] ),
    .ZN(_04556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05559_ (.A1(_04371_),
    .A2(_04545_),
    .B(_04556_),
    .ZN(_00811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05560_ (.A1(_04551_),
    .A2(\mem[52][9] ),
    .ZN(_04557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05561_ (.A1(_04373_),
    .A2(_04545_),
    .B(_04557_),
    .ZN(_00812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05562_ (.A1(_04551_),
    .A2(\mem[52][10] ),
    .ZN(_04558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05563_ (.A1(_04375_),
    .A2(_04546_),
    .B(_04558_),
    .ZN(_00813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05564_ (.A1(_04551_),
    .A2(\mem[52][11] ),
    .ZN(_04559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05565_ (.A1(_04377_),
    .A2(_04546_),
    .B(_04559_),
    .ZN(_00814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05566_ (.A1(_04551_),
    .A2(\mem[52][12] ),
    .ZN(_04560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05567_ (.A1(_04379_),
    .A2(_04546_),
    .B(_04560_),
    .ZN(_00815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05568_ (.I(_03438_),
    .Z(_04561_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05569_ (.A1(_04551_),
    .A2(\mem[52][13] ),
    .ZN(_04562_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05570_ (.A1(_04561_),
    .A2(_04546_),
    .B(_04562_),
    .ZN(_00816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05571_ (.I(_03446_),
    .Z(_04563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05572_ (.A1(_04544_),
    .A2(\mem[52][14] ),
    .ZN(_04564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05573_ (.A1(_04563_),
    .A2(_04546_),
    .B(_04564_),
    .ZN(_00817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05574_ (.I(_03449_),
    .Z(_04565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05575_ (.A1(_04544_),
    .A2(\mem[52][15] ),
    .ZN(_04566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05576_ (.A1(_04565_),
    .A2(_04546_),
    .B(_04566_),
    .ZN(_00818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05577_ (.I(_03452_),
    .Z(_04567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05578_ (.A1(_04226_),
    .A2(net70),
    .ZN(_04568_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05579_ (.I(_04568_),
    .Z(_04569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05580_ (.I(_04568_),
    .Z(_04570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05581_ (.A1(_04570_),
    .A2(\mem[53][0] ),
    .ZN(_04571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05582_ (.A1(_04567_),
    .A2(_04569_),
    .B(_04571_),
    .ZN(_00819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05583_ (.I(_03461_),
    .Z(_04572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05584_ (.A1(_04570_),
    .A2(\mem[53][1] ),
    .ZN(_04573_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05585_ (.A1(_04572_),
    .A2(_04569_),
    .B(_04573_),
    .ZN(_00820_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05586_ (.I(_03464_),
    .Z(_04574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05587_ (.A1(_04570_),
    .A2(\mem[53][2] ),
    .ZN(_04575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05588_ (.A1(_04574_),
    .A2(_04569_),
    .B(_04575_),
    .ZN(_00821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05589_ (.I(_03467_),
    .Z(_04576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05590_ (.A1(_04570_),
    .A2(\mem[53][3] ),
    .ZN(_04577_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05591_ (.A1(_04576_),
    .A2(_04569_),
    .B(_04577_),
    .ZN(_00822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05592_ (.I(_03470_),
    .Z(_04578_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05593_ (.I(_04568_),
    .Z(_04579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05594_ (.A1(_04579_),
    .A2(\mem[53][4] ),
    .ZN(_04580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05595_ (.A1(_04578_),
    .A2(_04569_),
    .B(_04580_),
    .ZN(_00823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05596_ (.I(_03474_),
    .Z(_04581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05597_ (.A1(_04579_),
    .A2(\mem[53][5] ),
    .ZN(_04582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05598_ (.A1(_04581_),
    .A2(_04569_),
    .B(_04582_),
    .ZN(_00824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05599_ (.I(_03477_),
    .Z(_04583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05600_ (.A1(_04579_),
    .A2(\mem[53][6] ),
    .ZN(_04584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05601_ (.A1(_04583_),
    .A2(_04569_),
    .B(_04584_),
    .ZN(_00825_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05602_ (.I(_03480_),
    .Z(_04585_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05603_ (.A1(_04579_),
    .A2(\mem[53][7] ),
    .ZN(_04586_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05604_ (.A1(_04585_),
    .A2(_04569_),
    .B(_04586_),
    .ZN(_00826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05605_ (.I(_03483_),
    .Z(_04587_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05606_ (.A1(_04579_),
    .A2(\mem[53][8] ),
    .ZN(_04588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05607_ (.A1(_04587_),
    .A2(_04569_),
    .B(_04588_),
    .ZN(_00827_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05608_ (.I(_03486_),
    .Z(_04589_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05609_ (.A1(_04579_),
    .A2(\mem[53][9] ),
    .ZN(_04590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05610_ (.A1(_04589_),
    .A2(_04569_),
    .B(_04590_),
    .ZN(_00828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05611_ (.I(_03489_),
    .Z(_04591_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05612_ (.A1(_04579_),
    .A2(\mem[53][10] ),
    .ZN(_04592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05613_ (.A1(_04591_),
    .A2(_04570_),
    .B(_04592_),
    .ZN(_00829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05614_ (.I(_03492_),
    .Z(_04593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05615_ (.A1(_04579_),
    .A2(\mem[53][11] ),
    .ZN(_04594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05616_ (.A1(_04593_),
    .A2(_04570_),
    .B(_04594_),
    .ZN(_00830_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05617_ (.I(_03495_),
    .Z(_04595_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05618_ (.A1(_04579_),
    .A2(\mem[53][12] ),
    .ZN(_04596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05619_ (.A1(_04595_),
    .A2(_04570_),
    .B(_04596_),
    .ZN(_00831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05620_ (.A1(_04579_),
    .A2(\mem[53][13] ),
    .ZN(_04597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05621_ (.A1(_04561_),
    .A2(_04570_),
    .B(_04597_),
    .ZN(_00832_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05622_ (.A1(_04568_),
    .A2(\mem[53][14] ),
    .ZN(_04598_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05623_ (.A1(_04563_),
    .A2(_04570_),
    .B(_04598_),
    .ZN(_00833_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05624_ (.A1(_04568_),
    .A2(\mem[53][15] ),
    .ZN(_04599_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05625_ (.A1(_04565_),
    .A2(_04570_),
    .B(_04599_),
    .ZN(_00834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05626_ (.A1(_04247_),
    .A2(net70),
    .ZN(_04600_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05627_ (.I(_04600_),
    .Z(_04601_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05628_ (.I(_04600_),
    .Z(_04602_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05629_ (.A1(_04602_),
    .A2(\mem[54][0] ),
    .ZN(_04603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05630_ (.A1(_04567_),
    .A2(_04601_),
    .B(_04603_),
    .ZN(_00835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05631_ (.A1(_04602_),
    .A2(\mem[54][1] ),
    .ZN(_04604_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05632_ (.A1(_04572_),
    .A2(_04601_),
    .B(_04604_),
    .ZN(_00836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05633_ (.A1(_04602_),
    .A2(\mem[54][2] ),
    .ZN(_04605_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05634_ (.A1(_04574_),
    .A2(_04601_),
    .B(_04605_),
    .ZN(_00837_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05635_ (.A1(_04602_),
    .A2(\mem[54][3] ),
    .ZN(_04606_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05636_ (.A1(_04576_),
    .A2(_04601_),
    .B(_04606_),
    .ZN(_00838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05637_ (.I(_04600_),
    .Z(_04607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05638_ (.A1(_04607_),
    .A2(\mem[54][4] ),
    .ZN(_04608_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05639_ (.A1(_04578_),
    .A2(_04601_),
    .B(_04608_),
    .ZN(_00839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05640_ (.A1(_04607_),
    .A2(\mem[54][5] ),
    .ZN(_04609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05641_ (.A1(_04581_),
    .A2(_04601_),
    .B(_04609_),
    .ZN(_00840_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05642_ (.A1(_04607_),
    .A2(\mem[54][6] ),
    .ZN(_04610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05643_ (.A1(_04583_),
    .A2(_04601_),
    .B(_04610_),
    .ZN(_00841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05644_ (.A1(_04607_),
    .A2(\mem[54][7] ),
    .ZN(_04611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05645_ (.A1(_04585_),
    .A2(_04601_),
    .B(_04611_),
    .ZN(_00842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05646_ (.A1(_04607_),
    .A2(\mem[54][8] ),
    .ZN(_04612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05647_ (.A1(_04587_),
    .A2(_04601_),
    .B(_04612_),
    .ZN(_00843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05648_ (.A1(_04607_),
    .A2(\mem[54][9] ),
    .ZN(_04613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05649_ (.A1(_04589_),
    .A2(_04601_),
    .B(_04613_),
    .ZN(_00844_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05650_ (.A1(_04607_),
    .A2(\mem[54][10] ),
    .ZN(_04614_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05651_ (.A1(_04591_),
    .A2(_04602_),
    .B(_04614_),
    .ZN(_00845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05652_ (.A1(_04607_),
    .A2(\mem[54][11] ),
    .ZN(_04615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05653_ (.A1(_04593_),
    .A2(_04602_),
    .B(_04615_),
    .ZN(_00846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05654_ (.A1(_04607_),
    .A2(\mem[54][12] ),
    .ZN(_04616_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05655_ (.A1(_04595_),
    .A2(_04602_),
    .B(_04616_),
    .ZN(_00847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05656_ (.A1(_04607_),
    .A2(\mem[54][13] ),
    .ZN(_04617_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05657_ (.A1(_04561_),
    .A2(_04602_),
    .B(_04617_),
    .ZN(_00848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05658_ (.A1(_04600_),
    .A2(\mem[54][14] ),
    .ZN(_04618_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05659_ (.A1(_04563_),
    .A2(_04602_),
    .B(_04618_),
    .ZN(_00849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05660_ (.A1(_04600_),
    .A2(\mem[54][15] ),
    .ZN(_04619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05661_ (.A1(_04565_),
    .A2(_04602_),
    .B(_04619_),
    .ZN(_00850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05662_ (.A1(net60),
    .A2(net70),
    .ZN(_04620_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05663_ (.I(_04620_),
    .Z(_04621_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05664_ (.I(_04620_),
    .Z(_04622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05665_ (.A1(_04622_),
    .A2(\mem[55][0] ),
    .ZN(_04623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05666_ (.A1(_04567_),
    .A2(_04621_),
    .B(_04623_),
    .ZN(_00851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05667_ (.A1(_04622_),
    .A2(\mem[55][1] ),
    .ZN(_04624_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05668_ (.A1(_04572_),
    .A2(_04621_),
    .B(_04624_),
    .ZN(_00852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05669_ (.A1(_04622_),
    .A2(\mem[55][2] ),
    .ZN(_04625_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05670_ (.A1(_04574_),
    .A2(_04621_),
    .B(_04625_),
    .ZN(_00853_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05671_ (.A1(_04622_),
    .A2(\mem[55][3] ),
    .ZN(_04626_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05672_ (.A1(_04576_),
    .A2(_04621_),
    .B(_04626_),
    .ZN(_00854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05673_ (.I(_04620_),
    .Z(_04627_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05674_ (.A1(_04627_),
    .A2(\mem[55][4] ),
    .ZN(_04628_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05675_ (.A1(_04578_),
    .A2(_04621_),
    .B(_04628_),
    .ZN(_00855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05676_ (.A1(_04627_),
    .A2(\mem[55][5] ),
    .ZN(_04629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05677_ (.A1(_04581_),
    .A2(_04621_),
    .B(_04629_),
    .ZN(_00856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05678_ (.A1(_04627_),
    .A2(\mem[55][6] ),
    .ZN(_04630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05679_ (.A1(_04583_),
    .A2(_04621_),
    .B(_04630_),
    .ZN(_00857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05680_ (.A1(_04627_),
    .A2(\mem[55][7] ),
    .ZN(_04631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05681_ (.A1(_04585_),
    .A2(_04621_),
    .B(_04631_),
    .ZN(_00858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05682_ (.A1(_04627_),
    .A2(\mem[55][8] ),
    .ZN(_04632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05683_ (.A1(_04587_),
    .A2(_04621_),
    .B(_04632_),
    .ZN(_00859_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05684_ (.A1(_04627_),
    .A2(\mem[55][9] ),
    .ZN(_04633_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05685_ (.A1(_04589_),
    .A2(_04621_),
    .B(_04633_),
    .ZN(_00860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05686_ (.A1(_04627_),
    .A2(\mem[55][10] ),
    .ZN(_04634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05687_ (.A1(_04591_),
    .A2(_04622_),
    .B(_04634_),
    .ZN(_00861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05688_ (.A1(_04627_),
    .A2(\mem[55][11] ),
    .ZN(_04635_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05689_ (.A1(_04593_),
    .A2(_04622_),
    .B(_04635_),
    .ZN(_00862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05690_ (.A1(_04627_),
    .A2(\mem[55][12] ),
    .ZN(_04636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05691_ (.A1(_04595_),
    .A2(_04622_),
    .B(_04636_),
    .ZN(_00863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05692_ (.A1(_04627_),
    .A2(\mem[55][13] ),
    .ZN(_04637_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05693_ (.A1(_04561_),
    .A2(_04622_),
    .B(_04637_),
    .ZN(_00864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05694_ (.A1(_04620_),
    .A2(\mem[55][14] ),
    .ZN(_04638_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05695_ (.A1(_04563_),
    .A2(_04622_),
    .B(_04638_),
    .ZN(_00865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05696_ (.A1(_04620_),
    .A2(\mem[55][15] ),
    .ZN(_04639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05697_ (.A1(_04565_),
    .A2(_04622_),
    .B(_04639_),
    .ZN(_00866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05698_ (.A1(_03588_),
    .A2(_01364_),
    .ZN(_04640_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05699_ (.I(_04640_),
    .Z(_04641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05700_ (.I(_04640_),
    .Z(_04642_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05701_ (.A1(_04642_),
    .A2(\mem[56][0] ),
    .ZN(_04643_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05702_ (.A1(_04567_),
    .A2(_04641_),
    .B(_04643_),
    .ZN(_00867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05703_ (.A1(_04642_),
    .A2(\mem[56][1] ),
    .ZN(_04644_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05704_ (.A1(_04572_),
    .A2(_04641_),
    .B(_04644_),
    .ZN(_00868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05705_ (.A1(_04642_),
    .A2(\mem[56][2] ),
    .ZN(_04645_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05706_ (.A1(_04574_),
    .A2(_04641_),
    .B(_04645_),
    .ZN(_00869_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05707_ (.A1(_04642_),
    .A2(\mem[56][3] ),
    .ZN(_04646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05708_ (.A1(_04576_),
    .A2(_04641_),
    .B(_04646_),
    .ZN(_00870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05709_ (.I(_04640_),
    .Z(_04647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05710_ (.A1(_04647_),
    .A2(\mem[56][4] ),
    .ZN(_04648_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05711_ (.A1(_04578_),
    .A2(_04641_),
    .B(_04648_),
    .ZN(_00871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05712_ (.A1(_04647_),
    .A2(\mem[56][5] ),
    .ZN(_04649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05713_ (.A1(_04581_),
    .A2(_04641_),
    .B(_04649_),
    .ZN(_00872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05714_ (.A1(_04647_),
    .A2(\mem[56][6] ),
    .ZN(_04650_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05715_ (.A1(_04583_),
    .A2(_04641_),
    .B(_04650_),
    .ZN(_00873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05716_ (.A1(_04647_),
    .A2(\mem[56][7] ),
    .ZN(_04651_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05717_ (.A1(_04585_),
    .A2(_04641_),
    .B(_04651_),
    .ZN(_00874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05718_ (.A1(_04647_),
    .A2(\mem[56][8] ),
    .ZN(_04652_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05719_ (.A1(_04587_),
    .A2(_04641_),
    .B(_04652_),
    .ZN(_00875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05720_ (.A1(_04647_),
    .A2(\mem[56][9] ),
    .ZN(_04653_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05721_ (.A1(_04589_),
    .A2(_04641_),
    .B(_04653_),
    .ZN(_00876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05722_ (.A1(_04647_),
    .A2(\mem[56][10] ),
    .ZN(_04654_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05723_ (.A1(_04591_),
    .A2(_04642_),
    .B(_04654_),
    .ZN(_00877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05724_ (.A1(_04647_),
    .A2(\mem[56][11] ),
    .ZN(_04655_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05725_ (.A1(_04593_),
    .A2(_04642_),
    .B(_04655_),
    .ZN(_00878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05726_ (.A1(_04647_),
    .A2(\mem[56][12] ),
    .ZN(_04656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05727_ (.A1(_04595_),
    .A2(_04642_),
    .B(_04656_),
    .ZN(_00879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05728_ (.A1(_04647_),
    .A2(\mem[56][13] ),
    .ZN(_04657_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05729_ (.A1(_04561_),
    .A2(_04642_),
    .B(_04657_),
    .ZN(_00880_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05730_ (.A1(_04640_),
    .A2(\mem[56][14] ),
    .ZN(_04658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05731_ (.A1(_04563_),
    .A2(_04642_),
    .B(_04658_),
    .ZN(_00881_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05732_ (.A1(_04640_),
    .A2(\mem[56][15] ),
    .ZN(_04659_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05733_ (.A1(_04565_),
    .A2(_04642_),
    .B(_04659_),
    .ZN(_00882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05734_ (.A1(net93),
    .A2(_01364_),
    .ZN(_04660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05735_ (.I(_04660_),
    .Z(_04661_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05736_ (.I(_04660_),
    .Z(_04662_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05737_ (.A1(_04662_),
    .A2(\mem[57][0] ),
    .ZN(_04663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05738_ (.A1(_04567_),
    .A2(_04661_),
    .B(_04663_),
    .ZN(_00883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05739_ (.A1(_04662_),
    .A2(\mem[57][1] ),
    .ZN(_04664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05740_ (.A1(_04572_),
    .A2(_04661_),
    .B(_04664_),
    .ZN(_00884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05741_ (.A1(_04662_),
    .A2(\mem[57][2] ),
    .ZN(_04665_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05742_ (.A1(_04574_),
    .A2(_04661_),
    .B(_04665_),
    .ZN(_00885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05743_ (.A1(_04662_),
    .A2(\mem[57][3] ),
    .ZN(_04666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05744_ (.A1(_04576_),
    .A2(_04661_),
    .B(_04666_),
    .ZN(_00886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05745_ (.I(_04660_),
    .Z(_04667_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05746_ (.A1(_04667_),
    .A2(\mem[57][4] ),
    .ZN(_04668_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05747_ (.A1(_04578_),
    .A2(_04661_),
    .B(_04668_),
    .ZN(_00887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05748_ (.A1(_04667_),
    .A2(\mem[57][5] ),
    .ZN(_04669_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05749_ (.A1(_04581_),
    .A2(_04661_),
    .B(_04669_),
    .ZN(_00888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05750_ (.A1(_04667_),
    .A2(\mem[57][6] ),
    .ZN(_04670_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05751_ (.A1(_04583_),
    .A2(_04661_),
    .B(_04670_),
    .ZN(_00889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05752_ (.A1(_04667_),
    .A2(\mem[57][7] ),
    .ZN(_04671_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05753_ (.A1(_04585_),
    .A2(_04661_),
    .B(_04671_),
    .ZN(_00890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05754_ (.A1(_04667_),
    .A2(\mem[57][8] ),
    .ZN(_04672_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05755_ (.A1(_04587_),
    .A2(_04661_),
    .B(_04672_),
    .ZN(_00891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05756_ (.A1(_04667_),
    .A2(\mem[57][9] ),
    .ZN(_04673_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05757_ (.A1(_04589_),
    .A2(_04661_),
    .B(_04673_),
    .ZN(_00892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05758_ (.A1(_04667_),
    .A2(\mem[57][10] ),
    .ZN(_04674_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05759_ (.A1(_04591_),
    .A2(_04662_),
    .B(_04674_),
    .ZN(_00893_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05760_ (.A1(_04667_),
    .A2(\mem[57][11] ),
    .ZN(_04675_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05761_ (.A1(_04593_),
    .A2(_04662_),
    .B(_04675_),
    .ZN(_00894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05762_ (.A1(_04667_),
    .A2(\mem[57][12] ),
    .ZN(_04676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05763_ (.A1(_04595_),
    .A2(_04662_),
    .B(_04676_),
    .ZN(_00895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05764_ (.A1(_04667_),
    .A2(\mem[57][13] ),
    .ZN(_04677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05765_ (.A1(_04561_),
    .A2(_04662_),
    .B(_04677_),
    .ZN(_00896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05766_ (.A1(_04660_),
    .A2(\mem[57][14] ),
    .ZN(_04678_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05767_ (.A1(_04563_),
    .A2(_04662_),
    .B(_04678_),
    .ZN(_00897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05768_ (.A1(_04660_),
    .A2(\mem[57][15] ),
    .ZN(_04679_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05769_ (.A1(_04565_),
    .A2(_04662_),
    .B(_04679_),
    .ZN(_00898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05770_ (.A1(net88),
    .A2(_03632_),
    .ZN(_04680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05771_ (.I(_04680_),
    .Z(_04681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05772_ (.I(_04680_),
    .Z(_04682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05773_ (.A1(_04682_),
    .A2(\mem[58][0] ),
    .ZN(_04683_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05774_ (.A1(_04567_),
    .A2(_04681_),
    .B(_04683_),
    .ZN(_00899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05775_ (.A1(_04682_),
    .A2(\mem[58][1] ),
    .ZN(_04684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05776_ (.A1(_04572_),
    .A2(_04681_),
    .B(_04684_),
    .ZN(_00900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05777_ (.A1(_04682_),
    .A2(\mem[58][2] ),
    .ZN(_04685_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05778_ (.A1(_04574_),
    .A2(_04681_),
    .B(_04685_),
    .ZN(_00901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05779_ (.A1(_04682_),
    .A2(\mem[58][3] ),
    .ZN(_04686_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05780_ (.A1(_04576_),
    .A2(_04681_),
    .B(_04686_),
    .ZN(_00902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05781_ (.I(_04680_),
    .Z(_04687_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05782_ (.A1(_04687_),
    .A2(\mem[58][4] ),
    .ZN(_04688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05783_ (.A1(_04578_),
    .A2(_04681_),
    .B(_04688_),
    .ZN(_00903_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05784_ (.A1(_04687_),
    .A2(\mem[58][5] ),
    .ZN(_04689_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05785_ (.A1(_04581_),
    .A2(_04681_),
    .B(_04689_),
    .ZN(_00904_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05786_ (.A1(_04687_),
    .A2(\mem[58][6] ),
    .ZN(_04690_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05787_ (.A1(_04583_),
    .A2(_04681_),
    .B(_04690_),
    .ZN(_00905_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05788_ (.A1(_04687_),
    .A2(\mem[58][7] ),
    .ZN(_04691_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05789_ (.A1(_04585_),
    .A2(_04681_),
    .B(_04691_),
    .ZN(_00906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05790_ (.A1(_04687_),
    .A2(\mem[58][8] ),
    .ZN(_04692_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05791_ (.A1(_04587_),
    .A2(_04681_),
    .B(_04692_),
    .ZN(_00907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05792_ (.A1(_04687_),
    .A2(\mem[58][9] ),
    .ZN(_04693_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05793_ (.A1(_04589_),
    .A2(_04681_),
    .B(_04693_),
    .ZN(_00908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05794_ (.A1(_04687_),
    .A2(\mem[58][10] ),
    .ZN(_04694_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05795_ (.A1(_04591_),
    .A2(_04682_),
    .B(_04694_),
    .ZN(_00909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05796_ (.A1(_04687_),
    .A2(\mem[58][11] ),
    .ZN(_04695_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05797_ (.A1(_04593_),
    .A2(_04682_),
    .B(_04695_),
    .ZN(_00910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05798_ (.A1(_04687_),
    .A2(\mem[58][12] ),
    .ZN(_04696_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05799_ (.A1(_04595_),
    .A2(_04682_),
    .B(_04696_),
    .ZN(_00911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05800_ (.A1(_04687_),
    .A2(\mem[58][13] ),
    .ZN(_04697_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05801_ (.A1(_04561_),
    .A2(_04682_),
    .B(_04697_),
    .ZN(_00912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05802_ (.A1(_04680_),
    .A2(\mem[58][14] ),
    .ZN(_04698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05803_ (.A1(_04563_),
    .A2(_04682_),
    .B(_04698_),
    .ZN(_00913_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05804_ (.A1(_04680_),
    .A2(\mem[58][15] ),
    .ZN(_04699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05805_ (.A1(_04565_),
    .A2(_04682_),
    .B(_04699_),
    .ZN(_00914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05806_ (.A1(_03522_),
    .A2(_03566_),
    .ZN(_04700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05807_ (.I(_04700_),
    .Z(_04701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05808_ (.I(_04700_),
    .Z(_04702_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05809_ (.A1(_04702_),
    .A2(\mem[5][0] ),
    .ZN(_04703_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05810_ (.A1(_04567_),
    .A2(_04701_),
    .B(_04703_),
    .ZN(_00915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05811_ (.A1(_04702_),
    .A2(\mem[5][1] ),
    .ZN(_04704_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05812_ (.A1(_04572_),
    .A2(_04701_),
    .B(_04704_),
    .ZN(_00916_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05813_ (.A1(_04702_),
    .A2(\mem[5][2] ),
    .ZN(_04705_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05814_ (.A1(_04574_),
    .A2(_04701_),
    .B(_04705_),
    .ZN(_00917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05815_ (.A1(_04702_),
    .A2(\mem[5][3] ),
    .ZN(_04706_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05816_ (.A1(_04576_),
    .A2(_04701_),
    .B(_04706_),
    .ZN(_00918_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05817_ (.I(_04700_),
    .Z(_04707_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05818_ (.A1(_04707_),
    .A2(\mem[5][4] ),
    .ZN(_04708_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05819_ (.A1(_04578_),
    .A2(_04701_),
    .B(_04708_),
    .ZN(_00919_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05820_ (.A1(_04707_),
    .A2(\mem[5][5] ),
    .ZN(_04709_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05821_ (.A1(_04581_),
    .A2(_04701_),
    .B(_04709_),
    .ZN(_00920_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05822_ (.A1(_04707_),
    .A2(\mem[5][6] ),
    .ZN(_04710_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05823_ (.A1(_04583_),
    .A2(_04701_),
    .B(_04710_),
    .ZN(_00921_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05824_ (.A1(_04707_),
    .A2(\mem[5][7] ),
    .ZN(_04711_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05825_ (.A1(_04585_),
    .A2(_04701_),
    .B(_04711_),
    .ZN(_00922_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05826_ (.A1(_04707_),
    .A2(\mem[5][8] ),
    .ZN(_04712_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05827_ (.A1(_04587_),
    .A2(_04701_),
    .B(_04712_),
    .ZN(_00923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05828_ (.A1(_04707_),
    .A2(\mem[5][9] ),
    .ZN(_04713_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05829_ (.A1(_04589_),
    .A2(_04701_),
    .B(_04713_),
    .ZN(_00924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05830_ (.A1(_04707_),
    .A2(\mem[5][10] ),
    .ZN(_04714_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05831_ (.A1(_04591_),
    .A2(_04702_),
    .B(_04714_),
    .ZN(_00925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05832_ (.A1(_04707_),
    .A2(\mem[5][11] ),
    .ZN(_04715_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05833_ (.A1(_04593_),
    .A2(_04702_),
    .B(_04715_),
    .ZN(_00926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05834_ (.A1(_04707_),
    .A2(\mem[5][12] ),
    .ZN(_04716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05835_ (.A1(_04595_),
    .A2(_04702_),
    .B(_04716_),
    .ZN(_00927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05836_ (.A1(_04707_),
    .A2(\mem[5][13] ),
    .ZN(_04717_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05837_ (.A1(_04561_),
    .A2(_04702_),
    .B(_04717_),
    .ZN(_00928_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05838_ (.A1(_04700_),
    .A2(\mem[5][14] ),
    .ZN(_04718_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05839_ (.A1(_04563_),
    .A2(_04702_),
    .B(_04718_),
    .ZN(_00929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05840_ (.A1(_04700_),
    .A2(\mem[5][15] ),
    .ZN(_04719_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05841_ (.A1(_04565_),
    .A2(_04702_),
    .B(_04719_),
    .ZN(_00930_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05842_ (.A1(net88),
    .A2(net41),
    .ZN(_04720_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05843_ (.I(_04720_),
    .Z(_04721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05844_ (.I(_04720_),
    .Z(_04722_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05845_ (.A1(_04722_),
    .A2(\mem[60][0] ),
    .ZN(_04723_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05846_ (.A1(_04567_),
    .A2(_04721_),
    .B(_04723_),
    .ZN(_00931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05847_ (.A1(_04722_),
    .A2(\mem[60][1] ),
    .ZN(_04724_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05848_ (.A1(_04572_),
    .A2(_04721_),
    .B(_04724_),
    .ZN(_00932_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05849_ (.A1(_04722_),
    .A2(\mem[60][2] ),
    .ZN(_04725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05850_ (.A1(_04574_),
    .A2(_04721_),
    .B(_04725_),
    .ZN(_00933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05851_ (.A1(_04722_),
    .A2(\mem[60][3] ),
    .ZN(_04726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05852_ (.A1(_04576_),
    .A2(_04721_),
    .B(_04726_),
    .ZN(_00934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05853_ (.I(_04720_),
    .Z(_04727_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05854_ (.A1(_04727_),
    .A2(\mem[60][4] ),
    .ZN(_04728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05855_ (.A1(_04578_),
    .A2(_04721_),
    .B(_04728_),
    .ZN(_00935_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05856_ (.A1(_04727_),
    .A2(\mem[60][5] ),
    .ZN(_04729_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05857_ (.A1(_04581_),
    .A2(_04721_),
    .B(_04729_),
    .ZN(_00936_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05858_ (.A1(_04727_),
    .A2(\mem[60][6] ),
    .ZN(_04730_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05859_ (.A1(_04583_),
    .A2(_04721_),
    .B(_04730_),
    .ZN(_00937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05860_ (.A1(_04727_),
    .A2(\mem[60][7] ),
    .ZN(_04731_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05861_ (.A1(_04585_),
    .A2(_04721_),
    .B(_04731_),
    .ZN(_00938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05862_ (.A1(_04727_),
    .A2(\mem[60][8] ),
    .ZN(_04732_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05863_ (.A1(_04587_),
    .A2(_04721_),
    .B(_04732_),
    .ZN(_00939_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05864_ (.A1(_04727_),
    .A2(\mem[60][9] ),
    .ZN(_04733_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05865_ (.A1(_04589_),
    .A2(_04721_),
    .B(_04733_),
    .ZN(_00940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05866_ (.A1(_04727_),
    .A2(\mem[60][10] ),
    .ZN(_04734_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05867_ (.A1(_04591_),
    .A2(_04722_),
    .B(_04734_),
    .ZN(_00941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05868_ (.A1(_04727_),
    .A2(\mem[60][11] ),
    .ZN(_04735_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05869_ (.A1(_04593_),
    .A2(_04722_),
    .B(_04735_),
    .ZN(_00942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05870_ (.A1(_04727_),
    .A2(\mem[60][12] ),
    .ZN(_04736_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05871_ (.A1(_04595_),
    .A2(_04722_),
    .B(_04736_),
    .ZN(_00943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05872_ (.A1(_04727_),
    .A2(\mem[60][13] ),
    .ZN(_04737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05873_ (.A1(_04561_),
    .A2(_04722_),
    .B(_04737_),
    .ZN(_00944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05874_ (.A1(_04720_),
    .A2(\mem[60][14] ),
    .ZN(_04738_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05875_ (.A1(_04563_),
    .A2(_04722_),
    .B(_04738_),
    .ZN(_00945_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05876_ (.A1(_04720_),
    .A2(\mem[60][15] ),
    .ZN(_04739_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05877_ (.A1(_04565_),
    .A2(_04722_),
    .B(_04739_),
    .ZN(_00946_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05878_ (.A1(net88),
    .A2(_03566_),
    .ZN(_04740_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05879_ (.I(_04740_),
    .Z(_04741_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05880_ (.I(_04740_),
    .Z(_04742_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05881_ (.A1(_04742_),
    .A2(\mem[61][0] ),
    .ZN(_04743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05882_ (.A1(_04567_),
    .A2(_04741_),
    .B(_04743_),
    .ZN(_00947_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05883_ (.A1(_04742_),
    .A2(\mem[61][1] ),
    .ZN(_04744_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05884_ (.A1(_04572_),
    .A2(_04741_),
    .B(_04744_),
    .ZN(_00948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05885_ (.A1(_04742_),
    .A2(\mem[61][2] ),
    .ZN(_04745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05886_ (.A1(_04574_),
    .A2(_04741_),
    .B(_04745_),
    .ZN(_00949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05887_ (.A1(_04742_),
    .A2(\mem[61][3] ),
    .ZN(_04746_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05888_ (.A1(_04576_),
    .A2(_04741_),
    .B(_04746_),
    .ZN(_00950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05889_ (.I(_04740_),
    .Z(_04747_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05890_ (.A1(_04747_),
    .A2(\mem[61][4] ),
    .ZN(_04748_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05891_ (.A1(_04578_),
    .A2(_04741_),
    .B(_04748_),
    .ZN(_00951_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05892_ (.A1(_04747_),
    .A2(\mem[61][5] ),
    .ZN(_04749_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05893_ (.A1(_04581_),
    .A2(_04741_),
    .B(_04749_),
    .ZN(_00952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05894_ (.A1(_04747_),
    .A2(\mem[61][6] ),
    .ZN(_04750_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05895_ (.A1(_04583_),
    .A2(_04741_),
    .B(_04750_),
    .ZN(_00953_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05896_ (.A1(_04747_),
    .A2(\mem[61][7] ),
    .ZN(_04751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05897_ (.A1(_04585_),
    .A2(_04741_),
    .B(_04751_),
    .ZN(_00954_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05898_ (.A1(_04747_),
    .A2(\mem[61][8] ),
    .ZN(_04752_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05899_ (.A1(_04587_),
    .A2(_04741_),
    .B(_04752_),
    .ZN(_00955_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05900_ (.A1(_04747_),
    .A2(\mem[61][9] ),
    .ZN(_04753_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05901_ (.A1(_04589_),
    .A2(_04741_),
    .B(_04753_),
    .ZN(_00956_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05902_ (.A1(_04747_),
    .A2(\mem[61][10] ),
    .ZN(_04754_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05903_ (.A1(_04591_),
    .A2(_04742_),
    .B(_04754_),
    .ZN(_00957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05904_ (.A1(_04747_),
    .A2(\mem[61][11] ),
    .ZN(_04755_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05905_ (.A1(_04593_),
    .A2(_04742_),
    .B(_04755_),
    .ZN(_00958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05906_ (.A1(_04747_),
    .A2(\mem[61][12] ),
    .ZN(_04756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05907_ (.A1(_04595_),
    .A2(_04742_),
    .B(_04756_),
    .ZN(_00959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05908_ (.A1(_04747_),
    .A2(\mem[61][13] ),
    .ZN(_04757_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05909_ (.A1(_04561_),
    .A2(_04742_),
    .B(_04757_),
    .ZN(_00960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05910_ (.A1(_04740_),
    .A2(\mem[61][14] ),
    .ZN(_04758_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05911_ (.A1(_04563_),
    .A2(_04742_),
    .B(_04758_),
    .ZN(_00961_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05912_ (.A1(_04740_),
    .A2(\mem[61][15] ),
    .ZN(_04759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05913_ (.A1(_04565_),
    .A2(_04742_),
    .B(_04759_),
    .ZN(_00962_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05914_ (.A1(net88),
    .A2(_01162_),
    .ZN(_04760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05915_ (.I(net89),
    .Z(_04761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05916_ (.I(net89),
    .Z(_04762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05917_ (.A1(_04762_),
    .A2(\mem[62][0] ),
    .ZN(_04763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05918_ (.A1(_04567_),
    .A2(_04761_),
    .B(_04763_),
    .ZN(_00963_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05919_ (.A1(_04762_),
    .A2(\mem[62][1] ),
    .ZN(_04764_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05920_ (.A1(_04572_),
    .A2(_04761_),
    .B(_04764_),
    .ZN(_00964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05921_ (.A1(_04762_),
    .A2(\mem[62][2] ),
    .ZN(_04765_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05922_ (.A1(_04574_),
    .A2(_04761_),
    .B(_04765_),
    .ZN(_00965_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05923_ (.A1(_04762_),
    .A2(\mem[62][3] ),
    .ZN(_04766_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05924_ (.A1(_04576_),
    .A2(_04761_),
    .B(_04766_),
    .ZN(_00966_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05925_ (.I(net89),
    .Z(_04767_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05926_ (.A1(_04767_),
    .A2(\mem[62][4] ),
    .ZN(_04768_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05927_ (.A1(_04578_),
    .A2(_04761_),
    .B(_04768_),
    .ZN(_00967_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05928_ (.A1(_04767_),
    .A2(\mem[62][5] ),
    .ZN(_04769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05929_ (.A1(_04581_),
    .A2(_04761_),
    .B(_04769_),
    .ZN(_00968_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05930_ (.A1(_04767_),
    .A2(\mem[62][6] ),
    .ZN(_04770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05931_ (.A1(_04583_),
    .A2(_04761_),
    .B(_04770_),
    .ZN(_00969_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05932_ (.A1(_04767_),
    .A2(\mem[62][7] ),
    .ZN(_04771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05933_ (.A1(_04585_),
    .A2(_04761_),
    .B(_04771_),
    .ZN(_00970_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05934_ (.A1(_04767_),
    .A2(\mem[62][8] ),
    .ZN(_04772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05935_ (.A1(_04587_),
    .A2(_04761_),
    .B(_04772_),
    .ZN(_00971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05936_ (.A1(_04767_),
    .A2(\mem[62][9] ),
    .ZN(_04773_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05937_ (.A1(_04589_),
    .A2(_04761_),
    .B(_04773_),
    .ZN(_00972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05938_ (.A1(_04767_),
    .A2(\mem[62][10] ),
    .ZN(_04774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05939_ (.A1(_04591_),
    .A2(_04762_),
    .B(_04774_),
    .ZN(_00973_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05940_ (.A1(_04767_),
    .A2(\mem[62][11] ),
    .ZN(_04775_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05941_ (.A1(_04593_),
    .A2(_04762_),
    .B(_04775_),
    .ZN(_00974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05942_ (.A1(_04767_),
    .A2(\mem[62][12] ),
    .ZN(_04776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05943_ (.A1(_04595_),
    .A2(_04762_),
    .B(_04776_),
    .ZN(_00975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05944_ (.A1(_04767_),
    .A2(\mem[62][13] ),
    .ZN(_04777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05945_ (.A1(_03438_),
    .A2(_04762_),
    .B(_04777_),
    .ZN(_00976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05946_ (.A1(net89),
    .A2(\mem[62][14] ),
    .ZN(_04778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05947_ (.A1(_03446_),
    .A2(_04762_),
    .B(_04778_),
    .ZN(_00977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05948_ (.A1(net89),
    .A2(\mem[62][15] ),
    .ZN(_04779_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05949_ (.A1(_03449_),
    .A2(_04762_),
    .B(_04779_),
    .ZN(_00978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05950_ (.A1(net93),
    .A2(_01431_),
    .ZN(_04780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05951_ (.I(_04780_),
    .Z(_04781_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05952_ (.I(_04780_),
    .Z(_04782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05953_ (.A1(_04782_),
    .A2(\mem[9][0] ),
    .ZN(_04783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05954_ (.A1(_03452_),
    .A2(_04781_),
    .B(_04783_),
    .ZN(_00979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05955_ (.A1(_04782_),
    .A2(\mem[9][1] ),
    .ZN(_04784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05956_ (.A1(_03461_),
    .A2(_04781_),
    .B(_04784_),
    .ZN(_00980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05957_ (.A1(_04782_),
    .A2(\mem[9][2] ),
    .ZN(_04785_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05958_ (.A1(_03464_),
    .A2(_04781_),
    .B(_04785_),
    .ZN(_00981_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05959_ (.A1(_04782_),
    .A2(\mem[9][3] ),
    .ZN(_04786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05960_ (.A1(_03467_),
    .A2(_04781_),
    .B(_04786_),
    .ZN(_00982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05961_ (.I(_04780_),
    .Z(_04787_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05962_ (.A1(_04787_),
    .A2(\mem[9][4] ),
    .ZN(_04788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05963_ (.A1(_03470_),
    .A2(_04781_),
    .B(_04788_),
    .ZN(_00983_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05964_ (.A1(_04787_),
    .A2(\mem[9][5] ),
    .ZN(_04789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05965_ (.A1(_03474_),
    .A2(_04781_),
    .B(_04789_),
    .ZN(_00984_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05966_ (.A1(_04787_),
    .A2(\mem[9][6] ),
    .ZN(_04790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05967_ (.A1(_03477_),
    .A2(_04781_),
    .B(_04790_),
    .ZN(_00985_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05968_ (.A1(_04787_),
    .A2(\mem[9][7] ),
    .ZN(_04791_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05969_ (.A1(_03480_),
    .A2(_04781_),
    .B(_04791_),
    .ZN(_00986_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05970_ (.A1(_04787_),
    .A2(\mem[9][8] ),
    .ZN(_04792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05971_ (.A1(_03483_),
    .A2(_04781_),
    .B(_04792_),
    .ZN(_00987_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05972_ (.A1(_04787_),
    .A2(\mem[9][9] ),
    .ZN(_04793_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05973_ (.A1(_03486_),
    .A2(_04781_),
    .B(_04793_),
    .ZN(_00988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05974_ (.A1(_04787_),
    .A2(\mem[9][10] ),
    .ZN(_04794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05975_ (.A1(_03489_),
    .A2(_04782_),
    .B(_04794_),
    .ZN(_00989_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05976_ (.A1(_04787_),
    .A2(\mem[9][11] ),
    .ZN(_04795_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05977_ (.A1(_03492_),
    .A2(_04782_),
    .B(_04795_),
    .ZN(_00990_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05978_ (.A1(_04787_),
    .A2(\mem[9][12] ),
    .ZN(_04796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05979_ (.A1(_03495_),
    .A2(_04782_),
    .B(_04796_),
    .ZN(_00991_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05980_ (.A1(_04787_),
    .A2(\mem[9][13] ),
    .ZN(_04797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05981_ (.A1(_03438_),
    .A2(_04782_),
    .B(_04797_),
    .ZN(_00992_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05982_ (.A1(_04780_),
    .A2(\mem[9][14] ),
    .ZN(_04798_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05983_ (.A1(_03446_),
    .A2(_04782_),
    .B(_04798_),
    .ZN(_00993_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05984_ (.A1(_04780_),
    .A2(\mem[9][15] ),
    .ZN(_04799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05985_ (.A1(_03449_),
    .A2(_04782_),
    .B(_04799_),
    .ZN(_00994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05986_ (.A1(_03790_),
    .A2(net70),
    .ZN(_04800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05987_ (.I(net71),
    .Z(_04801_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05988_ (.I(net71),
    .Z(_04802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05989_ (.A1(_04802_),
    .A2(\mem[49][0] ),
    .ZN(_04803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05990_ (.A1(_03452_),
    .A2(net72),
    .B(_04803_),
    .ZN(_00995_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05991_ (.A1(_04802_),
    .A2(\mem[49][1] ),
    .ZN(_04804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05992_ (.A1(_03461_),
    .A2(net72),
    .B(_04804_),
    .ZN(_00996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05993_ (.A1(_04802_),
    .A2(\mem[49][2] ),
    .ZN(_04805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05994_ (.A1(_03464_),
    .A2(net72),
    .B(_04805_),
    .ZN(_00997_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05995_ (.A1(_04802_),
    .A2(\mem[49][3] ),
    .ZN(_04806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05996_ (.A1(_03467_),
    .A2(net72),
    .B(_04806_),
    .ZN(_00998_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05997_ (.I(net71),
    .Z(_04807_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05998_ (.A1(_04807_),
    .A2(\mem[49][4] ),
    .ZN(_04808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05999_ (.A1(_03470_),
    .A2(net72),
    .B(_04808_),
    .ZN(_00999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06000_ (.A1(_04807_),
    .A2(\mem[49][5] ),
    .ZN(_04809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06001_ (.A1(_03474_),
    .A2(net72),
    .B(_04809_),
    .ZN(_01000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06002_ (.A1(_04807_),
    .A2(\mem[49][6] ),
    .ZN(_04810_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06003_ (.A1(_03477_),
    .A2(net72),
    .B(_04810_),
    .ZN(_01001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06004_ (.A1(_04807_),
    .A2(\mem[49][7] ),
    .ZN(_04811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06005_ (.A1(_03480_),
    .A2(net72),
    .B(_04811_),
    .ZN(_01002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06006_ (.A1(_04807_),
    .A2(\mem[49][8] ),
    .ZN(_04812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06007_ (.A1(_03483_),
    .A2(net72),
    .B(_04812_),
    .ZN(_01003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06008_ (.A1(_04807_),
    .A2(\mem[49][9] ),
    .ZN(_04813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06009_ (.A1(_03486_),
    .A2(net72),
    .B(_04813_),
    .ZN(_01004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06010_ (.A1(_04807_),
    .A2(\mem[49][10] ),
    .ZN(_04814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06011_ (.A1(_03489_),
    .A2(_04802_),
    .B(_04814_),
    .ZN(_01005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06012_ (.A1(_04807_),
    .A2(\mem[49][11] ),
    .ZN(_04815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06013_ (.A1(_03492_),
    .A2(_04802_),
    .B(_04815_),
    .ZN(_01006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06014_ (.A1(_04807_),
    .A2(\mem[49][12] ),
    .ZN(_04816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06015_ (.A1(_03495_),
    .A2(_04802_),
    .B(_04816_),
    .ZN(_01007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06016_ (.A1(_04807_),
    .A2(\mem[49][13] ),
    .ZN(_04817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06017_ (.A1(_03438_),
    .A2(_04802_),
    .B(_04817_),
    .ZN(_01008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06018_ (.A1(net71),
    .A2(\mem[49][14] ),
    .ZN(_04818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06019_ (.A1(_03446_),
    .A2(_04802_),
    .B(_04818_),
    .ZN(_01009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06020_ (.A1(net71),
    .A2(\mem[49][15] ),
    .ZN(_04819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06021_ (.A1(_03449_),
    .A2(_04802_),
    .B(_04819_),
    .ZN(_01010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06022_ (.A1(net60),
    .A2(net76),
    .ZN(_04820_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06023_ (.I(net77),
    .Z(_04821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06024_ (.I(net77),
    .Z(_04822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06025_ (.A1(_04822_),
    .A2(\mem[39][0] ),
    .ZN(_04823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06026_ (.A1(_03452_),
    .A2(_04821_),
    .B(_04823_),
    .ZN(_01011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06027_ (.A1(_04822_),
    .A2(\mem[39][1] ),
    .ZN(_04824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06028_ (.A1(_03461_),
    .A2(_04821_),
    .B(_04824_),
    .ZN(_01012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06029_ (.A1(_04822_),
    .A2(\mem[39][2] ),
    .ZN(_04825_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06030_ (.A1(_03464_),
    .A2(_04821_),
    .B(_04825_),
    .ZN(_01013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06031_ (.A1(_04822_),
    .A2(\mem[39][3] ),
    .ZN(_04826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06032_ (.A1(_03467_),
    .A2(_04821_),
    .B(_04826_),
    .ZN(_01014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06033_ (.I(_04820_),
    .Z(_04827_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06034_ (.A1(_04827_),
    .A2(\mem[39][4] ),
    .ZN(_04828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06035_ (.A1(_03470_),
    .A2(_04821_),
    .B(_04828_),
    .ZN(_01015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06036_ (.A1(_04827_),
    .A2(\mem[39][5] ),
    .ZN(_04829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06037_ (.A1(_03474_),
    .A2(_04821_),
    .B(_04829_),
    .ZN(_01016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06038_ (.A1(_04827_),
    .A2(\mem[39][6] ),
    .ZN(_04830_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06039_ (.A1(_03477_),
    .A2(_04821_),
    .B(_04830_),
    .ZN(_01017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06040_ (.A1(_04827_),
    .A2(\mem[39][7] ),
    .ZN(_04831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06041_ (.A1(_03480_),
    .A2(_04821_),
    .B(_04831_),
    .ZN(_01018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06042_ (.A1(_04827_),
    .A2(\mem[39][8] ),
    .ZN(_04832_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06043_ (.A1(_03483_),
    .A2(_04821_),
    .B(_04832_),
    .ZN(_01019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06044_ (.A1(_04827_),
    .A2(\mem[39][9] ),
    .ZN(_04833_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06045_ (.A1(_03486_),
    .A2(_04821_),
    .B(_04833_),
    .ZN(_01020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06046_ (.A1(_04827_),
    .A2(\mem[39][10] ),
    .ZN(_04834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06047_ (.A1(_03489_),
    .A2(_04822_),
    .B(_04834_),
    .ZN(_01021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06048_ (.A1(_04827_),
    .A2(\mem[39][11] ),
    .ZN(_04835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06049_ (.A1(_03492_),
    .A2(_04822_),
    .B(_04835_),
    .ZN(_01022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06050_ (.A1(_04827_),
    .A2(\mem[39][12] ),
    .ZN(_04836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06051_ (.A1(_03495_),
    .A2(_04822_),
    .B(_04836_),
    .ZN(_01023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06052_ (.A1(_04827_),
    .A2(\mem[39][13] ),
    .ZN(_04837_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06053_ (.A1(_03438_),
    .A2(_04822_),
    .B(_04837_),
    .ZN(_01024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06054_ (.A1(net77),
    .A2(\mem[39][14] ),
    .ZN(_04838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06055_ (.A1(_03446_),
    .A2(_04822_),
    .B(_04838_),
    .ZN(_01025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06056_ (.A1(_04820_),
    .A2(\mem[39][15] ),
    .ZN(_04839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06057_ (.A1(_03449_),
    .A2(_04822_),
    .B(_04839_),
    .ZN(_01026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06058_ (.A1(_03444_),
    .A2(\mem[7][0] ),
    .ZN(_04840_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06059_ (.A1(_03452_),
    .A2(net62),
    .B(_04840_),
    .ZN(_01027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06060_ (.I(net61),
    .Z(_04841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06061_ (.A1(_04841_),
    .A2(\mem[7][1] ),
    .ZN(_04842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06062_ (.A1(_03461_),
    .A2(net62),
    .B(_04842_),
    .ZN(_01028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06063_ (.A1(_04841_),
    .A2(\mem[7][2] ),
    .ZN(_04843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06064_ (.A1(_03464_),
    .A2(net62),
    .B(_04843_),
    .ZN(_01029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06065_ (.A1(_04841_),
    .A2(\mem[7][3] ),
    .ZN(_04844_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06066_ (.A1(_03467_),
    .A2(net62),
    .B(_04844_),
    .ZN(_01030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06067_ (.A1(_04841_),
    .A2(\mem[7][4] ),
    .ZN(_04845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06068_ (.A1(_03470_),
    .A2(net62),
    .B(_04845_),
    .ZN(_01031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06069_ (.A1(_04841_),
    .A2(\mem[7][5] ),
    .ZN(_04846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06070_ (.A1(_03474_),
    .A2(_03443_),
    .B(_04846_),
    .ZN(_01032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06071_ (.A1(_04841_),
    .A2(\mem[7][6] ),
    .ZN(_04847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06072_ (.A1(_03477_),
    .A2(net62),
    .B(_04847_),
    .ZN(_01033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06073_ (.A1(_04841_),
    .A2(\mem[7][7] ),
    .ZN(_04848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06074_ (.A1(_03480_),
    .A2(_03444_),
    .B(_04848_),
    .ZN(_01034_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06075_ (.A1(_04841_),
    .A2(\mem[7][8] ),
    .ZN(_04849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06076_ (.A1(_03483_),
    .A2(_03444_),
    .B(_04849_),
    .ZN(_01035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06077_ (.A1(_04841_),
    .A2(\mem[7][9] ),
    .ZN(_04850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06078_ (.A1(_03486_),
    .A2(_03444_),
    .B(_04850_),
    .ZN(_01036_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06079_ (.A1(_04841_),
    .A2(\mem[7][10] ),
    .ZN(_04851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06080_ (.A1(_03489_),
    .A2(_03444_),
    .B(_04851_),
    .ZN(_01037_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06081_ (.A1(net61),
    .A2(\mem[7][11] ),
    .ZN(_04852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06082_ (.A1(_03492_),
    .A2(_03444_),
    .B(_04852_),
    .ZN(_01038_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06083_ (.A1(net61),
    .A2(\mem[7][12] ),
    .ZN(_04853_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06084_ (.A1(_03495_),
    .A2(_03444_),
    .B(_04853_),
    .ZN(_01039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _06085_ (.I(net97),
    .ZN(_01040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06086_ (.I(_01040_),
    .Z(_01041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06087_ (.A1(_01041_),
    .A2(\mem[16][0] ),
    .ZN(_01042_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06088_ (.I(net131),
    .Z(_01043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06089_ (.I(_01043_),
    .Z(_01044_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06090_ (.A1(_01044_),
    .A2(\mem[17][0] ),
    .ZN(_01045_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06091_ (.A1(_01042_),
    .A2(_01045_),
    .ZN(_01046_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06092_ (.I(net3),
    .Z(_01047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06093_ (.A1(net58),
    .A2(_01047_),
    .ZN(_01048_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06094_ (.I(_01048_),
    .Z(_01049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06095_ (.I(_01049_),
    .Z(_01050_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06096_ (.A1(_01046_),
    .A2(_01050_),
    .ZN(_01051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06097_ (.A1(_01041_),
    .A2(\mem[18][0] ),
    .ZN(_01052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06098_ (.A1(_01044_),
    .A2(\mem[19][0] ),
    .ZN(_01053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06099_ (.A1(_01052_),
    .A2(_01053_),
    .ZN(_01054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06100_ (.I(net58),
    .ZN(_01055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06101_ (.A1(_01055_),
    .A2(net3),
    .ZN(_01056_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06102_ (.I(_01056_),
    .Z(_01057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06103_ (.I(_01057_),
    .Z(_01058_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06104_ (.A1(_01054_),
    .A2(_01058_),
    .ZN(_01059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06105_ (.A1(_01051_),
    .A2(_01059_),
    .ZN(_01060_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06106_ (.A1(_01041_),
    .A2(\mem[20][0] ),
    .ZN(_01061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06107_ (.I(_01043_),
    .Z(_01062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06108_ (.A1(_01062_),
    .A2(\mem[21][0] ),
    .ZN(_01063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06109_ (.A1(_01061_),
    .A2(_01063_),
    .ZN(_01064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06110_ (.I(net3),
    .ZN(_01065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06111_ (.A1(_01065_),
    .A2(net58),
    .ZN(_01066_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06112_ (.I(_01066_),
    .Z(_01067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06113_ (.I(_01067_),
    .Z(_01068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06114_ (.A1(_01064_),
    .A2(_01068_),
    .ZN(_01069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06115_ (.I(_01040_),
    .Z(_01070_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06116_ (.A1(_01070_),
    .A2(\mem[22][0] ),
    .ZN(_01071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06117_ (.A1(_01062_),
    .A2(\mem[23][0] ),
    .ZN(_01072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06118_ (.A1(_01071_),
    .A2(_01072_),
    .ZN(_01073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06119_ (.A1(net58),
    .A2(net3),
    .ZN(_01074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06120_ (.I(net59),
    .ZN(_01075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06121_ (.A1(_01073_),
    .A2(_01075_),
    .ZN(_01076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06122_ (.A1(_01069_),
    .A2(_01076_),
    .ZN(_01077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06123_ (.I(net4),
    .ZN(_01078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06124_ (.I(net86),
    .ZN(_01079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06125_ (.A1(_01078_),
    .A2(_01079_),
    .A3(net136),
    .ZN(_01080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06126_ (.I(net137),
    .ZN(_01081_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06127_ (.I(_01081_),
    .Z(_01082_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06128_ (.A1(_01060_),
    .A2(_01077_),
    .B(_01082_),
    .ZN(_01083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06129_ (.A1(_01041_),
    .A2(\mem[24][0] ),
    .ZN(_01084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06130_ (.A1(_01044_),
    .A2(\mem[25][0] ),
    .ZN(_01085_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06131_ (.A1(_01084_),
    .A2(_01085_),
    .ZN(_01086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06132_ (.A1(_01086_),
    .A2(_01050_),
    .ZN(_01087_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06133_ (.A1(_01041_),
    .A2(\mem[26][0] ),
    .ZN(_01088_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06134_ (.A1(_01062_),
    .A2(\mem[27][0] ),
    .ZN(_01089_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06135_ (.A1(_01088_),
    .A2(_01089_),
    .ZN(_01090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06136_ (.A1(_01090_),
    .A2(_01058_),
    .ZN(_01091_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06137_ (.A1(_01087_),
    .A2(_01091_),
    .ZN(_01092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06138_ (.A1(_01070_),
    .A2(\mem[28][0] ),
    .ZN(_01093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06139_ (.A1(_01062_),
    .A2(\mem[29][0] ),
    .ZN(_01094_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06140_ (.A1(_01093_),
    .A2(_01094_),
    .ZN(_01095_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06141_ (.A1(_01095_),
    .A2(_01068_),
    .ZN(_01096_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06142_ (.A1(_01070_),
    .A2(\mem[30][0] ),
    .ZN(_01097_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06143_ (.A1(_01062_),
    .A2(\mem[31][0] ),
    .ZN(_01098_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06144_ (.A1(_01097_),
    .A2(_01098_),
    .ZN(_01099_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06145_ (.A1(_01099_),
    .A2(_01075_),
    .ZN(_01100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06146_ (.A1(_01096_),
    .A2(_01100_),
    .ZN(_01101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06147_ (.A1(_01079_),
    .A2(net4),
    .A3(net68),
    .ZN(_01102_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06148_ (.I(net118),
    .ZN(_01103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06149_ (.I(_01103_),
    .Z(_01104_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06150_ (.A1(_01092_),
    .A2(_01101_),
    .B(_01104_),
    .ZN(_01105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06151_ (.A1(_01083_),
    .A2(_01105_),
    .ZN(_01106_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06152_ (.A1(_01041_),
    .A2(\mem[32][0] ),
    .ZN(_01107_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06153_ (.A1(_01062_),
    .A2(\mem[33][0] ),
    .ZN(_01108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06154_ (.A1(_01107_),
    .A2(_01108_),
    .ZN(_01109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06155_ (.A1(_01109_),
    .A2(_01050_),
    .ZN(_01110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06156_ (.A1(_01070_),
    .A2(\mem[34][0] ),
    .ZN(_01111_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06157_ (.A1(_01062_),
    .A2(\mem[35][0] ),
    .ZN(_01112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06158_ (.A1(_01111_),
    .A2(_01112_),
    .ZN(_01113_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06159_ (.A1(_01113_),
    .A2(_01058_),
    .ZN(_01114_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06160_ (.A1(_01110_),
    .A2(_01114_),
    .ZN(_01115_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06161_ (.A1(_01070_),
    .A2(\mem[36][0] ),
    .ZN(_01116_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06162_ (.A1(_01062_),
    .A2(\mem[37][0] ),
    .ZN(_01117_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06163_ (.A1(_01116_),
    .A2(_01117_),
    .ZN(_01118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06164_ (.A1(_01118_),
    .A2(_01068_),
    .ZN(_01119_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06165_ (.A1(_01070_),
    .A2(\mem[38][0] ),
    .ZN(_01120_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06166_ (.I(net131),
    .Z(_01121_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06167_ (.A1(_01121_),
    .A2(\mem[39][0] ),
    .ZN(_01122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06168_ (.A1(_01120_),
    .A2(_01122_),
    .ZN(_01123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06169_ (.A1(_01123_),
    .A2(_01075_),
    .ZN(_01124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06170_ (.A1(_01119_),
    .A2(_01124_),
    .ZN(_01125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06171_ (.A1(_01079_),
    .A2(net4),
    .A3(net68),
    .ZN(_01126_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06172_ (.I(net76),
    .Z(_01127_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06173_ (.A1(_01115_),
    .A2(_01125_),
    .B(_01127_),
    .ZN(_01128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06174_ (.A1(_01070_),
    .A2(\mem[40][0] ),
    .ZN(_01129_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06175_ (.A1(_01062_),
    .A2(\mem[41][0] ),
    .ZN(_01130_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06176_ (.A1(_01129_),
    .A2(_01130_),
    .ZN(_01131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06177_ (.A1(_01131_),
    .A2(_01050_),
    .ZN(_01132_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06178_ (.A1(_01070_),
    .A2(\mem[42][0] ),
    .ZN(_01133_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06179_ (.A1(_01062_),
    .A2(\mem[43][0] ),
    .ZN(_01134_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06180_ (.A1(_01133_),
    .A2(_01134_),
    .ZN(_01135_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06181_ (.A1(_01135_),
    .A2(_01058_),
    .ZN(_01136_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06182_ (.A1(_01132_),
    .A2(_01136_),
    .ZN(_01137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06183_ (.A1(_01070_),
    .A2(\mem[44][0] ),
    .ZN(_01138_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06184_ (.A1(_01121_),
    .A2(\mem[45][0] ),
    .ZN(_01139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06185_ (.A1(_01138_),
    .A2(_01139_),
    .ZN(_01140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06186_ (.A1(_01140_),
    .A2(_01068_),
    .ZN(_01141_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06187_ (.A1(_01070_),
    .A2(\mem[46][0] ),
    .ZN(_01142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06188_ (.A1(_01121_),
    .A2(\mem[47][0] ),
    .ZN(_01143_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06189_ (.A1(_01142_),
    .A2(_01143_),
    .ZN(_01144_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06190_ (.A1(_01144_),
    .A2(_01075_),
    .ZN(_01145_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06191_ (.A1(_01141_),
    .A2(_01145_),
    .ZN(_01146_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06192_ (.A1(net142),
    .A2(_01079_),
    .A3(net136),
    .Z(_01147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06193_ (.I(_01147_),
    .ZN(_01148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06194_ (.I(_01148_),
    .Z(_01149_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06195_ (.A1(_01137_),
    .A2(_01146_),
    .B(_01149_),
    .ZN(_01150_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06196_ (.A1(_01128_),
    .A2(_01150_),
    .ZN(_01151_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06197_ (.A1(_01106_),
    .A2(_01151_),
    .ZN(_01152_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06198_ (.I(net58),
    .Z(_01153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06199_ (.A1(_01065_),
    .A2(net131),
    .A3(_01153_),
    .ZN(_01154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06200_ (.A1(net132),
    .A2(\mem[4][0] ),
    .ZN(_01155_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06201_ (.I(_01121_),
    .Z(_01156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06202_ (.A1(_01050_),
    .A2(\mem[1][0] ),
    .A3(_01156_),
    .ZN(_01157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06203_ (.A1(_01155_),
    .A2(_01157_),
    .ZN(_01158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06204_ (.A1(_01068_),
    .A2(_01156_),
    .A3(\mem[5][0] ),
    .ZN(_01159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06205_ (.A1(net59),
    .A2(net97),
    .ZN(_01160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06206_ (.I(net98),
    .Z(_01161_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06207_ (.I(_01161_),
    .Z(_01162_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06208_ (.A1(_01162_),
    .A2(\mem[6][0] ),
    .ZN(_01163_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06209_ (.A1(_01159_),
    .A2(_01163_),
    .ZN(_01164_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06210_ (.A1(_01158_),
    .A2(_01164_),
    .ZN(_01165_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06211_ (.I(_01040_),
    .Z(_01166_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06212_ (.I(_01166_),
    .Z(_01167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06213_ (.A1(_01058_),
    .A2(_01167_),
    .A3(\mem[2][0] ),
    .ZN(_01168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06214_ (.A1(_01058_),
    .A2(_01156_),
    .A3(\mem[3][0] ),
    .ZN(_01169_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06215_ (.A1(_01168_),
    .A2(_01169_),
    .ZN(_01170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06216_ (.A1(net59),
    .A2(_01040_),
    .ZN(_01171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06217_ (.I(_01171_),
    .Z(_01172_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06218_ (.I(_01172_),
    .Z(_01173_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06219_ (.A1(_01173_),
    .A2(\mem[7][0] ),
    .ZN(_01174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06220_ (.A1(_01050_),
    .A2(\mem[0][0] ),
    .A3(_01167_),
    .ZN(_01175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06221_ (.A1(_01174_),
    .A2(_01175_),
    .ZN(_01176_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06222_ (.A1(_01170_),
    .A2(_01176_),
    .ZN(_01177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06223_ (.A1(net136),
    .A2(net86),
    .ZN(_01178_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06224_ (.A1(net134),
    .A2(net142),
    .ZN(_01179_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06225_ (.A1(_01165_),
    .A2(_01177_),
    .B(_01179_),
    .ZN(_01180_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06226_ (.A1(net41),
    .A2(\mem[12][0] ),
    .ZN(_01181_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06227_ (.A1(_01068_),
    .A2(_01156_),
    .A3(\mem[13][0] ),
    .ZN(_01182_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06228_ (.A1(_01181_),
    .A2(_01182_),
    .ZN(_01183_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06229_ (.A1(_01162_),
    .A2(\mem[14][0] ),
    .ZN(_01184_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06230_ (.A1(_01173_),
    .A2(\mem[15][0] ),
    .ZN(_01185_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06231_ (.A1(_01184_),
    .A2(_01185_),
    .ZN(_01186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06232_ (.A1(_01183_),
    .A2(_01186_),
    .ZN(_01187_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06233_ (.A1(_01167_),
    .A2(\mem[8][0] ),
    .ZN(_01188_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06234_ (.A1(_01156_),
    .A2(\mem[9][0] ),
    .ZN(_01189_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06235_ (.I(_01153_),
    .Z(_01190_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06236_ (.A1(_01188_),
    .A2(_01189_),
    .B(_01190_),
    .ZN(_01191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06237_ (.A1(_01167_),
    .A2(\mem[10][0] ),
    .ZN(_01192_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06238_ (.A1(_01156_),
    .A2(\mem[11][0] ),
    .ZN(_01193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06239_ (.I(_01055_),
    .Z(_01194_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06240_ (.A1(_01192_),
    .A2(_01193_),
    .B(_01194_),
    .ZN(_01195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06241_ (.I(_01065_),
    .Z(_01196_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06242_ (.A1(_01191_),
    .A2(_01195_),
    .B(_01196_),
    .ZN(_01197_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06243_ (.A1(net134),
    .A2(net4),
    .ZN(_01198_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06244_ (.A1(_01187_),
    .A2(_01197_),
    .B(net110),
    .ZN(_01199_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06245_ (.A1(_01180_),
    .A2(_01199_),
    .ZN(_01200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06246_ (.A1(net41),
    .A2(\mem[52][0] ),
    .ZN(_01201_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06247_ (.A1(_01068_),
    .A2(_01156_),
    .A3(\mem[53][0] ),
    .ZN(_01202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06248_ (.A1(_01201_),
    .A2(_01202_),
    .ZN(_01203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06249_ (.A1(_01162_),
    .A2(\mem[54][0] ),
    .ZN(_01204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06250_ (.A1(_01173_),
    .A2(\mem[55][0] ),
    .ZN(_01205_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06251_ (.A1(_01204_),
    .A2(_01205_),
    .ZN(_01206_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06252_ (.A1(_01203_),
    .A2(_01206_),
    .ZN(_01207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06253_ (.A1(_01167_),
    .A2(\mem[48][0] ),
    .ZN(_01208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06254_ (.A1(_01156_),
    .A2(\mem[49][0] ),
    .ZN(_01209_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06255_ (.A1(_01208_),
    .A2(_01209_),
    .B(_01190_),
    .ZN(_01210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06256_ (.A1(_01167_),
    .A2(\mem[50][0] ),
    .ZN(_01211_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06257_ (.I(_01043_),
    .Z(_01212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06258_ (.I(_01212_),
    .Z(_01213_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06259_ (.A1(_01213_),
    .A2(\mem[51][0] ),
    .ZN(_01214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06260_ (.A1(_01211_),
    .A2(_01214_),
    .B(_01194_),
    .ZN(_01215_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06261_ (.A1(_01210_),
    .A2(_01215_),
    .B(_01196_),
    .ZN(_01216_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06262_ (.A1(_01078_),
    .A2(net68),
    .A3(net6),
    .ZN(_01217_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06263_ (.A1(_01207_),
    .A2(_01216_),
    .B(net69),
    .ZN(_01218_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06264_ (.A1(_01068_),
    .A2(_01167_),
    .A3(\mem[60][0] ),
    .ZN(_01219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06265_ (.A1(_01068_),
    .A2(_01156_),
    .A3(\mem[61][0] ),
    .ZN(_01220_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06266_ (.A1(_01219_),
    .A2(_01220_),
    .ZN(_01221_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06267_ (.A1(_01162_),
    .A2(\mem[62][0] ),
    .ZN(_01222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06268_ (.A1(_01173_),
    .A2(\mem[63][0] ),
    .ZN(_01223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06269_ (.A1(_01222_),
    .A2(_01223_),
    .ZN(_01224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06270_ (.A1(_01221_),
    .A2(_01224_),
    .ZN(_01225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06271_ (.A1(_01167_),
    .A2(\mem[56][0] ),
    .ZN(_01226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06272_ (.A1(_01156_),
    .A2(\mem[57][0] ),
    .ZN(_01227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06273_ (.A1(_01226_),
    .A2(_01227_),
    .B(_01190_),
    .ZN(_01228_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06274_ (.A1(_01167_),
    .A2(\mem[58][0] ),
    .ZN(_01229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06275_ (.A1(_01213_),
    .A2(\mem[59][0] ),
    .ZN(_01230_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06276_ (.A1(_01229_),
    .A2(_01230_),
    .B(_01194_),
    .ZN(_01231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06277_ (.A1(_01228_),
    .A2(_01231_),
    .B(_01196_),
    .ZN(_01232_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06278_ (.A1(net4),
    .A2(net68),
    .A3(net86),
    .ZN(_01233_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06279_ (.A1(_01225_),
    .A2(_01232_),
    .B(net87),
    .ZN(_01234_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06280_ (.A1(_01218_),
    .A2(_01234_),
    .ZN(_01235_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06281_ (.A1(_01152_),
    .A2(_01200_),
    .A3(_01235_),
    .ZN(_00000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06282_ (.A1(_01068_),
    .A2(_01167_),
    .A3(\mem[36][1] ),
    .ZN(_01236_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06283_ (.I(_01057_),
    .Z(_01237_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06284_ (.A1(_01237_),
    .A2(_01213_),
    .A3(\mem[35][1] ),
    .ZN(_01238_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06285_ (.A1(_01236_),
    .A2(_01238_),
    .ZN(_01239_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06286_ (.I(_01066_),
    .Z(_01240_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06287_ (.I(_01240_),
    .Z(_01241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06288_ (.I(_01121_),
    .Z(_01242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06289_ (.A1(_01241_),
    .A2(_01242_),
    .A3(\mem[37][1] ),
    .ZN(_01243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06290_ (.A1(_01162_),
    .A2(\mem[38][1] ),
    .ZN(_01244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06291_ (.A1(_01243_),
    .A2(_01244_),
    .ZN(_01245_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06292_ (.A1(_01239_),
    .A2(_01245_),
    .ZN(_01246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06293_ (.I(_01166_),
    .Z(_01247_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06294_ (.A1(_01058_),
    .A2(_01247_),
    .A3(\mem[34][1] ),
    .ZN(_01248_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06295_ (.I(_01121_),
    .Z(_01249_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06296_ (.A1(_01050_),
    .A2(_01249_),
    .A3(\mem[33][1] ),
    .ZN(_01250_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06297_ (.A1(_01248_),
    .A2(_01250_),
    .ZN(_01251_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06298_ (.A1(_01173_),
    .A2(\mem[39][1] ),
    .ZN(_01252_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06299_ (.I(_01048_),
    .Z(_01253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06300_ (.I(_01253_),
    .Z(_01254_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06301_ (.I(_01040_),
    .Z(_01255_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06302_ (.I(_01255_),
    .Z(_01256_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06303_ (.A1(_01254_),
    .A2(_01256_),
    .A3(\mem[32][1] ),
    .ZN(_01257_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06304_ (.A1(_01252_),
    .A2(_01257_),
    .ZN(_01258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06305_ (.A1(_01251_),
    .A2(_01258_),
    .ZN(_01259_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06306_ (.A1(_01246_),
    .A2(_01259_),
    .ZN(_01260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06307_ (.I(_01127_),
    .Z(_01261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06308_ (.A1(_01260_),
    .A2(_01261_),
    .ZN(_01262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06309_ (.I(_01067_),
    .Z(_01263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06310_ (.I(_01166_),
    .Z(_01264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06311_ (.A1(_01263_),
    .A2(_01264_),
    .A3(\mem[44][1] ),
    .ZN(_01265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06312_ (.I(net122),
    .Z(_01266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06313_ (.I(_01266_),
    .Z(_01267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06314_ (.I(_01267_),
    .Z(_01268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06315_ (.I(_01121_),
    .Z(_01269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06316_ (.A1(_01268_),
    .A2(_01269_),
    .A3(\mem[43][1] ),
    .ZN(_01270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06317_ (.A1(_01265_),
    .A2(_01270_),
    .ZN(_01271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06318_ (.I(_01240_),
    .Z(_01272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06319_ (.I(_01212_),
    .Z(_01273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06320_ (.A1(_01272_),
    .A2(_01273_),
    .A3(\mem[45][1] ),
    .ZN(_01274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06321_ (.I(_01161_),
    .Z(_01275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06322_ (.A1(_01275_),
    .A2(\mem[46][1] ),
    .ZN(_01276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06323_ (.A1(_01274_),
    .A2(_01276_),
    .ZN(_01277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06324_ (.A1(_01271_),
    .A2(_01277_),
    .ZN(_01278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06325_ (.I(_01057_),
    .Z(_01279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06326_ (.I(_01166_),
    .Z(_01280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06327_ (.A1(_01279_),
    .A2(_01280_),
    .A3(\mem[42][1] ),
    .ZN(_01281_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06328_ (.I(_01049_),
    .Z(_01282_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06329_ (.I(_01212_),
    .Z(_01283_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06330_ (.A1(_01282_),
    .A2(_01283_),
    .A3(\mem[41][1] ),
    .ZN(_01284_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06331_ (.A1(_01281_),
    .A2(_01284_),
    .ZN(_01285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06332_ (.I(_01171_),
    .Z(_01286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06333_ (.A1(_01286_),
    .A2(\mem[47][1] ),
    .ZN(_01287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06334_ (.I(_01253_),
    .Z(_01288_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06335_ (.I(_01255_),
    .Z(_01289_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06336_ (.A1(_01288_),
    .A2(_01289_),
    .A3(\mem[40][1] ),
    .ZN(_01290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06337_ (.A1(_01287_),
    .A2(_01290_),
    .ZN(_01291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06338_ (.A1(_01285_),
    .A2(_01291_),
    .ZN(_01292_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06339_ (.A1(_01278_),
    .A2(_01292_),
    .ZN(_01293_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06340_ (.I(_01149_),
    .Z(_01294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06341_ (.A1(_01293_),
    .A2(_01294_),
    .ZN(_01295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06342_ (.A1(_01262_),
    .A2(_01295_),
    .ZN(_01296_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06343_ (.I(_01067_),
    .Z(_01297_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06344_ (.I(_01166_),
    .Z(_01298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06345_ (.A1(_01297_),
    .A2(_01298_),
    .A3(\mem[52][1] ),
    .ZN(_01299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06346_ (.I(_01267_),
    .Z(_01300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06347_ (.I(_01212_),
    .Z(_01301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06348_ (.A1(_01300_),
    .A2(_01301_),
    .A3(\mem[51][1] ),
    .ZN(_01302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06349_ (.A1(_01299_),
    .A2(_01302_),
    .ZN(_01303_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06350_ (.I(_01240_),
    .Z(_01304_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06351_ (.I(_01043_),
    .Z(_01305_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06352_ (.I(_01305_),
    .Z(_01306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06353_ (.A1(_01304_),
    .A2(_01306_),
    .A3(\mem[53][1] ),
    .ZN(_01307_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06354_ (.I(_01161_),
    .Z(_01308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06355_ (.A1(_01308_),
    .A2(\mem[54][1] ),
    .ZN(_01309_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06356_ (.A1(_01307_),
    .A2(_01309_),
    .ZN(_01310_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06357_ (.A1(_01303_),
    .A2(_01310_),
    .ZN(_01311_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06358_ (.I(_01267_),
    .Z(_01312_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06359_ (.I(_01040_),
    .Z(_01313_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06360_ (.I(_01313_),
    .Z(_01314_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06361_ (.A1(_01312_),
    .A2(_01314_),
    .A3(\mem[50][1] ),
    .ZN(_01315_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06362_ (.I(_01253_),
    .Z(_01316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06363_ (.I(_01305_),
    .Z(_01317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06364_ (.A1(_01316_),
    .A2(_01317_),
    .A3(\mem[49][1] ),
    .ZN(_01318_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06365_ (.A1(_01315_),
    .A2(_01318_),
    .ZN(_01319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06366_ (.I(_01171_),
    .Z(_01320_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06367_ (.A1(_01320_),
    .A2(\mem[55][1] ),
    .ZN(_01321_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06368_ (.I(_01048_),
    .Z(_01322_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06369_ (.I(_01322_),
    .Z(_01323_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06370_ (.I(_01255_),
    .Z(_01324_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06371_ (.A1(_01323_),
    .A2(_01324_),
    .A3(\mem[48][1] ),
    .ZN(_01325_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06372_ (.A1(_01321_),
    .A2(_01325_),
    .ZN(_01326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06373_ (.A1(_01319_),
    .A2(_01326_),
    .ZN(_01327_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06374_ (.A1(_01311_),
    .A2(_01327_),
    .ZN(_01328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06375_ (.I(net69),
    .ZN(_01329_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06376_ (.I(net70),
    .Z(_01330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06377_ (.I(_01330_),
    .Z(_01331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06378_ (.A1(_01328_),
    .A2(_01331_),
    .ZN(_01332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06379_ (.I(_01240_),
    .Z(_01333_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06380_ (.I(_01313_),
    .Z(_01334_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06381_ (.A1(_01333_),
    .A2(_01334_),
    .A3(\mem[60][1] ),
    .ZN(_01335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06382_ (.I(_01266_),
    .Z(_01336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06383_ (.I(_01305_),
    .Z(_01337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06384_ (.A1(_01336_),
    .A2(_01337_),
    .A3(\mem[59][1] ),
    .ZN(_01338_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06385_ (.A1(_01335_),
    .A2(_01338_),
    .ZN(_01339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06386_ (.I(_01066_),
    .Z(_01340_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06387_ (.I(_01043_),
    .Z(_01341_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06388_ (.I(_01341_),
    .Z(_01342_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06389_ (.A1(_01340_),
    .A2(_01342_),
    .A3(\mem[61][1] ),
    .ZN(_01343_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06390_ (.I(net98),
    .Z(_01344_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06391_ (.A1(_01344_),
    .A2(\mem[62][1] ),
    .ZN(_01345_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06392_ (.A1(_01343_),
    .A2(_01345_),
    .ZN(_01346_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06393_ (.A1(_01339_),
    .A2(_01346_),
    .ZN(_01347_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06394_ (.I(_01266_),
    .Z(_01348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06395_ (.I(_01313_),
    .Z(_01349_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06396_ (.A1(_01348_),
    .A2(_01349_),
    .A3(\mem[58][1] ),
    .ZN(_01350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06397_ (.I(_01253_),
    .Z(_01351_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06398_ (.I(_01341_),
    .Z(_01352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06399_ (.A1(_01351_),
    .A2(_01352_),
    .A3(\mem[57][1] ),
    .ZN(_01353_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06400_ (.A1(_01350_),
    .A2(_01353_),
    .ZN(_01354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06401_ (.I(_01171_),
    .Z(_01355_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06402_ (.A1(_01355_),
    .A2(\mem[63][1] ),
    .ZN(_01356_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06403_ (.I(_01322_),
    .Z(_01357_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06404_ (.I(_01040_),
    .Z(_01358_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06405_ (.I(_01358_),
    .Z(_01359_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06406_ (.A1(_01357_),
    .A2(_01359_),
    .A3(\mem[56][1] ),
    .ZN(_01360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06407_ (.A1(_01356_),
    .A2(_01360_),
    .ZN(_01361_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06408_ (.A1(_01354_),
    .A2(_01361_),
    .ZN(_01362_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06409_ (.A1(_01347_),
    .A2(_01362_),
    .ZN(_01363_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06410_ (.I(net87),
    .ZN(_01364_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06411_ (.I(_01364_),
    .Z(_01365_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06412_ (.A1(_01363_),
    .A2(_01365_),
    .ZN(_01366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06413_ (.A1(_01332_),
    .A2(_01366_),
    .ZN(_01367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06414_ (.A1(_01296_),
    .A2(_01367_),
    .ZN(_01368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06415_ (.I(_01067_),
    .Z(_01369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06416_ (.I(_01166_),
    .Z(_01370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06417_ (.A1(_01369_),
    .A2(_01370_),
    .A3(\mem[4][1] ),
    .ZN(_01371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06418_ (.I(_01267_),
    .Z(_01372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06419_ (.I(_01212_),
    .Z(_01373_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06420_ (.A1(_01372_),
    .A2(_01373_),
    .A3(\mem[3][1] ),
    .ZN(_01374_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06421_ (.A1(_01371_),
    .A2(_01374_),
    .ZN(_01375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06422_ (.I(_01240_),
    .Z(_01376_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06423_ (.I(_01212_),
    .Z(_01377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06424_ (.A1(_01376_),
    .A2(_01377_),
    .A3(\mem[5][1] ),
    .ZN(_01378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06425_ (.I(_01161_),
    .Z(_01379_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06426_ (.A1(_01379_),
    .A2(\mem[6][1] ),
    .ZN(_01380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06427_ (.A1(_01378_),
    .A2(_01380_),
    .ZN(_01381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06428_ (.A1(_01375_),
    .A2(_01381_),
    .ZN(_01382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06429_ (.I(_01267_),
    .Z(_01383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06430_ (.I(_01166_),
    .Z(_01384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06431_ (.A1(_01383_),
    .A2(_01384_),
    .A3(\mem[2][1] ),
    .ZN(_01385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06432_ (.I(_01049_),
    .Z(_01386_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06433_ (.I(_01212_),
    .Z(_01387_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06434_ (.A1(_01386_),
    .A2(_01387_),
    .A3(\mem[1][1] ),
    .ZN(_01388_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06435_ (.A1(_01385_),
    .A2(_01388_),
    .ZN(_01389_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06436_ (.I(_01171_),
    .Z(_01390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06437_ (.A1(_01390_),
    .A2(\mem[7][1] ),
    .ZN(_01391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06438_ (.I(_01322_),
    .Z(_01392_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06439_ (.I(_01255_),
    .Z(_01393_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06440_ (.A1(_01392_),
    .A2(_01393_),
    .A3(\mem[0][1] ),
    .ZN(_01394_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06441_ (.A1(_01391_),
    .A2(_01394_),
    .ZN(_01395_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06442_ (.A1(_01389_),
    .A2(_01395_),
    .ZN(_01396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06443_ (.A1(_01382_),
    .A2(_01396_),
    .ZN(_01397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06444_ (.I(_01179_),
    .ZN(_01398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06445_ (.I(_01398_),
    .Z(_01399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06446_ (.A1(_01397_),
    .A2(_01399_),
    .ZN(_01400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06447_ (.I(_01240_),
    .Z(_01401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06448_ (.I(_01313_),
    .Z(_01402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06449_ (.A1(_01401_),
    .A2(_01402_),
    .A3(\mem[12][1] ),
    .ZN(_01403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06450_ (.I(_01266_),
    .Z(_01404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06451_ (.I(_01305_),
    .Z(_01405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06452_ (.A1(_01404_),
    .A2(_01405_),
    .A3(\mem[11][1] ),
    .ZN(_01406_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06453_ (.A1(_01403_),
    .A2(_01406_),
    .ZN(_01407_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06454_ (.I(_01066_),
    .Z(_01408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06455_ (.I(_01305_),
    .Z(_01409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06456_ (.A1(_01408_),
    .A2(_01409_),
    .A3(\mem[13][1] ),
    .ZN(_01410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06457_ (.I(net98),
    .Z(_01411_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06458_ (.A1(_01411_),
    .A2(\mem[14][1] ),
    .ZN(_01412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06459_ (.A1(_01410_),
    .A2(_01412_),
    .ZN(_01413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06460_ (.A1(_01407_),
    .A2(_01413_),
    .ZN(_01414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06461_ (.I(_01267_),
    .Z(_01415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06462_ (.I(_01313_),
    .Z(_01416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06463_ (.A1(_01415_),
    .A2(_01416_),
    .A3(\mem[10][1] ),
    .ZN(_01417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06464_ (.I(_01253_),
    .Z(_01418_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06465_ (.I(_01305_),
    .Z(_01419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06466_ (.A1(_01418_),
    .A2(_01419_),
    .A3(\mem[9][1] ),
    .ZN(_01420_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06467_ (.A1(_01417_),
    .A2(_01420_),
    .ZN(_01421_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06468_ (.I(_01171_),
    .Z(_01422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06469_ (.A1(_01422_),
    .A2(\mem[15][1] ),
    .ZN(_01423_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06470_ (.I(_01322_),
    .Z(_01424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06471_ (.I(_01358_),
    .Z(_01425_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06472_ (.A1(_01424_),
    .A2(_01425_),
    .A3(\mem[8][1] ),
    .ZN(_01426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06473_ (.A1(_01423_),
    .A2(_01426_),
    .ZN(_01427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06474_ (.A1(_01421_),
    .A2(_01427_),
    .ZN(_01428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06475_ (.A1(_01414_),
    .A2(_01428_),
    .ZN(_01429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06476_ (.I(net110),
    .ZN(_01430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06477_ (.I(_01430_),
    .Z(_01431_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06478_ (.I(_01431_),
    .Z(_01432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06479_ (.A1(_01429_),
    .A2(_01432_),
    .ZN(_01433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06480_ (.A1(_01400_),
    .A2(_01433_),
    .ZN(_01434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06481_ (.I(_01240_),
    .Z(_01435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06482_ (.I(_01313_),
    .Z(_01436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06483_ (.A1(_01435_),
    .A2(_01436_),
    .A3(\mem[20][1] ),
    .ZN(_01437_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06484_ (.I(_01266_),
    .Z(_01438_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06485_ (.I(_01305_),
    .Z(_01439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06486_ (.A1(_01438_),
    .A2(_01439_),
    .A3(\mem[19][1] ),
    .ZN(_01440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06487_ (.A1(_01437_),
    .A2(_01440_),
    .ZN(_01441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06488_ (.I(_01066_),
    .Z(_01442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06489_ (.I(_01341_),
    .Z(_01443_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06490_ (.A1(_01442_),
    .A2(_01443_),
    .A3(\mem[21][1] ),
    .ZN(_01444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06491_ (.I(net98),
    .Z(_01445_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06492_ (.A1(_01445_),
    .A2(\mem[22][1] ),
    .ZN(_01446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06493_ (.A1(_01444_),
    .A2(_01446_),
    .ZN(_01447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06494_ (.A1(_01441_),
    .A2(_01447_),
    .ZN(_01448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06495_ (.I(_01266_),
    .Z(_01449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06496_ (.I(_01255_),
    .Z(_01450_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06497_ (.A1(_01449_),
    .A2(_01450_),
    .A3(\mem[18][1] ),
    .ZN(_01451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06498_ (.I(_01253_),
    .Z(_01452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06499_ (.I(_01341_),
    .Z(_01453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06500_ (.A1(_01452_),
    .A2(_01453_),
    .A3(\mem[17][1] ),
    .ZN(_01454_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06501_ (.A1(_01451_),
    .A2(_01454_),
    .ZN(_01455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06502_ (.I(_01171_),
    .Z(_01456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06503_ (.A1(_01456_),
    .A2(\mem[23][1] ),
    .ZN(_01457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06504_ (.I(_01322_),
    .Z(_01458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06505_ (.I(_01358_),
    .Z(_01459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06506_ (.A1(_01458_),
    .A2(_01459_),
    .A3(\mem[16][1] ),
    .ZN(_01460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06507_ (.A1(_01457_),
    .A2(_01460_),
    .ZN(_01461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06508_ (.A1(_01455_),
    .A2(_01461_),
    .ZN(_01462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06509_ (.A1(_01448_),
    .A2(_01462_),
    .ZN(_01463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06510_ (.I(_01082_),
    .Z(_01464_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06511_ (.A1(_01463_),
    .A2(_01464_),
    .ZN(_01465_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06512_ (.I(_01066_),
    .Z(_01466_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06513_ (.I(_01255_),
    .Z(_01467_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06514_ (.A1(_01466_),
    .A2(_01467_),
    .A3(\mem[28][1] ),
    .ZN(_01468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06515_ (.I(_01043_),
    .Z(_01469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06516_ (.I(_01153_),
    .Z(_01470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06517_ (.A1(_01196_),
    .A2(_01469_),
    .A3(_01470_),
    .A4(\mem[27][1] ),
    .ZN(_01471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06518_ (.A1(_01468_),
    .A2(_01471_),
    .ZN(_01472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06519_ (.I(_01043_),
    .Z(_01473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06520_ (.I(_01047_),
    .Z(_01474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06521_ (.A1(_01194_),
    .A2(_01473_),
    .A3(_01474_),
    .A4(\mem[29][1] ),
    .ZN(_01475_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06522_ (.I(_01358_),
    .Z(_01476_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06523_ (.I(_01153_),
    .Z(_01477_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06524_ (.I(_01047_),
    .Z(_01478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06525_ (.A1(_01476_),
    .A2(_01477_),
    .A3(_01478_),
    .A4(\mem[30][1] ),
    .ZN(_01479_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06526_ (.A1(_01475_),
    .A2(_01479_),
    .ZN(_01480_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06527_ (.A1(_01472_),
    .A2(_01480_),
    .ZN(_01481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06528_ (.I(_01358_),
    .Z(_01482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06529_ (.I(_01065_),
    .Z(_01483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06530_ (.I(_01153_),
    .Z(_01484_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06531_ (.A1(_01482_),
    .A2(_01483_),
    .A3(_01484_),
    .A4(\mem[26][1] ),
    .ZN(_01485_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06532_ (.I(_01322_),
    .Z(_01486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06533_ (.I(_01341_),
    .Z(_01487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06534_ (.A1(_01486_),
    .A2(_01487_),
    .A3(\mem[25][1] ),
    .ZN(_01488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06535_ (.A1(_01485_),
    .A2(_01488_),
    .ZN(_01489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06536_ (.I(_01341_),
    .Z(_01490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06537_ (.I(_01047_),
    .Z(_01491_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06538_ (.A1(_01490_),
    .A2(_01190_),
    .A3(_01491_),
    .A4(\mem[31][1] ),
    .ZN(_01492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06539_ (.I(_01322_),
    .Z(_01493_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06540_ (.I(_01358_),
    .Z(_01494_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06541_ (.A1(_01493_),
    .A2(_01494_),
    .A3(\mem[24][1] ),
    .ZN(_01495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06542_ (.A1(_01492_),
    .A2(_01495_),
    .ZN(_01496_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06543_ (.A1(_01489_),
    .A2(_01496_),
    .ZN(_01497_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06544_ (.A1(_01481_),
    .A2(_01497_),
    .ZN(_01498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06545_ (.I(_01104_),
    .Z(_01499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06546_ (.A1(_01498_),
    .A2(_01499_),
    .ZN(_01500_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06547_ (.A1(_01465_),
    .A2(_01500_),
    .ZN(_01501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06548_ (.A1(_01434_),
    .A2(_01501_),
    .ZN(_01502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06549_ (.A1(_01368_),
    .A2(_01502_),
    .ZN(_00007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06550_ (.I(_01067_),
    .Z(_01503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06551_ (.I(_01166_),
    .Z(_01504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06552_ (.A1(_01503_),
    .A2(_01504_),
    .A3(\mem[36][2] ),
    .ZN(_01505_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06553_ (.A1(_01237_),
    .A2(_01213_),
    .A3(\mem[35][2] ),
    .ZN(_01506_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06554_ (.A1(_01505_),
    .A2(_01506_),
    .ZN(_01507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06555_ (.I(_01240_),
    .Z(_01508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06556_ (.A1(_01508_),
    .A2(_01242_),
    .A3(\mem[37][2] ),
    .ZN(_01509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06557_ (.I(_01161_),
    .Z(_01510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06558_ (.A1(_01510_),
    .A2(\mem[38][2] ),
    .ZN(_01511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06559_ (.A1(_01509_),
    .A2(_01511_),
    .ZN(_01512_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06560_ (.A1(_01507_),
    .A2(_01512_),
    .ZN(_01513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06561_ (.A1(_01058_),
    .A2(_01247_),
    .A3(\mem[34][2] ),
    .ZN(_01514_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06562_ (.A1(_01050_),
    .A2(_01249_),
    .A3(\mem[33][2] ),
    .ZN(_01515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06563_ (.A1(_01514_),
    .A2(_01515_),
    .ZN(_01516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06564_ (.A1(_01173_),
    .A2(\mem[39][2] ),
    .ZN(_01517_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06565_ (.A1(_01254_),
    .A2(_01256_),
    .A3(\mem[32][2] ),
    .ZN(_01518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06566_ (.A1(_01517_),
    .A2(_01518_),
    .ZN(_01519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06567_ (.A1(_01516_),
    .A2(_01519_),
    .ZN(_01520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06568_ (.A1(_01513_),
    .A2(_01520_),
    .ZN(_01521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06569_ (.A1(_01521_),
    .A2(_01261_),
    .ZN(_01522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06570_ (.I(_01166_),
    .Z(_01523_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06571_ (.A1(_01263_),
    .A2(_01523_),
    .A3(\mem[44][2] ),
    .ZN(_01524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06572_ (.A1(_01268_),
    .A2(_01269_),
    .A3(\mem[43][2] ),
    .ZN(_01525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06573_ (.A1(_01524_),
    .A2(_01525_),
    .ZN(_01526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06574_ (.A1(_01272_),
    .A2(_01273_),
    .A3(\mem[45][2] ),
    .ZN(_01527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06575_ (.A1(_01275_),
    .A2(\mem[46][2] ),
    .ZN(_01528_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06576_ (.A1(_01527_),
    .A2(_01528_),
    .ZN(_01529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06577_ (.A1(_01526_),
    .A2(_01529_),
    .ZN(_01530_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06578_ (.I(_01166_),
    .Z(_01531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06579_ (.A1(_01279_),
    .A2(_01531_),
    .A3(\mem[42][2] ),
    .ZN(_01532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06580_ (.A1(_01282_),
    .A2(_01283_),
    .A3(\mem[41][2] ),
    .ZN(_01533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06581_ (.A1(_01532_),
    .A2(_01533_),
    .ZN(_01534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06582_ (.I(_01171_),
    .Z(_01535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06583_ (.A1(_01535_),
    .A2(\mem[47][2] ),
    .ZN(_01536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06584_ (.I(_01255_),
    .Z(_01537_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06585_ (.A1(_01288_),
    .A2(_01537_),
    .A3(\mem[40][2] ),
    .ZN(_01538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06586_ (.A1(_01536_),
    .A2(_01538_),
    .ZN(_01539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06587_ (.A1(_01534_),
    .A2(_01539_),
    .ZN(_01540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06588_ (.A1(_01530_),
    .A2(_01540_),
    .ZN(_01541_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06589_ (.A1(_01541_),
    .A2(_01294_),
    .ZN(_01542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06590_ (.A1(_01522_),
    .A2(_01542_),
    .ZN(_01543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06591_ (.A1(_01297_),
    .A2(_01298_),
    .A3(\mem[52][2] ),
    .ZN(_01544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06592_ (.A1(_01300_),
    .A2(_01301_),
    .A3(\mem[51][2] ),
    .ZN(_01545_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06593_ (.A1(_01544_),
    .A2(_01545_),
    .ZN(_01546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06594_ (.I(_01066_),
    .Z(_01547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06595_ (.A1(_01547_),
    .A2(_01306_),
    .A3(\mem[53][2] ),
    .ZN(_01548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06596_ (.A1(_01308_),
    .A2(\mem[54][2] ),
    .ZN(_01549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06597_ (.A1(_01548_),
    .A2(_01549_),
    .ZN(_01550_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06598_ (.A1(_01546_),
    .A2(_01550_),
    .ZN(_01551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06599_ (.A1(_01312_),
    .A2(_01314_),
    .A3(\mem[50][2] ),
    .ZN(_01552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06600_ (.A1(_01316_),
    .A2(_01317_),
    .A3(\mem[49][2] ),
    .ZN(_01553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06601_ (.A1(_01552_),
    .A2(_01553_),
    .ZN(_01554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06602_ (.I(_01171_),
    .Z(_01555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06603_ (.A1(_01555_),
    .A2(\mem[55][2] ),
    .ZN(_01556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06604_ (.I(_01255_),
    .Z(_01557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06605_ (.A1(_01323_),
    .A2(_01557_),
    .A3(\mem[48][2] ),
    .ZN(_01558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06606_ (.A1(_01556_),
    .A2(_01558_),
    .ZN(_01559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06607_ (.A1(_01554_),
    .A2(_01559_),
    .ZN(_01560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06608_ (.A1(_01551_),
    .A2(_01560_),
    .ZN(_01561_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06609_ (.A1(_01561_),
    .A2(_01331_),
    .ZN(_01562_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06610_ (.I(_01240_),
    .Z(_01563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06611_ (.A1(_01563_),
    .A2(_01334_),
    .A3(\mem[60][2] ),
    .ZN(_01564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06612_ (.A1(_01336_),
    .A2(_01337_),
    .A3(\mem[59][2] ),
    .ZN(_01565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06613_ (.A1(_01564_),
    .A2(_01565_),
    .ZN(_01566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06614_ (.A1(_01340_),
    .A2(_01342_),
    .A3(\mem[61][2] ),
    .ZN(_01567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06615_ (.A1(_01344_),
    .A2(\mem[62][2] ),
    .ZN(_01568_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06616_ (.A1(_01567_),
    .A2(_01568_),
    .ZN(_01569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06617_ (.A1(_01566_),
    .A2(_01569_),
    .ZN(_01570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06618_ (.I(_01255_),
    .Z(_01571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06619_ (.A1(_01348_),
    .A2(_01571_),
    .A3(\mem[58][2] ),
    .ZN(_01572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06620_ (.A1(_01351_),
    .A2(_01352_),
    .A3(\mem[57][2] ),
    .ZN(_01573_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06621_ (.A1(_01572_),
    .A2(_01573_),
    .ZN(_01574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06622_ (.I(_01171_),
    .Z(_01575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06623_ (.A1(_01575_),
    .A2(\mem[63][2] ),
    .ZN(_01576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06624_ (.I(_01358_),
    .Z(_01577_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06625_ (.A1(_01357_),
    .A2(_01577_),
    .A3(\mem[56][2] ),
    .ZN(_01578_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06626_ (.A1(_01576_),
    .A2(_01578_),
    .ZN(_01579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06627_ (.A1(_01574_),
    .A2(_01579_),
    .ZN(_01580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06628_ (.A1(_01570_),
    .A2(_01580_),
    .ZN(_01581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06629_ (.A1(_01581_),
    .A2(_01365_),
    .ZN(_01582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06630_ (.A1(_01562_),
    .A2(_01582_),
    .ZN(_01583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06631_ (.A1(_01543_),
    .A2(_01583_),
    .ZN(_01584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06632_ (.I(_01067_),
    .Z(_01585_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06633_ (.A1(_01585_),
    .A2(_01370_),
    .A3(\mem[4][2] ),
    .ZN(_01586_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06634_ (.A1(_01372_),
    .A2(_01373_),
    .A3(\mem[3][2] ),
    .ZN(_01587_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06635_ (.A1(_01586_),
    .A2(_01587_),
    .ZN(_01588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06636_ (.A1(_01376_),
    .A2(_01377_),
    .A3(\mem[5][2] ),
    .ZN(_01589_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06637_ (.I(_01161_),
    .Z(_01590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06638_ (.A1(_01590_),
    .A2(\mem[6][2] ),
    .ZN(_01591_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06639_ (.A1(_01589_),
    .A2(_01591_),
    .ZN(_01592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06640_ (.A1(_01588_),
    .A2(_01592_),
    .ZN(_01593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06641_ (.I(_01313_),
    .Z(_01594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06642_ (.A1(_01383_),
    .A2(_01594_),
    .A3(\mem[2][2] ),
    .ZN(_01595_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06643_ (.A1(_01386_),
    .A2(_01387_),
    .A3(\mem[1][2] ),
    .ZN(_01596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06644_ (.A1(_01595_),
    .A2(_01596_),
    .ZN(_01597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06645_ (.A1(_01390_),
    .A2(\mem[7][2] ),
    .ZN(_01598_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06646_ (.A1(_01392_),
    .A2(_01393_),
    .A3(\mem[0][2] ),
    .ZN(_01599_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06647_ (.A1(_01598_),
    .A2(_01599_),
    .ZN(_01600_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06648_ (.A1(_01597_),
    .A2(_01600_),
    .ZN(_01601_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06649_ (.A1(_01593_),
    .A2(_01601_),
    .ZN(_01602_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06650_ (.A1(_01602_),
    .A2(_01399_),
    .ZN(_01603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06651_ (.I(_01313_),
    .Z(_01604_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06652_ (.A1(_01401_),
    .A2(_01604_),
    .A3(\mem[12][2] ),
    .ZN(_01605_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06653_ (.A1(_01404_),
    .A2(_01405_),
    .A3(\mem[11][2] ),
    .ZN(_01606_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06654_ (.A1(_01605_),
    .A2(_01606_),
    .ZN(_01607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06655_ (.I(_01066_),
    .Z(_01608_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06656_ (.A1(_01608_),
    .A2(_01409_),
    .A3(\mem[13][2] ),
    .ZN(_01609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06657_ (.I(net98),
    .Z(_01610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06658_ (.A1(_01610_),
    .A2(\mem[14][2] ),
    .ZN(_01611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06659_ (.A1(_01609_),
    .A2(_01611_),
    .ZN(_01612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06660_ (.A1(_01607_),
    .A2(_01612_),
    .ZN(_01613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06661_ (.I(_01313_),
    .Z(_01614_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06662_ (.A1(_01415_),
    .A2(_01614_),
    .A3(\mem[10][2] ),
    .ZN(_01615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06663_ (.A1(_01418_),
    .A2(_01419_),
    .A3(\mem[9][2] ),
    .ZN(_01616_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06664_ (.A1(_01615_),
    .A2(_01616_),
    .ZN(_01617_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06665_ (.A1(_01422_),
    .A2(\mem[15][2] ),
    .ZN(_01618_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06666_ (.A1(_01424_),
    .A2(_01425_),
    .A3(\mem[8][2] ),
    .ZN(_01619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06667_ (.A1(_01618_),
    .A2(_01619_),
    .ZN(_01620_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06668_ (.A1(_01617_),
    .A2(_01620_),
    .ZN(_01621_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06669_ (.A1(_01613_),
    .A2(_01621_),
    .ZN(_01622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06670_ (.A1(_01622_),
    .A2(_01432_),
    .ZN(_01623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06671_ (.A1(_01603_),
    .A2(_01623_),
    .ZN(_01624_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06672_ (.I(_01240_),
    .Z(_01625_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06673_ (.A1(_01625_),
    .A2(_01436_),
    .A3(\mem[20][2] ),
    .ZN(_01626_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06674_ (.A1(_01438_),
    .A2(_01439_),
    .A3(\mem[19][2] ),
    .ZN(_01627_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06675_ (.A1(_01626_),
    .A2(_01627_),
    .ZN(_01628_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06676_ (.I(_01066_),
    .Z(_01629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06677_ (.A1(_01629_),
    .A2(_01443_),
    .A3(\mem[21][2] ),
    .ZN(_01630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06678_ (.I(net98),
    .Z(_01631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06679_ (.A1(_01631_),
    .A2(\mem[22][2] ),
    .ZN(_01632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06680_ (.A1(_01630_),
    .A2(_01632_),
    .ZN(_01633_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06681_ (.A1(_01628_),
    .A2(_01633_),
    .ZN(_01634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06682_ (.I(_01255_),
    .Z(_01635_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06683_ (.A1(_01449_),
    .A2(_01635_),
    .A3(\mem[18][2] ),
    .ZN(_01636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06684_ (.A1(_01452_),
    .A2(_01453_),
    .A3(\mem[17][2] ),
    .ZN(_01637_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06685_ (.A1(_01636_),
    .A2(_01637_),
    .ZN(_01638_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06686_ (.A1(_01456_),
    .A2(\mem[23][2] ),
    .ZN(_01639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06687_ (.A1(_01458_),
    .A2(_01459_),
    .A3(\mem[16][2] ),
    .ZN(_01640_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06688_ (.A1(_01639_),
    .A2(_01640_),
    .ZN(_01641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06689_ (.A1(_01638_),
    .A2(_01641_),
    .ZN(_01642_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06690_ (.A1(_01634_),
    .A2(_01642_),
    .ZN(_01643_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06691_ (.A1(_01643_),
    .A2(_01464_),
    .ZN(_01644_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06692_ (.A1(_01466_),
    .A2(_01467_),
    .A3(\mem[28][2] ),
    .ZN(_01645_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06693_ (.A1(_01196_),
    .A2(_01469_),
    .A3(_01470_),
    .A4(\mem[27][2] ),
    .ZN(_01646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06694_ (.A1(_01645_),
    .A2(_01646_),
    .ZN(_01647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06695_ (.A1(_01194_),
    .A2(_01473_),
    .A3(_01474_),
    .A4(\mem[29][2] ),
    .ZN(_01648_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06696_ (.I(_01358_),
    .Z(_01649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06697_ (.A1(_01649_),
    .A2(_01477_),
    .A3(_01478_),
    .A4(\mem[30][2] ),
    .ZN(_01650_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06698_ (.A1(_01648_),
    .A2(_01650_),
    .ZN(_01651_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06699_ (.A1(_01647_),
    .A2(_01651_),
    .ZN(_01652_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06700_ (.A1(_01482_),
    .A2(_01483_),
    .A3(_01484_),
    .A4(\mem[26][2] ),
    .ZN(_01653_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06701_ (.A1(_01486_),
    .A2(_01487_),
    .A3(\mem[25][2] ),
    .ZN(_01654_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06702_ (.A1(_01653_),
    .A2(_01654_),
    .ZN(_01655_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06703_ (.A1(_01490_),
    .A2(_01190_),
    .A3(_01491_),
    .A4(\mem[31][2] ),
    .ZN(_01656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06704_ (.I(_01358_),
    .Z(_01657_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06705_ (.A1(_01493_),
    .A2(_01657_),
    .A3(\mem[24][2] ),
    .ZN(_01658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06706_ (.A1(_01656_),
    .A2(_01658_),
    .ZN(_01659_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06707_ (.A1(_01655_),
    .A2(_01659_),
    .ZN(_01660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06708_ (.A1(_01652_),
    .A2(_01660_),
    .ZN(_01661_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06709_ (.A1(_01661_),
    .A2(_01499_),
    .ZN(_01662_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06710_ (.A1(_01644_),
    .A2(_01662_),
    .ZN(_01663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06711_ (.A1(_01624_),
    .A2(_01663_),
    .ZN(_01664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06712_ (.A1(_01584_),
    .A2(_01664_),
    .ZN(_00008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06713_ (.A1(_01503_),
    .A2(_01504_),
    .A3(\mem[36][3] ),
    .ZN(_01665_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06714_ (.A1(_01237_),
    .A2(_01213_),
    .A3(\mem[35][3] ),
    .ZN(_01666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06715_ (.A1(_01665_),
    .A2(_01666_),
    .ZN(_01667_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06716_ (.A1(_01508_),
    .A2(_01242_),
    .A3(\mem[37][3] ),
    .ZN(_01668_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06717_ (.A1(_01510_),
    .A2(\mem[38][3] ),
    .ZN(_01669_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06718_ (.A1(_01668_),
    .A2(_01669_),
    .ZN(_01670_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06719_ (.A1(_01667_),
    .A2(_01670_),
    .ZN(_01671_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06720_ (.A1(_01058_),
    .A2(_01247_),
    .A3(\mem[34][3] ),
    .ZN(_01672_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06721_ (.A1(_01050_),
    .A2(_01249_),
    .A3(\mem[33][3] ),
    .ZN(_01673_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06722_ (.A1(_01672_),
    .A2(_01673_),
    .ZN(_01674_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06723_ (.A1(_01173_),
    .A2(\mem[39][3] ),
    .ZN(_01675_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06724_ (.A1(_01254_),
    .A2(_01256_),
    .A3(\mem[32][3] ),
    .ZN(_01676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06725_ (.A1(_01675_),
    .A2(_01676_),
    .ZN(_01677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06726_ (.A1(_01674_),
    .A2(_01677_),
    .ZN(_01678_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06727_ (.A1(_01671_),
    .A2(_01678_),
    .ZN(_01679_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06728_ (.A1(_01679_),
    .A2(_01261_),
    .ZN(_01680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06729_ (.A1(_01263_),
    .A2(_01523_),
    .A3(\mem[44][3] ),
    .ZN(_01681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06730_ (.A1(_01268_),
    .A2(_01269_),
    .A3(\mem[43][3] ),
    .ZN(_01682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06731_ (.A1(_01681_),
    .A2(_01682_),
    .ZN(_01683_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06732_ (.A1(_01272_),
    .A2(_01273_),
    .A3(\mem[45][3] ),
    .ZN(_01684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06733_ (.A1(_01275_),
    .A2(\mem[46][3] ),
    .ZN(_01685_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06734_ (.A1(_01684_),
    .A2(_01685_),
    .ZN(_01686_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06735_ (.A1(_01683_),
    .A2(_01686_),
    .ZN(_01687_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06736_ (.A1(_01279_),
    .A2(_01531_),
    .A3(\mem[42][3] ),
    .ZN(_01688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06737_ (.A1(_01282_),
    .A2(_01283_),
    .A3(\mem[41][3] ),
    .ZN(_01689_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06738_ (.A1(_01688_),
    .A2(_01689_),
    .ZN(_01690_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06739_ (.A1(_01535_),
    .A2(\mem[47][3] ),
    .ZN(_01691_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06740_ (.A1(_01288_),
    .A2(_01537_),
    .A3(\mem[40][3] ),
    .ZN(_01692_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06741_ (.A1(_01691_),
    .A2(_01692_),
    .ZN(_01693_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06742_ (.A1(_01690_),
    .A2(_01693_),
    .ZN(_01694_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06743_ (.A1(_01687_),
    .A2(_01694_),
    .ZN(_01695_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06744_ (.A1(_01695_),
    .A2(_01294_),
    .ZN(_01696_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06745_ (.A1(_01680_),
    .A2(_01696_),
    .ZN(_01697_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06746_ (.A1(_01297_),
    .A2(_01298_),
    .A3(\mem[52][3] ),
    .ZN(_01698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06747_ (.A1(_01300_),
    .A2(_01301_),
    .A3(\mem[51][3] ),
    .ZN(_01699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06748_ (.A1(_01698_),
    .A2(_01699_),
    .ZN(_01700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06749_ (.A1(_01547_),
    .A2(_01306_),
    .A3(\mem[53][3] ),
    .ZN(_01701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06750_ (.A1(_01308_),
    .A2(\mem[54][3] ),
    .ZN(_01702_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06751_ (.A1(_01701_),
    .A2(_01702_),
    .ZN(_01703_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06752_ (.A1(_01700_),
    .A2(_01703_),
    .ZN(_01704_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06753_ (.A1(_01312_),
    .A2(_01314_),
    .A3(\mem[50][3] ),
    .ZN(_01705_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06754_ (.A1(_01316_),
    .A2(_01317_),
    .A3(\mem[49][3] ),
    .ZN(_01706_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06755_ (.A1(_01705_),
    .A2(_01706_),
    .ZN(_01707_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06756_ (.A1(_01555_),
    .A2(\mem[55][3] ),
    .ZN(_01708_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06757_ (.A1(_01323_),
    .A2(_01557_),
    .A3(\mem[48][3] ),
    .ZN(_01709_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06758_ (.A1(_01708_),
    .A2(_01709_),
    .ZN(_01710_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06759_ (.A1(_01707_),
    .A2(_01710_),
    .ZN(_01711_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06760_ (.A1(_01704_),
    .A2(_01711_),
    .ZN(_01712_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06761_ (.A1(_01712_),
    .A2(_01331_),
    .ZN(_01713_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06762_ (.A1(_01563_),
    .A2(_01334_),
    .A3(\mem[60][3] ),
    .ZN(_01714_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06763_ (.A1(_01336_),
    .A2(_01337_),
    .A3(\mem[59][3] ),
    .ZN(_01715_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06764_ (.A1(_01714_),
    .A2(_01715_),
    .ZN(_01716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06765_ (.A1(_01340_),
    .A2(_01342_),
    .A3(\mem[61][3] ),
    .ZN(_01717_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06766_ (.A1(_01344_),
    .A2(\mem[62][3] ),
    .ZN(_01718_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06767_ (.A1(_01717_),
    .A2(_01718_),
    .ZN(_01719_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06768_ (.A1(_01716_),
    .A2(_01719_),
    .ZN(_01720_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06769_ (.A1(_01348_),
    .A2(_01571_),
    .A3(\mem[58][3] ),
    .ZN(_01721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06770_ (.A1(_01351_),
    .A2(_01352_),
    .A3(\mem[57][3] ),
    .ZN(_01722_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06771_ (.A1(_01721_),
    .A2(_01722_),
    .ZN(_01723_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06772_ (.A1(_01575_),
    .A2(\mem[63][3] ),
    .ZN(_01724_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06773_ (.A1(_01357_),
    .A2(_01577_),
    .A3(\mem[56][3] ),
    .ZN(_01725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06774_ (.A1(_01724_),
    .A2(_01725_),
    .ZN(_01726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06775_ (.A1(_01723_),
    .A2(_01726_),
    .ZN(_01727_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06776_ (.A1(_01720_),
    .A2(_01727_),
    .ZN(_01728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06777_ (.A1(_01728_),
    .A2(_01365_),
    .ZN(_01729_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06778_ (.A1(_01713_),
    .A2(_01729_),
    .ZN(_01730_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06779_ (.A1(_01697_),
    .A2(_01730_),
    .ZN(_01731_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06780_ (.A1(_01585_),
    .A2(_01370_),
    .A3(\mem[4][3] ),
    .ZN(_01732_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06781_ (.A1(_01372_),
    .A2(_01373_),
    .A3(\mem[3][3] ),
    .ZN(_01733_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06782_ (.A1(_01732_),
    .A2(_01733_),
    .ZN(_01734_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06783_ (.A1(_01376_),
    .A2(_01377_),
    .A3(\mem[5][3] ),
    .ZN(_01735_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06784_ (.A1(_01590_),
    .A2(\mem[6][3] ),
    .ZN(_01736_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06785_ (.A1(_01735_),
    .A2(_01736_),
    .ZN(_01737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06786_ (.A1(_01734_),
    .A2(_01737_),
    .ZN(_01738_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06787_ (.A1(_01383_),
    .A2(_01594_),
    .A3(\mem[2][3] ),
    .ZN(_01739_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06788_ (.A1(_01386_),
    .A2(_01387_),
    .A3(\mem[1][3] ),
    .ZN(_01740_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06789_ (.A1(_01739_),
    .A2(_01740_),
    .ZN(_01741_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06790_ (.A1(_01390_),
    .A2(\mem[7][3] ),
    .ZN(_01742_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06791_ (.A1(_01392_),
    .A2(_01393_),
    .A3(\mem[0][3] ),
    .ZN(_01743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06792_ (.A1(_01742_),
    .A2(_01743_),
    .ZN(_01744_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06793_ (.A1(_01741_),
    .A2(_01744_),
    .ZN(_01745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06794_ (.A1(_01738_),
    .A2(_01745_),
    .ZN(_01746_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06795_ (.A1(_01746_),
    .A2(_01399_),
    .ZN(_01747_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06796_ (.A1(_01401_),
    .A2(_01604_),
    .A3(\mem[12][3] ),
    .ZN(_01748_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06797_ (.A1(_01404_),
    .A2(_01405_),
    .A3(\mem[11][3] ),
    .ZN(_01749_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06798_ (.A1(_01748_),
    .A2(_01749_),
    .ZN(_01750_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06799_ (.A1(_01608_),
    .A2(_01409_),
    .A3(\mem[13][3] ),
    .ZN(_01751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06800_ (.A1(_01610_),
    .A2(\mem[14][3] ),
    .ZN(_01752_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06801_ (.A1(_01751_),
    .A2(_01752_),
    .ZN(_01753_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06802_ (.A1(_01750_),
    .A2(_01753_),
    .ZN(_01754_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06803_ (.A1(_01415_),
    .A2(_01614_),
    .A3(\mem[10][3] ),
    .ZN(_01755_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06804_ (.A1(_01418_),
    .A2(_01419_),
    .A3(\mem[9][3] ),
    .ZN(_01756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06805_ (.A1(_01755_),
    .A2(_01756_),
    .ZN(_01757_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06806_ (.A1(_01422_),
    .A2(\mem[15][3] ),
    .ZN(_01758_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06807_ (.A1(_01424_),
    .A2(_01425_),
    .A3(\mem[8][3] ),
    .ZN(_01759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06808_ (.A1(_01758_),
    .A2(_01759_),
    .ZN(_01760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06809_ (.A1(_01757_),
    .A2(_01760_),
    .ZN(_01761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06810_ (.A1(_01754_),
    .A2(_01761_),
    .ZN(_01762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06811_ (.A1(_01762_),
    .A2(_01432_),
    .ZN(_01763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06812_ (.A1(_01747_),
    .A2(_01763_),
    .ZN(_01764_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06813_ (.A1(_01625_),
    .A2(_01436_),
    .A3(\mem[20][3] ),
    .ZN(_01765_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06814_ (.A1(_01438_),
    .A2(_01439_),
    .A3(\mem[19][3] ),
    .ZN(_01766_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06815_ (.A1(_01765_),
    .A2(_01766_),
    .ZN(_01767_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06816_ (.A1(_01629_),
    .A2(_01443_),
    .A3(\mem[21][3] ),
    .ZN(_01768_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06817_ (.A1(_01631_),
    .A2(\mem[22][3] ),
    .ZN(_01769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06818_ (.A1(_01768_),
    .A2(_01769_),
    .ZN(_01770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06819_ (.A1(_01767_),
    .A2(_01770_),
    .ZN(_01771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06820_ (.A1(_01449_),
    .A2(_01635_),
    .A3(\mem[18][3] ),
    .ZN(_01772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06821_ (.A1(_01452_),
    .A2(_01453_),
    .A3(\mem[17][3] ),
    .ZN(_01773_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06822_ (.A1(_01772_),
    .A2(_01773_),
    .ZN(_01774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06823_ (.A1(_01456_),
    .A2(\mem[23][3] ),
    .ZN(_01775_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06824_ (.A1(_01458_),
    .A2(_01459_),
    .A3(\mem[16][3] ),
    .ZN(_01776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06825_ (.A1(_01775_),
    .A2(_01776_),
    .ZN(_01777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06826_ (.A1(_01774_),
    .A2(_01777_),
    .ZN(_01778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06827_ (.A1(_01771_),
    .A2(_01778_),
    .ZN(_01779_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06828_ (.A1(_01779_),
    .A2(_01464_),
    .ZN(_01780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06829_ (.A1(_01466_),
    .A2(_01467_),
    .A3(\mem[28][3] ),
    .ZN(_01781_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06830_ (.I(_01153_),
    .Z(_01782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06831_ (.A1(_01196_),
    .A2(_01469_),
    .A3(_01782_),
    .A4(\mem[27][3] ),
    .ZN(_01783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06832_ (.A1(_01781_),
    .A2(_01783_),
    .ZN(_01784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06833_ (.A1(_01194_),
    .A2(_01473_),
    .A3(_01474_),
    .A4(\mem[29][3] ),
    .ZN(_01785_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06834_ (.I(_01153_),
    .Z(_01786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06835_ (.A1(_01649_),
    .A2(_01786_),
    .A3(_01478_),
    .A4(\mem[30][3] ),
    .ZN(_01787_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06836_ (.A1(_01785_),
    .A2(_01787_),
    .ZN(_01788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06837_ (.A1(_01784_),
    .A2(_01788_),
    .ZN(_01789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06838_ (.I(_01065_),
    .Z(_01790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06839_ (.A1(_01482_),
    .A2(_01790_),
    .A3(_01484_),
    .A4(\mem[26][3] ),
    .ZN(_01791_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06840_ (.A1(_01486_),
    .A2(_01487_),
    .A3(\mem[25][3] ),
    .ZN(_01792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06841_ (.A1(_01791_),
    .A2(_01792_),
    .ZN(_01793_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06842_ (.A1(_01490_),
    .A2(_01190_),
    .A3(_01491_),
    .A4(\mem[31][3] ),
    .ZN(_01794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06843_ (.A1(_01493_),
    .A2(_01657_),
    .A3(\mem[24][3] ),
    .ZN(_01795_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06844_ (.A1(_01794_),
    .A2(_01795_),
    .ZN(_01796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06845_ (.A1(_01793_),
    .A2(_01796_),
    .ZN(_01797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06846_ (.A1(_01789_),
    .A2(_01797_),
    .ZN(_01798_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06847_ (.A1(_01798_),
    .A2(_01499_),
    .ZN(_01799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06848_ (.A1(_01780_),
    .A2(_01799_),
    .ZN(_01800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06849_ (.A1(_01764_),
    .A2(_01800_),
    .ZN(_01801_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06850_ (.A1(_01731_),
    .A2(_01801_),
    .ZN(_00009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06851_ (.A1(_01503_),
    .A2(_01504_),
    .A3(\mem[36][4] ),
    .ZN(_01802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06852_ (.A1(_01237_),
    .A2(_01213_),
    .A3(\mem[35][4] ),
    .ZN(_01803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06853_ (.A1(_01802_),
    .A2(_01803_),
    .ZN(_01804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06854_ (.A1(_01508_),
    .A2(_01242_),
    .A3(\mem[37][4] ),
    .ZN(_01805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06855_ (.A1(_01510_),
    .A2(\mem[38][4] ),
    .ZN(_01806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06856_ (.A1(_01805_),
    .A2(_01806_),
    .ZN(_01807_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06857_ (.A1(_01804_),
    .A2(_01807_),
    .ZN(_01808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06858_ (.A1(_01058_),
    .A2(_01247_),
    .A3(\mem[34][4] ),
    .ZN(_01809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06859_ (.I(_01121_),
    .Z(_01810_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06860_ (.A1(_01050_),
    .A2(_01810_),
    .A3(\mem[33][4] ),
    .ZN(_01811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06861_ (.A1(_01809_),
    .A2(_01811_),
    .ZN(_01812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06862_ (.A1(_01173_),
    .A2(\mem[39][4] ),
    .ZN(_01813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06863_ (.A1(_01254_),
    .A2(_01256_),
    .A3(\mem[32][4] ),
    .ZN(_01814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06864_ (.A1(_01813_),
    .A2(_01814_),
    .ZN(_01815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06865_ (.A1(_01812_),
    .A2(_01815_),
    .ZN(_01816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06866_ (.A1(_01808_),
    .A2(_01816_),
    .ZN(_01817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06867_ (.A1(_01817_),
    .A2(_01261_),
    .ZN(_01818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06868_ (.A1(_01263_),
    .A2(_01523_),
    .A3(\mem[44][4] ),
    .ZN(_01819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06869_ (.I(_01121_),
    .Z(_01820_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06870_ (.A1(_01268_),
    .A2(_01820_),
    .A3(\mem[43][4] ),
    .ZN(_01821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06871_ (.A1(_01819_),
    .A2(_01821_),
    .ZN(_01822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06872_ (.I(_01212_),
    .Z(_01823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06873_ (.A1(_01272_),
    .A2(_01823_),
    .A3(\mem[45][4] ),
    .ZN(_01824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06874_ (.A1(_01275_),
    .A2(\mem[46][4] ),
    .ZN(_01825_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06875_ (.A1(_01824_),
    .A2(_01825_),
    .ZN(_01826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06876_ (.A1(_01822_),
    .A2(_01826_),
    .ZN(_01827_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06877_ (.A1(_01279_),
    .A2(_01531_),
    .A3(\mem[42][4] ),
    .ZN(_01828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06878_ (.I(_01212_),
    .Z(_01829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06879_ (.A1(_01282_),
    .A2(_01829_),
    .A3(\mem[41][4] ),
    .ZN(_01830_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06880_ (.A1(_01828_),
    .A2(_01830_),
    .ZN(_01831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06881_ (.A1(_01535_),
    .A2(\mem[47][4] ),
    .ZN(_01832_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06882_ (.A1(_01288_),
    .A2(_01537_),
    .A3(\mem[40][4] ),
    .ZN(_01833_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06883_ (.A1(_01832_),
    .A2(_01833_),
    .ZN(_01834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06884_ (.A1(_01831_),
    .A2(_01834_),
    .ZN(_01835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06885_ (.A1(_01827_),
    .A2(_01835_),
    .ZN(_01836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06886_ (.A1(_01836_),
    .A2(_01294_),
    .ZN(_01837_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06887_ (.A1(_01818_),
    .A2(_01837_),
    .ZN(_01838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06888_ (.A1(_01297_),
    .A2(_01298_),
    .A3(\mem[52][4] ),
    .ZN(_01839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06889_ (.A1(_01300_),
    .A2(_01301_),
    .A3(\mem[51][4] ),
    .ZN(_01840_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06890_ (.A1(_01839_),
    .A2(_01840_),
    .ZN(_01841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06891_ (.A1(_01547_),
    .A2(_01306_),
    .A3(\mem[53][4] ),
    .ZN(_01842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06892_ (.A1(_01308_),
    .A2(\mem[54][4] ),
    .ZN(_01843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06893_ (.A1(_01842_),
    .A2(_01843_),
    .ZN(_01844_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06894_ (.A1(_01841_),
    .A2(_01844_),
    .ZN(_01845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06895_ (.A1(_01312_),
    .A2(_01314_),
    .A3(\mem[50][4] ),
    .ZN(_01846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06896_ (.A1(_01316_),
    .A2(_01317_),
    .A3(\mem[49][4] ),
    .ZN(_01847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06897_ (.A1(_01846_),
    .A2(_01847_),
    .ZN(_01848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06898_ (.A1(_01555_),
    .A2(\mem[55][4] ),
    .ZN(_01849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06899_ (.A1(_01323_),
    .A2(_01557_),
    .A3(\mem[48][4] ),
    .ZN(_01850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06900_ (.A1(_01849_),
    .A2(_01850_),
    .ZN(_01851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06901_ (.A1(_01848_),
    .A2(_01851_),
    .ZN(_01852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06902_ (.A1(_01845_),
    .A2(_01852_),
    .ZN(_01853_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06903_ (.A1(_01853_),
    .A2(_01331_),
    .ZN(_01854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06904_ (.A1(_01563_),
    .A2(_01334_),
    .A3(\mem[60][4] ),
    .ZN(_01855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06905_ (.I(_01305_),
    .Z(_01856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06906_ (.A1(_01336_),
    .A2(_01856_),
    .A3(\mem[59][4] ),
    .ZN(_01857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06907_ (.A1(_01855_),
    .A2(_01857_),
    .ZN(_01858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06908_ (.A1(_01340_),
    .A2(_01342_),
    .A3(\mem[61][4] ),
    .ZN(_01859_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06909_ (.A1(_01344_),
    .A2(\mem[62][4] ),
    .ZN(_01860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06910_ (.A1(_01859_),
    .A2(_01860_),
    .ZN(_01861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06911_ (.A1(_01858_),
    .A2(_01861_),
    .ZN(_01862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06912_ (.A1(_01348_),
    .A2(_01571_),
    .A3(\mem[58][4] ),
    .ZN(_01863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06913_ (.I(_01341_),
    .Z(_01864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06914_ (.A1(_01351_),
    .A2(_01864_),
    .A3(\mem[57][4] ),
    .ZN(_01865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06915_ (.A1(_01863_),
    .A2(_01865_),
    .ZN(_01866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06916_ (.A1(_01575_),
    .A2(\mem[63][4] ),
    .ZN(_01867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06917_ (.A1(_01357_),
    .A2(_01577_),
    .A3(\mem[56][4] ),
    .ZN(_01868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06918_ (.A1(_01867_),
    .A2(_01868_),
    .ZN(_01869_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06919_ (.A1(_01866_),
    .A2(_01869_),
    .ZN(_01870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06920_ (.A1(_01862_),
    .A2(_01870_),
    .ZN(_01871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06921_ (.A1(_01871_),
    .A2(_01365_),
    .ZN(_01872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06922_ (.A1(_01854_),
    .A2(_01872_),
    .ZN(_01873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06923_ (.A1(_01838_),
    .A2(_01873_),
    .ZN(_01874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06924_ (.A1(_01585_),
    .A2(_01370_),
    .A3(\mem[4][4] ),
    .ZN(_01875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06925_ (.A1(_01372_),
    .A2(_01373_),
    .A3(\mem[3][4] ),
    .ZN(_01876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06926_ (.A1(_01875_),
    .A2(_01876_),
    .ZN(_01877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06927_ (.I(_01212_),
    .Z(_01878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06928_ (.A1(_01376_),
    .A2(_01878_),
    .A3(\mem[5][4] ),
    .ZN(_01879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06929_ (.A1(_01590_),
    .A2(\mem[6][4] ),
    .ZN(_01880_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06930_ (.A1(_01879_),
    .A2(_01880_),
    .ZN(_01881_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06931_ (.A1(_01877_),
    .A2(_01881_),
    .ZN(_01882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06932_ (.A1(_01383_),
    .A2(_01594_),
    .A3(\mem[2][4] ),
    .ZN(_01883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06933_ (.A1(_01386_),
    .A2(_01387_),
    .A3(\mem[1][4] ),
    .ZN(_01884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06934_ (.A1(_01883_),
    .A2(_01884_),
    .ZN(_01885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06935_ (.A1(_01390_),
    .A2(\mem[7][4] ),
    .ZN(_01886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06936_ (.A1(_01392_),
    .A2(_01393_),
    .A3(\mem[0][4] ),
    .ZN(_01887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06937_ (.A1(_01886_),
    .A2(_01887_),
    .ZN(_01888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06938_ (.A1(_01885_),
    .A2(_01888_),
    .ZN(_01889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06939_ (.A1(_01882_),
    .A2(_01889_),
    .ZN(_01890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06940_ (.A1(_01890_),
    .A2(_01399_),
    .ZN(_01891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06941_ (.A1(_01401_),
    .A2(_01604_),
    .A3(\mem[12][4] ),
    .ZN(_01892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06942_ (.I(_01305_),
    .Z(_01893_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06943_ (.A1(_01404_),
    .A2(_01893_),
    .A3(\mem[11][4] ),
    .ZN(_01894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06944_ (.A1(_01892_),
    .A2(_01894_),
    .ZN(_01895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06945_ (.A1(_01608_),
    .A2(_01409_),
    .A3(\mem[13][4] ),
    .ZN(_01896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06946_ (.A1(_01610_),
    .A2(\mem[14][4] ),
    .ZN(_01897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06947_ (.A1(_01896_),
    .A2(_01897_),
    .ZN(_01898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06948_ (.A1(_01895_),
    .A2(_01898_),
    .ZN(_01899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06949_ (.A1(_01415_),
    .A2(_01614_),
    .A3(\mem[10][4] ),
    .ZN(_01900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06950_ (.A1(_01418_),
    .A2(_01419_),
    .A3(\mem[9][4] ),
    .ZN(_01901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06951_ (.A1(_01900_),
    .A2(_01901_),
    .ZN(_01902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06952_ (.A1(_01422_),
    .A2(\mem[15][4] ),
    .ZN(_01903_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06953_ (.A1(_01424_),
    .A2(_01425_),
    .A3(\mem[8][4] ),
    .ZN(_01904_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06954_ (.A1(_01903_),
    .A2(_01904_),
    .ZN(_01905_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06955_ (.A1(_01902_),
    .A2(_01905_),
    .ZN(_01906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06956_ (.A1(_01899_),
    .A2(_01906_),
    .ZN(_01907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06957_ (.A1(_01907_),
    .A2(_01432_),
    .ZN(_01908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06958_ (.A1(_01891_),
    .A2(_01908_),
    .ZN(_01909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06959_ (.A1(_01625_),
    .A2(_01436_),
    .A3(\mem[20][4] ),
    .ZN(_01910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06960_ (.I(_01305_),
    .Z(_01911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06961_ (.A1(_01438_),
    .A2(_01911_),
    .A3(\mem[19][4] ),
    .ZN(_01912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06962_ (.A1(_01910_),
    .A2(_01912_),
    .ZN(_01913_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06963_ (.A1(_01629_),
    .A2(_01443_),
    .A3(\mem[21][4] ),
    .ZN(_01914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06964_ (.A1(_01631_),
    .A2(\mem[22][4] ),
    .ZN(_01915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06965_ (.A1(_01914_),
    .A2(_01915_),
    .ZN(_01916_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06966_ (.A1(_01913_),
    .A2(_01916_),
    .ZN(_01917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06967_ (.A1(_01449_),
    .A2(_01635_),
    .A3(\mem[18][4] ),
    .ZN(_01918_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06968_ (.I(_01341_),
    .Z(_01919_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06969_ (.A1(_01452_),
    .A2(_01919_),
    .A3(\mem[17][4] ),
    .ZN(_01920_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06970_ (.A1(_01918_),
    .A2(_01920_),
    .ZN(_01921_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06971_ (.A1(_01456_),
    .A2(\mem[23][4] ),
    .ZN(_01922_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06972_ (.A1(_01458_),
    .A2(_01459_),
    .A3(\mem[16][4] ),
    .ZN(_01923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06973_ (.A1(_01922_),
    .A2(_01923_),
    .ZN(_01924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06974_ (.A1(_01921_),
    .A2(_01924_),
    .ZN(_01925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06975_ (.A1(_01917_),
    .A2(_01925_),
    .ZN(_01926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06976_ (.A1(_01926_),
    .A2(_01464_),
    .ZN(_01927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06977_ (.A1(_01466_),
    .A2(_01467_),
    .A3(\mem[28][4] ),
    .ZN(_01928_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06978_ (.I(_01043_),
    .Z(_01929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06979_ (.A1(_01196_),
    .A2(_01929_),
    .A3(_01782_),
    .A4(\mem[27][4] ),
    .ZN(_01930_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06980_ (.A1(_01928_),
    .A2(_01930_),
    .ZN(_01931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06981_ (.A1(_01194_),
    .A2(_01473_),
    .A3(_01474_),
    .A4(\mem[29][4] ),
    .ZN(_01932_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06982_ (.A1(_01649_),
    .A2(_01786_),
    .A3(_01478_),
    .A4(\mem[30][4] ),
    .ZN(_01933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06983_ (.A1(_01932_),
    .A2(_01933_),
    .ZN(_01934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06984_ (.A1(_01931_),
    .A2(_01934_),
    .ZN(_01935_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06985_ (.A1(_01482_),
    .A2(_01790_),
    .A3(_01484_),
    .A4(\mem[26][4] ),
    .ZN(_01936_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06986_ (.I(_01341_),
    .Z(_01937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06987_ (.A1(_01486_),
    .A2(_01937_),
    .A3(\mem[25][4] ),
    .ZN(_01938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06988_ (.A1(_01936_),
    .A2(_01938_),
    .ZN(_01939_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06989_ (.A1(_01490_),
    .A2(_01190_),
    .A3(_01491_),
    .A4(\mem[31][4] ),
    .ZN(_01940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06990_ (.A1(_01493_),
    .A2(_01657_),
    .A3(\mem[24][4] ),
    .ZN(_01941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06991_ (.A1(_01940_),
    .A2(_01941_),
    .ZN(_01942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06992_ (.A1(_01939_),
    .A2(_01942_),
    .ZN(_01943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06993_ (.A1(_01935_),
    .A2(_01943_),
    .ZN(_01944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06994_ (.A1(_01944_),
    .A2(_01499_),
    .ZN(_01945_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06995_ (.A1(_01927_),
    .A2(_01945_),
    .ZN(_01946_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06996_ (.A1(_01909_),
    .A2(_01946_),
    .ZN(_01947_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06997_ (.A1(_01874_),
    .A2(_01947_),
    .ZN(_00010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06998_ (.A1(_01503_),
    .A2(_01504_),
    .A3(\mem[36][5] ),
    .ZN(_01948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06999_ (.A1(_01237_),
    .A2(_01213_),
    .A3(\mem[35][5] ),
    .ZN(_01949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07000_ (.A1(_01948_),
    .A2(_01949_),
    .ZN(_01950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07001_ (.A1(_01508_),
    .A2(_01242_),
    .A3(\mem[37][5] ),
    .ZN(_01951_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07002_ (.A1(_01510_),
    .A2(\mem[38][5] ),
    .ZN(_01952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07003_ (.A1(_01951_),
    .A2(_01952_),
    .ZN(_01953_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07004_ (.A1(_01950_),
    .A2(_01953_),
    .ZN(_01954_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07005_ (.I(_01057_),
    .Z(_01955_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07006_ (.A1(_01955_),
    .A2(_01247_),
    .A3(\mem[34][5] ),
    .ZN(_01956_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07007_ (.I(_01049_),
    .Z(_01957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07008_ (.A1(_01957_),
    .A2(_01810_),
    .A3(\mem[33][5] ),
    .ZN(_01958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07009_ (.A1(_01956_),
    .A2(_01958_),
    .ZN(_01959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07010_ (.A1(_01173_),
    .A2(\mem[39][5] ),
    .ZN(_01960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07011_ (.I(_01253_),
    .Z(_01961_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07012_ (.A1(_01961_),
    .A2(_01256_),
    .A3(\mem[32][5] ),
    .ZN(_01962_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07013_ (.A1(_01960_),
    .A2(_01962_),
    .ZN(_01963_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07014_ (.A1(_01959_),
    .A2(_01963_),
    .ZN(_01964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07015_ (.A1(_01954_),
    .A2(_01964_),
    .ZN(_01965_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07016_ (.A1(_01965_),
    .A2(_01261_),
    .ZN(_01966_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07017_ (.A1(_01263_),
    .A2(_01523_),
    .A3(\mem[44][5] ),
    .ZN(_01967_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07018_ (.A1(_01268_),
    .A2(_01820_),
    .A3(\mem[43][5] ),
    .ZN(_01968_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07019_ (.A1(_01967_),
    .A2(_01968_),
    .ZN(_01969_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07020_ (.A1(_01272_),
    .A2(_01823_),
    .A3(\mem[45][5] ),
    .ZN(_01970_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07021_ (.A1(_01275_),
    .A2(\mem[46][5] ),
    .ZN(_01971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07022_ (.A1(_01970_),
    .A2(_01971_),
    .ZN(_01972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07023_ (.A1(_01969_),
    .A2(_01972_),
    .ZN(_01973_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07024_ (.I(_01267_),
    .Z(_01974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07025_ (.A1(_01974_),
    .A2(_01531_),
    .A3(\mem[42][5] ),
    .ZN(_01975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07026_ (.A1(_01282_),
    .A2(_01829_),
    .A3(\mem[41][5] ),
    .ZN(_01976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07027_ (.A1(_01975_),
    .A2(_01976_),
    .ZN(_01977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07028_ (.A1(_01535_),
    .A2(\mem[47][5] ),
    .ZN(_01978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07029_ (.A1(_01288_),
    .A2(_01537_),
    .A3(\mem[40][5] ),
    .ZN(_01979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07030_ (.A1(_01978_),
    .A2(_01979_),
    .ZN(_01980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07031_ (.A1(_01977_),
    .A2(_01980_),
    .ZN(_01981_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07032_ (.A1(_01973_),
    .A2(_01981_),
    .ZN(_01982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07033_ (.A1(_01982_),
    .A2(_01294_),
    .ZN(_01983_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07034_ (.A1(_01966_),
    .A2(_01983_),
    .ZN(_01984_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07035_ (.A1(_01297_),
    .A2(_01298_),
    .A3(\mem[52][5] ),
    .ZN(_01985_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07036_ (.A1(_01300_),
    .A2(_01301_),
    .A3(\mem[51][5] ),
    .ZN(_01986_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07037_ (.A1(_01985_),
    .A2(_01986_),
    .ZN(_01987_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07038_ (.A1(_01547_),
    .A2(_01306_),
    .A3(\mem[53][5] ),
    .ZN(_01988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07039_ (.A1(_01308_),
    .A2(\mem[54][5] ),
    .ZN(_01989_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07040_ (.A1(_01988_),
    .A2(_01989_),
    .ZN(_01990_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07041_ (.A1(_01987_),
    .A2(_01990_),
    .ZN(_01991_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07042_ (.I(_01267_),
    .Z(_01992_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07043_ (.A1(_01992_),
    .A2(_01314_),
    .A3(\mem[50][5] ),
    .ZN(_01993_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07044_ (.A1(_01316_),
    .A2(_01317_),
    .A3(\mem[49][5] ),
    .ZN(_01994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07045_ (.A1(_01993_),
    .A2(_01994_),
    .ZN(_01995_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07046_ (.A1(_01555_),
    .A2(\mem[55][5] ),
    .ZN(_01996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07047_ (.I(_01322_),
    .Z(_01997_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07048_ (.A1(_01997_),
    .A2(_01557_),
    .A3(\mem[48][5] ),
    .ZN(_01998_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07049_ (.A1(_01996_),
    .A2(_01998_),
    .ZN(_01999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07050_ (.A1(_01995_),
    .A2(_01999_),
    .ZN(_02000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07051_ (.A1(_01991_),
    .A2(_02000_),
    .ZN(_02001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07052_ (.A1(_02001_),
    .A2(_01331_),
    .ZN(_02002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07053_ (.A1(_01563_),
    .A2(_01334_),
    .A3(\mem[60][5] ),
    .ZN(_02003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07054_ (.A1(_01336_),
    .A2(_01856_),
    .A3(\mem[59][5] ),
    .ZN(_02004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07055_ (.A1(_02003_),
    .A2(_02004_),
    .ZN(_02005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07056_ (.A1(_01340_),
    .A2(_01342_),
    .A3(\mem[61][5] ),
    .ZN(_02006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07057_ (.A1(_01344_),
    .A2(\mem[62][5] ),
    .ZN(_02007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07058_ (.A1(_02006_),
    .A2(_02007_),
    .ZN(_02008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07059_ (.A1(_02005_),
    .A2(_02008_),
    .ZN(_02009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07060_ (.I(_01266_),
    .Z(_02010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07061_ (.A1(_02010_),
    .A2(_01571_),
    .A3(\mem[58][5] ),
    .ZN(_02011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07062_ (.I(_01253_),
    .Z(_02012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07063_ (.A1(_02012_),
    .A2(_01864_),
    .A3(\mem[57][5] ),
    .ZN(_02013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07064_ (.A1(_02011_),
    .A2(_02013_),
    .ZN(_02014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07065_ (.A1(_01575_),
    .A2(\mem[63][5] ),
    .ZN(_02015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07066_ (.A1(_01357_),
    .A2(_01577_),
    .A3(\mem[56][5] ),
    .ZN(_02016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07067_ (.A1(_02015_),
    .A2(_02016_),
    .ZN(_02017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07068_ (.A1(_02014_),
    .A2(_02017_),
    .ZN(_02018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07069_ (.A1(_02009_),
    .A2(_02018_),
    .ZN(_02019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07070_ (.A1(_02019_),
    .A2(_01365_),
    .ZN(_02020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07071_ (.A1(_02002_),
    .A2(_02020_),
    .ZN(_02021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07072_ (.A1(_01984_),
    .A2(_02021_),
    .ZN(_02022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07073_ (.A1(_01585_),
    .A2(_01370_),
    .A3(\mem[4][5] ),
    .ZN(_02023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07074_ (.A1(_01372_),
    .A2(_01373_),
    .A3(\mem[3][5] ),
    .ZN(_02024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07075_ (.A1(_02023_),
    .A2(_02024_),
    .ZN(_02025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07076_ (.A1(_01376_),
    .A2(_01878_),
    .A3(\mem[5][5] ),
    .ZN(_02026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07077_ (.A1(_01590_),
    .A2(\mem[6][5] ),
    .ZN(_02027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07078_ (.A1(_02026_),
    .A2(_02027_),
    .ZN(_02028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07079_ (.A1(_02025_),
    .A2(_02028_),
    .ZN(_02029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07080_ (.I(_01267_),
    .Z(_02030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07081_ (.A1(_02030_),
    .A2(_01594_),
    .A3(\mem[2][5] ),
    .ZN(_02031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07082_ (.I(_01253_),
    .Z(_02032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07083_ (.A1(_02032_),
    .A2(_01387_),
    .A3(\mem[1][5] ),
    .ZN(_02033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07084_ (.A1(_02031_),
    .A2(_02033_),
    .ZN(_02034_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07085_ (.A1(_01390_),
    .A2(\mem[7][5] ),
    .ZN(_02035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07086_ (.A1(_01392_),
    .A2(_01393_),
    .A3(\mem[0][5] ),
    .ZN(_02036_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07087_ (.A1(_02035_),
    .A2(_02036_),
    .ZN(_02037_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07088_ (.A1(_02034_),
    .A2(_02037_),
    .ZN(_02038_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07089_ (.A1(_02029_),
    .A2(_02038_),
    .ZN(_02039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07090_ (.A1(_02039_),
    .A2(_01399_),
    .ZN(_02040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07091_ (.A1(_01401_),
    .A2(_01604_),
    .A3(\mem[12][5] ),
    .ZN(_02041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07092_ (.A1(_01404_),
    .A2(_01893_),
    .A3(\mem[11][5] ),
    .ZN(_02042_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07093_ (.A1(_02041_),
    .A2(_02042_),
    .ZN(_02043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07094_ (.A1(_01608_),
    .A2(_01409_),
    .A3(\mem[13][5] ),
    .ZN(_02044_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07095_ (.A1(_01610_),
    .A2(\mem[14][5] ),
    .ZN(_02045_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07096_ (.A1(_02044_),
    .A2(_02045_),
    .ZN(_02046_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07097_ (.A1(_02043_),
    .A2(_02046_),
    .ZN(_02047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07098_ (.I(_01267_),
    .Z(_02048_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07099_ (.A1(_02048_),
    .A2(_01614_),
    .A3(\mem[10][5] ),
    .ZN(_02049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07100_ (.A1(_01418_),
    .A2(_01419_),
    .A3(\mem[9][5] ),
    .ZN(_02050_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07101_ (.A1(_02049_),
    .A2(_02050_),
    .ZN(_02051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07102_ (.A1(_01422_),
    .A2(\mem[15][5] ),
    .ZN(_02052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07103_ (.I(_01322_),
    .Z(_02053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07104_ (.A1(_02053_),
    .A2(_01425_),
    .A3(\mem[8][5] ),
    .ZN(_02054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07105_ (.A1(_02052_),
    .A2(_02054_),
    .ZN(_02055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07106_ (.A1(_02051_),
    .A2(_02055_),
    .ZN(_02056_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07107_ (.A1(_02047_),
    .A2(_02056_),
    .ZN(_02057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07108_ (.A1(_02057_),
    .A2(_01432_),
    .ZN(_02058_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07109_ (.A1(_02040_),
    .A2(_02058_),
    .ZN(_02059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07110_ (.A1(_01625_),
    .A2(_01436_),
    .A3(\mem[20][5] ),
    .ZN(_02060_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07111_ (.A1(_01438_),
    .A2(_01911_),
    .A3(\mem[19][5] ),
    .ZN(_02061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07112_ (.A1(_02060_),
    .A2(_02061_),
    .ZN(_02062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07113_ (.A1(_01629_),
    .A2(_01443_),
    .A3(\mem[21][5] ),
    .ZN(_02063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07114_ (.A1(_01631_),
    .A2(\mem[22][5] ),
    .ZN(_02064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07115_ (.A1(_02063_),
    .A2(_02064_),
    .ZN(_02065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07116_ (.A1(_02062_),
    .A2(_02065_),
    .ZN(_02066_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07117_ (.I(_01266_),
    .Z(_02067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07118_ (.A1(_02067_),
    .A2(_01635_),
    .A3(\mem[18][5] ),
    .ZN(_02068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07119_ (.I(_01253_),
    .Z(_02069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07120_ (.A1(_02069_),
    .A2(_01919_),
    .A3(\mem[17][5] ),
    .ZN(_02070_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07121_ (.A1(_02068_),
    .A2(_02070_),
    .ZN(_02071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07122_ (.A1(_01456_),
    .A2(\mem[23][5] ),
    .ZN(_02072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07123_ (.I(_01322_),
    .Z(_02073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07124_ (.A1(_02073_),
    .A2(_01459_),
    .A3(\mem[16][5] ),
    .ZN(_02074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07125_ (.A1(_02072_),
    .A2(_02074_),
    .ZN(_02075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07126_ (.A1(_02071_),
    .A2(_02075_),
    .ZN(_02076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07127_ (.A1(_02066_),
    .A2(_02076_),
    .ZN(_02077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07128_ (.A1(_02077_),
    .A2(_01464_),
    .ZN(_02078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07129_ (.A1(_01466_),
    .A2(_01467_),
    .A3(\mem[28][5] ),
    .ZN(_02079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07130_ (.A1(_01196_),
    .A2(_01929_),
    .A3(_01782_),
    .A4(\mem[27][5] ),
    .ZN(_02080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07131_ (.A1(_02079_),
    .A2(_02080_),
    .ZN(_02081_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07132_ (.A1(_01194_),
    .A2(_01473_),
    .A3(_01474_),
    .A4(\mem[29][5] ),
    .ZN(_02082_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07133_ (.A1(_01649_),
    .A2(_01786_),
    .A3(_01478_),
    .A4(\mem[30][5] ),
    .ZN(_02083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07134_ (.A1(_02082_),
    .A2(_02083_),
    .ZN(_02084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07135_ (.A1(_02081_),
    .A2(_02084_),
    .ZN(_02085_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07136_ (.A1(_01482_),
    .A2(_01790_),
    .A3(_01484_),
    .A4(\mem[26][5] ),
    .ZN(_02086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07137_ (.A1(_01486_),
    .A2(_01937_),
    .A3(\mem[25][5] ),
    .ZN(_02087_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07138_ (.A1(_02086_),
    .A2(_02087_),
    .ZN(_02088_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07139_ (.A1(_01490_),
    .A2(_01190_),
    .A3(_01491_),
    .A4(\mem[31][5] ),
    .ZN(_02089_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07140_ (.A1(_01493_),
    .A2(_01657_),
    .A3(\mem[24][5] ),
    .ZN(_02090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07141_ (.A1(_02089_),
    .A2(_02090_),
    .ZN(_02091_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07142_ (.A1(_02088_),
    .A2(_02091_),
    .ZN(_02092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07143_ (.A1(_02085_),
    .A2(_02092_),
    .ZN(_02093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07144_ (.A1(_02093_),
    .A2(_01499_),
    .ZN(_02094_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07145_ (.A1(_02078_),
    .A2(_02094_),
    .ZN(_02095_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07146_ (.A1(_02059_),
    .A2(_02095_),
    .ZN(_02096_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07147_ (.A1(_02022_),
    .A2(_02096_),
    .ZN(_00011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07148_ (.A1(_01503_),
    .A2(_01504_),
    .A3(\mem[36][6] ),
    .ZN(_02097_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07149_ (.A1(_01237_),
    .A2(_01213_),
    .A3(\mem[35][6] ),
    .ZN(_02098_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07150_ (.A1(_02097_),
    .A2(_02098_),
    .ZN(_02099_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07151_ (.A1(_01508_),
    .A2(_01242_),
    .A3(\mem[37][6] ),
    .ZN(_02100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07152_ (.A1(_01510_),
    .A2(\mem[38][6] ),
    .ZN(_02101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07153_ (.A1(_02100_),
    .A2(_02101_),
    .ZN(_02102_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07154_ (.A1(_02099_),
    .A2(_02102_),
    .ZN(_02103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07155_ (.A1(_01955_),
    .A2(_01247_),
    .A3(\mem[34][6] ),
    .ZN(_02104_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07156_ (.A1(_01957_),
    .A2(_01810_),
    .A3(\mem[33][6] ),
    .ZN(_02105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07157_ (.A1(_02104_),
    .A2(_02105_),
    .ZN(_02106_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07158_ (.A1(_01173_),
    .A2(\mem[39][6] ),
    .ZN(_02107_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07159_ (.A1(_01961_),
    .A2(_01256_),
    .A3(\mem[32][6] ),
    .ZN(_02108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07160_ (.A1(_02107_),
    .A2(_02108_),
    .ZN(_02109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07161_ (.A1(_02106_),
    .A2(_02109_),
    .ZN(_02110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07162_ (.A1(_02103_),
    .A2(_02110_),
    .ZN(_02111_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07163_ (.A1(_02111_),
    .A2(_01261_),
    .ZN(_02112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07164_ (.A1(_01263_),
    .A2(_01523_),
    .A3(\mem[44][6] ),
    .ZN(_02113_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07165_ (.A1(_01268_),
    .A2(_01820_),
    .A3(\mem[43][6] ),
    .ZN(_02114_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07166_ (.A1(_02113_),
    .A2(_02114_),
    .ZN(_02115_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07167_ (.A1(_01272_),
    .A2(_01823_),
    .A3(\mem[45][6] ),
    .ZN(_02116_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07168_ (.A1(_01275_),
    .A2(\mem[46][6] ),
    .ZN(_02117_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07169_ (.A1(_02116_),
    .A2(_02117_),
    .ZN(_02118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07170_ (.A1(_02115_),
    .A2(_02118_),
    .ZN(_02119_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07171_ (.A1(_01974_),
    .A2(_01531_),
    .A3(\mem[42][6] ),
    .ZN(_02120_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07172_ (.A1(_01282_),
    .A2(_01829_),
    .A3(\mem[41][6] ),
    .ZN(_02121_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07173_ (.A1(_02120_),
    .A2(_02121_),
    .ZN(_02122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07174_ (.A1(_01535_),
    .A2(\mem[47][6] ),
    .ZN(_02123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07175_ (.A1(_01288_),
    .A2(_01537_),
    .A3(\mem[40][6] ),
    .ZN(_02124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07176_ (.A1(_02123_),
    .A2(_02124_),
    .ZN(_02125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07177_ (.A1(_02122_),
    .A2(_02125_),
    .ZN(_02126_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07178_ (.A1(_02119_),
    .A2(_02126_),
    .ZN(_02127_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07179_ (.A1(_02127_),
    .A2(_01294_),
    .ZN(_02128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07180_ (.A1(_02112_),
    .A2(_02128_),
    .ZN(_02129_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07181_ (.A1(_01297_),
    .A2(_01298_),
    .A3(\mem[52][6] ),
    .ZN(_02130_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07182_ (.A1(_01300_),
    .A2(_01301_),
    .A3(\mem[51][6] ),
    .ZN(_02131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07183_ (.A1(_02130_),
    .A2(_02131_),
    .ZN(_02132_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07184_ (.A1(_01547_),
    .A2(_01306_),
    .A3(\mem[53][6] ),
    .ZN(_02133_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07185_ (.A1(_01308_),
    .A2(\mem[54][6] ),
    .ZN(_02134_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07186_ (.A1(_02133_),
    .A2(_02134_),
    .ZN(_02135_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07187_ (.A1(_02132_),
    .A2(_02135_),
    .ZN(_02136_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07188_ (.A1(_01992_),
    .A2(_01314_),
    .A3(\mem[50][6] ),
    .ZN(_02137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07189_ (.A1(_01316_),
    .A2(_01317_),
    .A3(\mem[49][6] ),
    .ZN(_02138_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07190_ (.A1(_02137_),
    .A2(_02138_),
    .ZN(_02139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07191_ (.A1(_01555_),
    .A2(\mem[55][6] ),
    .ZN(_02140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07192_ (.A1(_01997_),
    .A2(_01557_),
    .A3(\mem[48][6] ),
    .ZN(_02141_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07193_ (.A1(_02140_),
    .A2(_02141_),
    .ZN(_02142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07194_ (.A1(_02139_),
    .A2(_02142_),
    .ZN(_02143_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07195_ (.A1(_02136_),
    .A2(_02143_),
    .ZN(_02144_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07196_ (.A1(_02144_),
    .A2(_01331_),
    .ZN(_02145_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07197_ (.A1(_01563_),
    .A2(_01334_),
    .A3(\mem[60][6] ),
    .ZN(_02146_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07198_ (.A1(_01336_),
    .A2(_01856_),
    .A3(\mem[59][6] ),
    .ZN(_02147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07199_ (.A1(_02146_),
    .A2(_02147_),
    .ZN(_02148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07200_ (.A1(_01340_),
    .A2(_01342_),
    .A3(\mem[61][6] ),
    .ZN(_02149_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07201_ (.A1(_01344_),
    .A2(\mem[62][6] ),
    .ZN(_02150_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07202_ (.A1(_02149_),
    .A2(_02150_),
    .ZN(_02151_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07203_ (.A1(_02148_),
    .A2(_02151_),
    .ZN(_02152_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07204_ (.A1(_02010_),
    .A2(_01571_),
    .A3(\mem[58][6] ),
    .ZN(_02153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07205_ (.A1(_02012_),
    .A2(_01864_),
    .A3(\mem[57][6] ),
    .ZN(_02154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07206_ (.A1(_02153_),
    .A2(_02154_),
    .ZN(_02155_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07207_ (.A1(_01575_),
    .A2(\mem[63][6] ),
    .ZN(_02156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07208_ (.A1(_01357_),
    .A2(_01577_),
    .A3(\mem[56][6] ),
    .ZN(_02157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07209_ (.A1(_02156_),
    .A2(_02157_),
    .ZN(_02158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07210_ (.A1(_02155_),
    .A2(_02158_),
    .ZN(_02159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07211_ (.A1(_02152_),
    .A2(_02159_),
    .ZN(_02160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07212_ (.A1(_02160_),
    .A2(_01365_),
    .ZN(_02161_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07213_ (.A1(_02145_),
    .A2(_02161_),
    .ZN(_02162_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07214_ (.A1(_02129_),
    .A2(_02162_),
    .ZN(_02163_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07215_ (.A1(_01585_),
    .A2(_01370_),
    .A3(\mem[4][6] ),
    .ZN(_02164_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07216_ (.A1(_01372_),
    .A2(_01373_),
    .A3(\mem[3][6] ),
    .ZN(_02165_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07217_ (.A1(_02164_),
    .A2(_02165_),
    .ZN(_02166_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07218_ (.A1(_01376_),
    .A2(_01878_),
    .A3(\mem[5][6] ),
    .ZN(_02167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07219_ (.A1(_01590_),
    .A2(\mem[6][6] ),
    .ZN(_02168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07220_ (.A1(_02167_),
    .A2(_02168_),
    .ZN(_02169_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07221_ (.A1(_02166_),
    .A2(_02169_),
    .ZN(_02170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07222_ (.A1(_02030_),
    .A2(_01594_),
    .A3(\mem[2][6] ),
    .ZN(_02171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07223_ (.A1(_02032_),
    .A2(_01387_),
    .A3(\mem[1][6] ),
    .ZN(_02172_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07224_ (.A1(_02171_),
    .A2(_02172_),
    .ZN(_02173_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07225_ (.A1(_01390_),
    .A2(\mem[7][6] ),
    .ZN(_02174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07226_ (.A1(_01392_),
    .A2(_01393_),
    .A3(\mem[0][6] ),
    .ZN(_02175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07227_ (.A1(_02174_),
    .A2(_02175_),
    .ZN(_02176_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07228_ (.A1(_02173_),
    .A2(_02176_),
    .ZN(_02177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07229_ (.A1(_02170_),
    .A2(_02177_),
    .ZN(_02178_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07230_ (.A1(_02178_),
    .A2(_01399_),
    .ZN(_02179_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07231_ (.A1(_01401_),
    .A2(_01604_),
    .A3(\mem[12][6] ),
    .ZN(_02180_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07232_ (.A1(_01404_),
    .A2(_01893_),
    .A3(\mem[11][6] ),
    .ZN(_02181_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07233_ (.A1(_02180_),
    .A2(_02181_),
    .ZN(_02182_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07234_ (.A1(_01608_),
    .A2(_01409_),
    .A3(\mem[13][6] ),
    .ZN(_02183_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07235_ (.A1(_01610_),
    .A2(\mem[14][6] ),
    .ZN(_02184_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07236_ (.A1(_02183_),
    .A2(_02184_),
    .ZN(_02185_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07237_ (.A1(_02182_),
    .A2(_02185_),
    .ZN(_02186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07238_ (.A1(_02048_),
    .A2(_01614_),
    .A3(\mem[10][6] ),
    .ZN(_02187_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07239_ (.A1(_01418_),
    .A2(_01419_),
    .A3(\mem[9][6] ),
    .ZN(_02188_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07240_ (.A1(_02187_),
    .A2(_02188_),
    .ZN(_02189_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07241_ (.A1(_01422_),
    .A2(\mem[15][6] ),
    .ZN(_02190_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07242_ (.A1(_02053_),
    .A2(_01425_),
    .A3(\mem[8][6] ),
    .ZN(_02191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07243_ (.A1(_02190_),
    .A2(_02191_),
    .ZN(_02192_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07244_ (.A1(_02189_),
    .A2(_02192_),
    .ZN(_02193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07245_ (.A1(_02186_),
    .A2(_02193_),
    .ZN(_02194_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07246_ (.A1(_02194_),
    .A2(_01432_),
    .ZN(_02195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07247_ (.A1(_02179_),
    .A2(_02195_),
    .ZN(_02196_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07248_ (.A1(_01625_),
    .A2(_01436_),
    .A3(\mem[20][6] ),
    .ZN(_02197_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07249_ (.A1(_01438_),
    .A2(_01911_),
    .A3(\mem[19][6] ),
    .ZN(_02198_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07250_ (.A1(_02197_),
    .A2(_02198_),
    .ZN(_02199_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07251_ (.A1(_01629_),
    .A2(_01443_),
    .A3(\mem[21][6] ),
    .ZN(_02200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07252_ (.A1(_01631_),
    .A2(\mem[22][6] ),
    .ZN(_02201_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07253_ (.A1(_02200_),
    .A2(_02201_),
    .ZN(_02202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07254_ (.A1(_02199_),
    .A2(_02202_),
    .ZN(_02203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07255_ (.A1(_02067_),
    .A2(_01635_),
    .A3(\mem[18][6] ),
    .ZN(_02204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07256_ (.A1(_02069_),
    .A2(_01919_),
    .A3(\mem[17][6] ),
    .ZN(_02205_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07257_ (.A1(_02204_),
    .A2(_02205_),
    .ZN(_02206_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07258_ (.A1(_01456_),
    .A2(\mem[23][6] ),
    .ZN(_02207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07259_ (.A1(_02073_),
    .A2(_01459_),
    .A3(\mem[16][6] ),
    .ZN(_02208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07260_ (.A1(_02207_),
    .A2(_02208_),
    .ZN(_02209_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07261_ (.A1(_02206_),
    .A2(_02209_),
    .ZN(_02210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07262_ (.A1(_02203_),
    .A2(_02210_),
    .ZN(_02211_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07263_ (.A1(_02211_),
    .A2(_01464_),
    .ZN(_02212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07264_ (.A1(_01466_),
    .A2(_01467_),
    .A3(\mem[28][6] ),
    .ZN(_02213_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07265_ (.A1(_01196_),
    .A2(_01929_),
    .A3(_01782_),
    .A4(\mem[27][6] ),
    .ZN(_02214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07266_ (.A1(_02213_),
    .A2(_02214_),
    .ZN(_02215_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07267_ (.A1(_01194_),
    .A2(_01473_),
    .A3(_01474_),
    .A4(\mem[29][6] ),
    .ZN(_02216_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07268_ (.A1(_01649_),
    .A2(_01786_),
    .A3(_01478_),
    .A4(\mem[30][6] ),
    .ZN(_02217_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07269_ (.A1(_02216_),
    .A2(_02217_),
    .ZN(_02218_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07270_ (.A1(_02215_),
    .A2(_02218_),
    .ZN(_02219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07271_ (.A1(_01482_),
    .A2(_01790_),
    .A3(_01484_),
    .A4(\mem[26][6] ),
    .ZN(_02220_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07272_ (.A1(_01486_),
    .A2(_01937_),
    .A3(\mem[25][6] ),
    .ZN(_02221_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07273_ (.A1(_02220_),
    .A2(_02221_),
    .ZN(_02222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07274_ (.I(_01047_),
    .Z(_02223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07275_ (.A1(_01490_),
    .A2(_01190_),
    .A3(_02223_),
    .A4(\mem[31][6] ),
    .ZN(_02224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07276_ (.A1(_01493_),
    .A2(_01657_),
    .A3(\mem[24][6] ),
    .ZN(_02225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07277_ (.A1(_02224_),
    .A2(_02225_),
    .ZN(_02226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07278_ (.A1(_02222_),
    .A2(_02226_),
    .ZN(_02227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07279_ (.A1(_02219_),
    .A2(_02227_),
    .ZN(_02228_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07280_ (.A1(_02228_),
    .A2(_01499_),
    .ZN(_02229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07281_ (.A1(_02212_),
    .A2(_02229_),
    .ZN(_02230_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07282_ (.A1(_02196_),
    .A2(_02230_),
    .ZN(_02231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07283_ (.A1(_02163_),
    .A2(_02231_),
    .ZN(_00012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07284_ (.A1(_01503_),
    .A2(_01504_),
    .A3(\mem[36][7] ),
    .ZN(_02232_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07285_ (.A1(_01237_),
    .A2(_01213_),
    .A3(\mem[35][7] ),
    .ZN(_02233_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07286_ (.A1(_02232_),
    .A2(_02233_),
    .ZN(_02234_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07287_ (.A1(_01508_),
    .A2(_01242_),
    .A3(\mem[37][7] ),
    .ZN(_02235_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07288_ (.A1(_01510_),
    .A2(\mem[38][7] ),
    .ZN(_02236_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07289_ (.A1(_02235_),
    .A2(_02236_),
    .ZN(_02237_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07290_ (.A1(_02234_),
    .A2(_02237_),
    .ZN(_02238_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07291_ (.A1(_01955_),
    .A2(_01264_),
    .A3(\mem[34][7] ),
    .ZN(_02239_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07292_ (.A1(_01957_),
    .A2(_01810_),
    .A3(\mem[33][7] ),
    .ZN(_02240_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07293_ (.A1(_02239_),
    .A2(_02240_),
    .ZN(_02241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07294_ (.A1(_01286_),
    .A2(\mem[39][7] ),
    .ZN(_02242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07295_ (.A1(_01961_),
    .A2(_01450_),
    .A3(\mem[32][7] ),
    .ZN(_02243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07296_ (.A1(_02242_),
    .A2(_02243_),
    .ZN(_02244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07297_ (.A1(_02241_),
    .A2(_02244_),
    .ZN(_02245_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07298_ (.A1(_02238_),
    .A2(_02245_),
    .ZN(_02246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07299_ (.A1(_02246_),
    .A2(_01261_),
    .ZN(_02247_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07300_ (.A1(_01369_),
    .A2(_01523_),
    .A3(\mem[44][7] ),
    .ZN(_02248_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07301_ (.A1(_01268_),
    .A2(_01820_),
    .A3(\mem[43][7] ),
    .ZN(_02249_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07302_ (.A1(_02248_),
    .A2(_02249_),
    .ZN(_02250_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07303_ (.A1(_01435_),
    .A2(_01823_),
    .A3(\mem[45][7] ),
    .ZN(_02251_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07304_ (.A1(_01379_),
    .A2(\mem[46][7] ),
    .ZN(_02252_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07305_ (.A1(_02251_),
    .A2(_02252_),
    .ZN(_02253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07306_ (.A1(_02250_),
    .A2(_02253_),
    .ZN(_02254_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07307_ (.A1(_01974_),
    .A2(_01531_),
    .A3(\mem[42][7] ),
    .ZN(_02255_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07308_ (.A1(_01282_),
    .A2(_01829_),
    .A3(\mem[41][7] ),
    .ZN(_02256_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07309_ (.A1(_02255_),
    .A2(_02256_),
    .ZN(_02257_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07310_ (.A1(_01535_),
    .A2(\mem[47][7] ),
    .ZN(_02258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07311_ (.A1(_01288_),
    .A2(_01537_),
    .A3(\mem[40][7] ),
    .ZN(_02259_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07312_ (.A1(_02258_),
    .A2(_02259_),
    .ZN(_02260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07313_ (.A1(_02257_),
    .A2(_02260_),
    .ZN(_02261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07314_ (.A1(_02254_),
    .A2(_02261_),
    .ZN(_02262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07315_ (.A1(_02262_),
    .A2(_01294_),
    .ZN(_02263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07316_ (.A1(_02247_),
    .A2(_02263_),
    .ZN(_02264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07317_ (.A1(_01241_),
    .A2(_01384_),
    .A3(\mem[52][7] ),
    .ZN(_02265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07318_ (.A1(_01300_),
    .A2(_01301_),
    .A3(\mem[51][7] ),
    .ZN(_02266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07319_ (.A1(_02265_),
    .A2(_02266_),
    .ZN(_02267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07320_ (.A1(_01547_),
    .A2(_01306_),
    .A3(\mem[53][7] ),
    .ZN(_02268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07321_ (.A1(_01411_),
    .A2(\mem[54][7] ),
    .ZN(_02269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07322_ (.A1(_02268_),
    .A2(_02269_),
    .ZN(_02270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07323_ (.A1(_02267_),
    .A2(_02270_),
    .ZN(_02271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07324_ (.A1(_01992_),
    .A2(_01402_),
    .A3(\mem[50][7] ),
    .ZN(_02272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07325_ (.A1(_01316_),
    .A2(_01317_),
    .A3(\mem[49][7] ),
    .ZN(_02273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07326_ (.A1(_02272_),
    .A2(_02273_),
    .ZN(_02274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07327_ (.A1(_01555_),
    .A2(\mem[55][7] ),
    .ZN(_02275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07328_ (.A1(_01997_),
    .A2(_01557_),
    .A3(\mem[48][7] ),
    .ZN(_02276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07329_ (.A1(_02275_),
    .A2(_02276_),
    .ZN(_02277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07330_ (.A1(_02274_),
    .A2(_02277_),
    .ZN(_02278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07331_ (.A1(_02271_),
    .A2(_02278_),
    .ZN(_02279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07332_ (.A1(_02279_),
    .A2(_01331_),
    .ZN(_02280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07333_ (.A1(_01563_),
    .A2(_01416_),
    .A3(\mem[60][7] ),
    .ZN(_02281_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07334_ (.A1(_01336_),
    .A2(_01856_),
    .A3(\mem[59][7] ),
    .ZN(_02282_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07335_ (.A1(_02281_),
    .A2(_02282_),
    .ZN(_02283_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07336_ (.A1(_01442_),
    .A2(_01342_),
    .A3(\mem[61][7] ),
    .ZN(_02284_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07337_ (.A1(_01445_),
    .A2(\mem[62][7] ),
    .ZN(_02285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07338_ (.A1(_02284_),
    .A2(_02285_),
    .ZN(_02286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07339_ (.A1(_02283_),
    .A2(_02286_),
    .ZN(_02287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07340_ (.A1(_02010_),
    .A2(_01571_),
    .A3(\mem[58][7] ),
    .ZN(_02288_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07341_ (.A1(_02012_),
    .A2(_01864_),
    .A3(\mem[57][7] ),
    .ZN(_02289_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07342_ (.A1(_02288_),
    .A2(_02289_),
    .ZN(_02290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07343_ (.A1(_01575_),
    .A2(\mem[63][7] ),
    .ZN(_02291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07344_ (.A1(_01357_),
    .A2(_01577_),
    .A3(\mem[56][7] ),
    .ZN(_02292_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07345_ (.A1(_02291_),
    .A2(_02292_),
    .ZN(_02293_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07346_ (.A1(_02290_),
    .A2(_02293_),
    .ZN(_02294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07347_ (.A1(_02287_),
    .A2(_02294_),
    .ZN(_02295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07348_ (.A1(_02295_),
    .A2(_01365_),
    .ZN(_02296_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07349_ (.A1(_02280_),
    .A2(_02296_),
    .ZN(_02297_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07350_ (.A1(_02264_),
    .A2(_02297_),
    .ZN(_02298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07351_ (.A1(_01585_),
    .A2(_01280_),
    .A3(\mem[4][7] ),
    .ZN(_02299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07352_ (.A1(_01372_),
    .A2(_01373_),
    .A3(\mem[3][7] ),
    .ZN(_02300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07353_ (.A1(_02299_),
    .A2(_02300_),
    .ZN(_02301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07354_ (.A1(_01304_),
    .A2(_01878_),
    .A3(\mem[5][7] ),
    .ZN(_02302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07355_ (.A1(_01590_),
    .A2(\mem[6][7] ),
    .ZN(_02303_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07356_ (.A1(_02302_),
    .A2(_02303_),
    .ZN(_02304_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07357_ (.A1(_02301_),
    .A2(_02304_),
    .ZN(_02305_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07358_ (.A1(_02030_),
    .A2(_01594_),
    .A3(\mem[2][7] ),
    .ZN(_02306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07359_ (.A1(_02032_),
    .A2(_01387_),
    .A3(\mem[1][7] ),
    .ZN(_02307_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07360_ (.A1(_02306_),
    .A2(_02307_),
    .ZN(_02308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07361_ (.A1(_01320_),
    .A2(\mem[7][7] ),
    .ZN(_02309_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07362_ (.A1(_01392_),
    .A2(_01324_),
    .A3(\mem[0][7] ),
    .ZN(_02310_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07363_ (.A1(_02309_),
    .A2(_02310_),
    .ZN(_02311_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07364_ (.A1(_02308_),
    .A2(_02311_),
    .ZN(_02312_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07365_ (.A1(_02305_),
    .A2(_02312_),
    .ZN(_02313_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07366_ (.A1(_02313_),
    .A2(_01399_),
    .ZN(_02314_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07367_ (.A1(_01333_),
    .A2(_01604_),
    .A3(\mem[12][7] ),
    .ZN(_02315_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07368_ (.A1(_01404_),
    .A2(_01893_),
    .A3(\mem[11][7] ),
    .ZN(_02316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07369_ (.A1(_02315_),
    .A2(_02316_),
    .ZN(_02317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07370_ (.A1(_01608_),
    .A2(_01409_),
    .A3(\mem[13][7] ),
    .ZN(_02318_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07371_ (.A1(_01610_),
    .A2(\mem[14][7] ),
    .ZN(_02319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07372_ (.A1(_02318_),
    .A2(_02319_),
    .ZN(_02320_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07373_ (.A1(_02317_),
    .A2(_02320_),
    .ZN(_02321_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07374_ (.A1(_02048_),
    .A2(_01614_),
    .A3(\mem[10][7] ),
    .ZN(_02322_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07375_ (.A1(_01418_),
    .A2(_01419_),
    .A3(\mem[9][7] ),
    .ZN(_02323_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07376_ (.A1(_02322_),
    .A2(_02323_),
    .ZN(_02324_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07377_ (.A1(_01355_),
    .A2(\mem[15][7] ),
    .ZN(_02325_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07378_ (.A1(_02053_),
    .A2(_01359_),
    .A3(\mem[8][7] ),
    .ZN(_02326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07379_ (.A1(_02325_),
    .A2(_02326_),
    .ZN(_02327_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07380_ (.A1(_02324_),
    .A2(_02327_),
    .ZN(_02328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07381_ (.A1(_02321_),
    .A2(_02328_),
    .ZN(_02329_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07382_ (.A1(_02329_),
    .A2(_01432_),
    .ZN(_02330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07383_ (.A1(_02314_),
    .A2(_02330_),
    .ZN(_02331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07384_ (.A1(_01625_),
    .A2(_01349_),
    .A3(\mem[20][7] ),
    .ZN(_02332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07385_ (.A1(_01438_),
    .A2(_01911_),
    .A3(\mem[19][7] ),
    .ZN(_02333_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07386_ (.A1(_02332_),
    .A2(_02333_),
    .ZN(_02334_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07387_ (.A1(_01629_),
    .A2(_01443_),
    .A3(\mem[21][7] ),
    .ZN(_02335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07388_ (.A1(_01631_),
    .A2(\mem[22][7] ),
    .ZN(_02336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07389_ (.A1(_02335_),
    .A2(_02336_),
    .ZN(_02337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07390_ (.A1(_02334_),
    .A2(_02337_),
    .ZN(_02338_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07391_ (.A1(_02067_),
    .A2(_01635_),
    .A3(\mem[18][7] ),
    .ZN(_02339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07392_ (.A1(_02069_),
    .A2(_01919_),
    .A3(\mem[17][7] ),
    .ZN(_02340_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07393_ (.A1(_02339_),
    .A2(_02340_),
    .ZN(_02341_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07394_ (.A1(_01172_),
    .A2(\mem[23][7] ),
    .ZN(_02342_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07395_ (.A1(_02073_),
    .A2(_01494_),
    .A3(\mem[16][7] ),
    .ZN(_02343_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07396_ (.A1(_02342_),
    .A2(_02343_),
    .ZN(_02344_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07397_ (.A1(_02341_),
    .A2(_02344_),
    .ZN(_02345_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07398_ (.A1(_02338_),
    .A2(_02345_),
    .ZN(_02346_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07399_ (.A1(_02346_),
    .A2(_01464_),
    .ZN(_02347_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07400_ (.A1(_01408_),
    .A2(_01289_),
    .A3(\mem[28][7] ),
    .ZN(_02348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07401_ (.A1(_01196_),
    .A2(_01929_),
    .A3(_01782_),
    .A4(\mem[27][7] ),
    .ZN(_02349_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07402_ (.A1(_02348_),
    .A2(_02349_),
    .ZN(_02350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07403_ (.A1(_01194_),
    .A2(_01473_),
    .A3(_01474_),
    .A4(\mem[29][7] ),
    .ZN(_02351_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07404_ (.A1(_01649_),
    .A2(_01786_),
    .A3(_01478_),
    .A4(\mem[30][7] ),
    .ZN(_02352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07405_ (.A1(_02351_),
    .A2(_02352_),
    .ZN(_02353_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07406_ (.A1(_02350_),
    .A2(_02353_),
    .ZN(_02354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07407_ (.A1(_01476_),
    .A2(_01790_),
    .A3(_01484_),
    .A4(\mem[26][7] ),
    .ZN(_02355_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07408_ (.A1(_01486_),
    .A2(_01937_),
    .A3(\mem[25][7] ),
    .ZN(_02356_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07409_ (.A1(_02355_),
    .A2(_02356_),
    .ZN(_02357_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07410_ (.A1(_01490_),
    .A2(_01190_),
    .A3(_02223_),
    .A4(\mem[31][7] ),
    .ZN(_02358_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07411_ (.A1(_01493_),
    .A2(_01657_),
    .A3(\mem[24][7] ),
    .ZN(_02359_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07412_ (.A1(_02358_),
    .A2(_02359_),
    .ZN(_02360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07413_ (.A1(_02357_),
    .A2(_02360_),
    .ZN(_02361_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07414_ (.A1(_02354_),
    .A2(_02361_),
    .ZN(_02362_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07415_ (.A1(_02362_),
    .A2(_01499_),
    .ZN(_02363_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07416_ (.A1(_02347_),
    .A2(_02363_),
    .ZN(_02364_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07417_ (.A1(_02331_),
    .A2(_02364_),
    .ZN(_02365_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07418_ (.A1(_02298_),
    .A2(_02365_),
    .ZN(_00013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07419_ (.A1(_01503_),
    .A2(_01504_),
    .A3(\mem[36][8] ),
    .ZN(_02366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07420_ (.A1(_01237_),
    .A2(_01213_),
    .A3(\mem[35][8] ),
    .ZN(_02367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07421_ (.A1(_02366_),
    .A2(_02367_),
    .ZN(_02368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07422_ (.A1(_01508_),
    .A2(_01242_),
    .A3(\mem[37][8] ),
    .ZN(_02369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07423_ (.A1(_01510_),
    .A2(\mem[38][8] ),
    .ZN(_02370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07424_ (.A1(_02369_),
    .A2(_02370_),
    .ZN(_02371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07425_ (.A1(_02368_),
    .A2(_02371_),
    .ZN(_02372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07426_ (.A1(_01955_),
    .A2(_01264_),
    .A3(\mem[34][8] ),
    .ZN(_02373_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07427_ (.A1(_01957_),
    .A2(_01810_),
    .A3(\mem[33][8] ),
    .ZN(_02374_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07428_ (.A1(_02373_),
    .A2(_02374_),
    .ZN(_02375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07429_ (.A1(_01286_),
    .A2(\mem[39][8] ),
    .ZN(_02376_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07430_ (.A1(_01961_),
    .A2(_01450_),
    .A3(\mem[32][8] ),
    .ZN(_02377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07431_ (.A1(_02376_),
    .A2(_02377_),
    .ZN(_02378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07432_ (.A1(_02375_),
    .A2(_02378_),
    .ZN(_02379_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07433_ (.A1(_02372_),
    .A2(_02379_),
    .ZN(_02380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07434_ (.A1(_02380_),
    .A2(_01261_),
    .ZN(_02381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07435_ (.A1(_01369_),
    .A2(_01523_),
    .A3(\mem[44][8] ),
    .ZN(_02382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07436_ (.A1(_01268_),
    .A2(_01820_),
    .A3(\mem[43][8] ),
    .ZN(_02383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07437_ (.A1(_02382_),
    .A2(_02383_),
    .ZN(_02384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07438_ (.A1(_01435_),
    .A2(_01823_),
    .A3(\mem[45][8] ),
    .ZN(_02385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07439_ (.A1(_01379_),
    .A2(\mem[46][8] ),
    .ZN(_02386_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07440_ (.A1(_02385_),
    .A2(_02386_),
    .ZN(_02387_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07441_ (.A1(_02384_),
    .A2(_02387_),
    .ZN(_02388_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07442_ (.A1(_01974_),
    .A2(_01531_),
    .A3(\mem[42][8] ),
    .ZN(_02389_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07443_ (.A1(_01282_),
    .A2(_01829_),
    .A3(\mem[41][8] ),
    .ZN(_02390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07444_ (.A1(_02389_),
    .A2(_02390_),
    .ZN(_02391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07445_ (.A1(_01535_),
    .A2(\mem[47][8] ),
    .ZN(_02392_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07446_ (.A1(_01288_),
    .A2(_01537_),
    .A3(\mem[40][8] ),
    .ZN(_02393_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07447_ (.A1(_02392_),
    .A2(_02393_),
    .ZN(_02394_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07448_ (.A1(_02391_),
    .A2(_02394_),
    .ZN(_02395_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07449_ (.A1(_02388_),
    .A2(_02395_),
    .ZN(_02396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07450_ (.A1(_02396_),
    .A2(_01294_),
    .ZN(_02397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07451_ (.A1(_02381_),
    .A2(_02397_),
    .ZN(_02398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07452_ (.A1(_01241_),
    .A2(_01384_),
    .A3(\mem[52][8] ),
    .ZN(_02399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07453_ (.A1(_01300_),
    .A2(_01301_),
    .A3(\mem[51][8] ),
    .ZN(_02400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07454_ (.A1(_02399_),
    .A2(_02400_),
    .ZN(_02401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07455_ (.A1(_01547_),
    .A2(_01306_),
    .A3(\mem[53][8] ),
    .ZN(_02402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07456_ (.A1(_01411_),
    .A2(\mem[54][8] ),
    .ZN(_02403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07457_ (.A1(_02402_),
    .A2(_02403_),
    .ZN(_02404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07458_ (.A1(_02401_),
    .A2(_02404_),
    .ZN(_02405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07459_ (.A1(_01992_),
    .A2(_01402_),
    .A3(\mem[50][8] ),
    .ZN(_02406_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07460_ (.A1(_01316_),
    .A2(_01317_),
    .A3(\mem[49][8] ),
    .ZN(_02407_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07461_ (.A1(_02406_),
    .A2(_02407_),
    .ZN(_02408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07462_ (.A1(_01555_),
    .A2(\mem[55][8] ),
    .ZN(_02409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07463_ (.A1(_01997_),
    .A2(_01557_),
    .A3(\mem[48][8] ),
    .ZN(_02410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07464_ (.A1(_02409_),
    .A2(_02410_),
    .ZN(_02411_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07465_ (.A1(_02408_),
    .A2(_02411_),
    .ZN(_02412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07466_ (.A1(_02405_),
    .A2(_02412_),
    .ZN(_02413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07467_ (.A1(_02413_),
    .A2(_01331_),
    .ZN(_02414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07468_ (.A1(_01563_),
    .A2(_01416_),
    .A3(\mem[60][8] ),
    .ZN(_02415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07469_ (.A1(_01336_),
    .A2(_01856_),
    .A3(\mem[59][8] ),
    .ZN(_02416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07470_ (.A1(_02415_),
    .A2(_02416_),
    .ZN(_02417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07471_ (.A1(_01442_),
    .A2(_01342_),
    .A3(\mem[61][8] ),
    .ZN(_02418_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07472_ (.A1(_01445_),
    .A2(\mem[62][8] ),
    .ZN(_02419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07473_ (.A1(_02418_),
    .A2(_02419_),
    .ZN(_02420_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07474_ (.A1(_02417_),
    .A2(_02420_),
    .ZN(_02421_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07475_ (.A1(_02010_),
    .A2(_01571_),
    .A3(\mem[58][8] ),
    .ZN(_02422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07476_ (.A1(_02012_),
    .A2(_01864_),
    .A3(\mem[57][8] ),
    .ZN(_02423_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07477_ (.A1(_02422_),
    .A2(_02423_),
    .ZN(_02424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07478_ (.A1(_01575_),
    .A2(\mem[63][8] ),
    .ZN(_02425_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07479_ (.A1(_01357_),
    .A2(_01577_),
    .A3(\mem[56][8] ),
    .ZN(_02426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07480_ (.A1(_02425_),
    .A2(_02426_),
    .ZN(_02427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07481_ (.A1(_02424_),
    .A2(_02427_),
    .ZN(_02428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07482_ (.A1(_02421_),
    .A2(_02428_),
    .ZN(_02429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07483_ (.A1(_02429_),
    .A2(_01365_),
    .ZN(_02430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07484_ (.A1(_02414_),
    .A2(_02430_),
    .ZN(_02431_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07485_ (.A1(_02398_),
    .A2(_02431_),
    .ZN(_02432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07486_ (.A1(_01585_),
    .A2(_01280_),
    .A3(\mem[4][8] ),
    .ZN(_02433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07487_ (.A1(_01372_),
    .A2(_01373_),
    .A3(\mem[3][8] ),
    .ZN(_02434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07488_ (.A1(_02433_),
    .A2(_02434_),
    .ZN(_02435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07489_ (.A1(_01304_),
    .A2(_01878_),
    .A3(\mem[5][8] ),
    .ZN(_02436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07490_ (.A1(_01590_),
    .A2(\mem[6][8] ),
    .ZN(_02437_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07491_ (.A1(_02436_),
    .A2(_02437_),
    .ZN(_02438_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07492_ (.A1(_02435_),
    .A2(_02438_),
    .ZN(_02439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07493_ (.A1(_02030_),
    .A2(_01594_),
    .A3(\mem[2][8] ),
    .ZN(_02440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07494_ (.A1(_02032_),
    .A2(_01387_),
    .A3(\mem[1][8] ),
    .ZN(_02441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07495_ (.A1(_02440_),
    .A2(_02441_),
    .ZN(_02442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07496_ (.A1(_01320_),
    .A2(\mem[7][8] ),
    .ZN(_02443_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07497_ (.A1(_01392_),
    .A2(_01324_),
    .A3(\mem[0][8] ),
    .ZN(_02444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07498_ (.A1(_02443_),
    .A2(_02444_),
    .ZN(_02445_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07499_ (.A1(_02442_),
    .A2(_02445_),
    .ZN(_02446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07500_ (.A1(_02439_),
    .A2(_02446_),
    .ZN(_02447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07501_ (.A1(_02447_),
    .A2(_01399_),
    .ZN(_02448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07502_ (.A1(_01333_),
    .A2(_01604_),
    .A3(\mem[12][8] ),
    .ZN(_02449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07503_ (.A1(_01404_),
    .A2(_01893_),
    .A3(\mem[11][8] ),
    .ZN(_02450_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07504_ (.A1(_02449_),
    .A2(_02450_),
    .ZN(_02451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07505_ (.A1(_01608_),
    .A2(_01409_),
    .A3(\mem[13][8] ),
    .ZN(_02452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07506_ (.A1(_01610_),
    .A2(\mem[14][8] ),
    .ZN(_02453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07507_ (.A1(_02452_),
    .A2(_02453_),
    .ZN(_02454_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07508_ (.A1(_02451_),
    .A2(_02454_),
    .ZN(_02455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07509_ (.A1(_02048_),
    .A2(_01614_),
    .A3(\mem[10][8] ),
    .ZN(_02456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07510_ (.A1(_01418_),
    .A2(_01419_),
    .A3(\mem[9][8] ),
    .ZN(_02457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07511_ (.A1(_02456_),
    .A2(_02457_),
    .ZN(_02458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07512_ (.A1(_01355_),
    .A2(\mem[15][8] ),
    .ZN(_02459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07513_ (.A1(_02053_),
    .A2(_01359_),
    .A3(\mem[8][8] ),
    .ZN(_02460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07514_ (.A1(_02459_),
    .A2(_02460_),
    .ZN(_02461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07515_ (.A1(_02458_),
    .A2(_02461_),
    .ZN(_02462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07516_ (.A1(_02455_),
    .A2(_02462_),
    .ZN(_02463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07517_ (.A1(_02463_),
    .A2(_01432_),
    .ZN(_02464_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07518_ (.A1(_02448_),
    .A2(_02464_),
    .ZN(_02465_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07519_ (.A1(_01625_),
    .A2(_01349_),
    .A3(\mem[20][8] ),
    .ZN(_02466_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07520_ (.A1(_01438_),
    .A2(_01911_),
    .A3(\mem[19][8] ),
    .ZN(_02467_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07521_ (.A1(_02466_),
    .A2(_02467_),
    .ZN(_02468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07522_ (.A1(_01629_),
    .A2(_01443_),
    .A3(\mem[21][8] ),
    .ZN(_02469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07523_ (.A1(_01631_),
    .A2(\mem[22][8] ),
    .ZN(_02470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07524_ (.A1(_02469_),
    .A2(_02470_),
    .ZN(_02471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07525_ (.A1(_02468_),
    .A2(_02471_),
    .ZN(_02472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07526_ (.A1(_02067_),
    .A2(_01635_),
    .A3(\mem[18][8] ),
    .ZN(_02473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07527_ (.A1(_02069_),
    .A2(_01919_),
    .A3(\mem[17][8] ),
    .ZN(_02474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07528_ (.A1(_02473_),
    .A2(_02474_),
    .ZN(_02475_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07529_ (.A1(_01172_),
    .A2(\mem[23][8] ),
    .ZN(_02476_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07530_ (.A1(_02073_),
    .A2(_01494_),
    .A3(\mem[16][8] ),
    .ZN(_02477_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07531_ (.A1(_02476_),
    .A2(_02477_),
    .ZN(_02478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07532_ (.A1(_02475_),
    .A2(_02478_),
    .ZN(_02479_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07533_ (.A1(_02472_),
    .A2(_02479_),
    .ZN(_02480_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07534_ (.A1(_02480_),
    .A2(_01464_),
    .ZN(_02481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07535_ (.A1(_01408_),
    .A2(_01289_),
    .A3(\mem[28][8] ),
    .ZN(_02482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07536_ (.A1(_01483_),
    .A2(_01929_),
    .A3(_01782_),
    .A4(\mem[27][8] ),
    .ZN(_02483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07537_ (.A1(_02482_),
    .A2(_02483_),
    .ZN(_02484_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07538_ (.A1(_01055_),
    .A2(_01473_),
    .A3(_01474_),
    .A4(\mem[29][8] ),
    .ZN(_02485_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07539_ (.A1(_01649_),
    .A2(_01786_),
    .A3(_01478_),
    .A4(\mem[30][8] ),
    .ZN(_02486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07540_ (.A1(_02485_),
    .A2(_02486_),
    .ZN(_02487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07541_ (.A1(_02484_),
    .A2(_02487_),
    .ZN(_02488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07542_ (.A1(_01476_),
    .A2(_01790_),
    .A3(_01470_),
    .A4(\mem[26][8] ),
    .ZN(_02489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07543_ (.A1(_01486_),
    .A2(_01937_),
    .A3(\mem[25][8] ),
    .ZN(_02490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07544_ (.A1(_02489_),
    .A2(_02490_),
    .ZN(_02491_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07545_ (.A1(_01490_),
    .A2(_01477_),
    .A3(_02223_),
    .A4(\mem[31][8] ),
    .ZN(_02492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07546_ (.A1(_01493_),
    .A2(_01657_),
    .A3(\mem[24][8] ),
    .ZN(_02493_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07547_ (.A1(_02492_),
    .A2(_02493_),
    .ZN(_02494_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07548_ (.A1(_02491_),
    .A2(_02494_),
    .ZN(_02495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07549_ (.A1(_02488_),
    .A2(_02495_),
    .ZN(_02496_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07550_ (.A1(_02496_),
    .A2(_01499_),
    .ZN(_02497_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07551_ (.A1(_02481_),
    .A2(_02497_),
    .ZN(_02498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07552_ (.A1(_02465_),
    .A2(_02498_),
    .ZN(_02499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07553_ (.A1(_02432_),
    .A2(_02499_),
    .ZN(_00014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07554_ (.A1(_01503_),
    .A2(_01504_),
    .A3(\mem[36][9] ),
    .ZN(_02500_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07555_ (.A1(_01237_),
    .A2(_01249_),
    .A3(\mem[35][9] ),
    .ZN(_02501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07556_ (.A1(_02500_),
    .A2(_02501_),
    .ZN(_02502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07557_ (.A1(_01508_),
    .A2(_01269_),
    .A3(\mem[37][9] ),
    .ZN(_02503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07558_ (.A1(_01510_),
    .A2(\mem[38][9] ),
    .ZN(_02504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07559_ (.A1(_02503_),
    .A2(_02504_),
    .ZN(_02505_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07560_ (.A1(_02502_),
    .A2(_02505_),
    .ZN(_02506_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07561_ (.A1(_01955_),
    .A2(_01264_),
    .A3(\mem[34][9] ),
    .ZN(_02507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07562_ (.A1(_01957_),
    .A2(_01810_),
    .A3(\mem[33][9] ),
    .ZN(_02508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07563_ (.A1(_02507_),
    .A2(_02508_),
    .ZN(_02509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07564_ (.A1(_01286_),
    .A2(\mem[39][9] ),
    .ZN(_02510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07565_ (.A1(_01961_),
    .A2(_01450_),
    .A3(\mem[32][9] ),
    .ZN(_02511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07566_ (.A1(_02510_),
    .A2(_02511_),
    .ZN(_02512_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07567_ (.A1(_02509_),
    .A2(_02512_),
    .ZN(_02513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07568_ (.A1(_02506_),
    .A2(_02513_),
    .ZN(_02514_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07569_ (.A1(_02514_),
    .A2(_01261_),
    .ZN(_02515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07570_ (.A1(_01369_),
    .A2(_01523_),
    .A3(\mem[44][9] ),
    .ZN(_02516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07571_ (.A1(_01268_),
    .A2(_01820_),
    .A3(\mem[43][9] ),
    .ZN(_02517_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07572_ (.A1(_02516_),
    .A2(_02517_),
    .ZN(_02518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07573_ (.A1(_01435_),
    .A2(_01823_),
    .A3(\mem[45][9] ),
    .ZN(_02519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07574_ (.A1(_01379_),
    .A2(\mem[46][9] ),
    .ZN(_02520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07575_ (.A1(_02519_),
    .A2(_02520_),
    .ZN(_02521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07576_ (.A1(_02518_),
    .A2(_02521_),
    .ZN(_02522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07577_ (.A1(_01974_),
    .A2(_01531_),
    .A3(\mem[42][9] ),
    .ZN(_02523_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07578_ (.A1(_01282_),
    .A2(_01829_),
    .A3(\mem[41][9] ),
    .ZN(_02524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07579_ (.A1(_02523_),
    .A2(_02524_),
    .ZN(_02525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07580_ (.A1(_01535_),
    .A2(\mem[47][9] ),
    .ZN(_02526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07581_ (.A1(_01288_),
    .A2(_01537_),
    .A3(\mem[40][9] ),
    .ZN(_02527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07582_ (.A1(_02526_),
    .A2(_02527_),
    .ZN(_02528_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07583_ (.A1(_02525_),
    .A2(_02528_),
    .ZN(_02529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07584_ (.A1(_02522_),
    .A2(_02529_),
    .ZN(_02530_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07585_ (.A1(_02530_),
    .A2(_01294_),
    .ZN(_02531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07586_ (.A1(_02515_),
    .A2(_02531_),
    .ZN(_02532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07587_ (.A1(_01241_),
    .A2(_01384_),
    .A3(\mem[52][9] ),
    .ZN(_02533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07588_ (.A1(_01300_),
    .A2(_01273_),
    .A3(\mem[51][9] ),
    .ZN(_02534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07589_ (.A1(_02533_),
    .A2(_02534_),
    .ZN(_02535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07590_ (.A1(_01547_),
    .A2(_01337_),
    .A3(\mem[53][9] ),
    .ZN(_02536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07591_ (.A1(_01411_),
    .A2(\mem[54][9] ),
    .ZN(_02537_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07592_ (.A1(_02536_),
    .A2(_02537_),
    .ZN(_02538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07593_ (.A1(_02535_),
    .A2(_02538_),
    .ZN(_02539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07594_ (.A1(_01992_),
    .A2(_01402_),
    .A3(\mem[50][9] ),
    .ZN(_02540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07595_ (.A1(_01316_),
    .A2(_01405_),
    .A3(\mem[49][9] ),
    .ZN(_02541_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07596_ (.A1(_02540_),
    .A2(_02541_),
    .ZN(_02542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07597_ (.A1(_01555_),
    .A2(\mem[55][9] ),
    .ZN(_02543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07598_ (.A1(_01997_),
    .A2(_01557_),
    .A3(\mem[48][9] ),
    .ZN(_02544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07599_ (.A1(_02543_),
    .A2(_02544_),
    .ZN(_02545_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07600_ (.A1(_02542_),
    .A2(_02545_),
    .ZN(_02546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07601_ (.A1(_02539_),
    .A2(_02546_),
    .ZN(_02547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07602_ (.A1(_02547_),
    .A2(_01331_),
    .ZN(_02548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07603_ (.A1(_01563_),
    .A2(_01416_),
    .A3(\mem[60][9] ),
    .ZN(_02549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07604_ (.A1(_01336_),
    .A2(_01856_),
    .A3(\mem[59][9] ),
    .ZN(_02550_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07605_ (.A1(_02549_),
    .A2(_02550_),
    .ZN(_02551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07606_ (.A1(_01442_),
    .A2(_01453_),
    .A3(\mem[61][9] ),
    .ZN(_02552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07607_ (.A1(_01445_),
    .A2(\mem[62][9] ),
    .ZN(_02553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07608_ (.A1(_02552_),
    .A2(_02553_),
    .ZN(_02554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07609_ (.A1(_02551_),
    .A2(_02554_),
    .ZN(_02555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07610_ (.A1(_02010_),
    .A2(_01571_),
    .A3(\mem[58][9] ),
    .ZN(_02556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07611_ (.A1(_02012_),
    .A2(_01864_),
    .A3(\mem[57][9] ),
    .ZN(_02557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07612_ (.A1(_02556_),
    .A2(_02557_),
    .ZN(_02558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07613_ (.A1(_01575_),
    .A2(\mem[63][9] ),
    .ZN(_02559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07614_ (.A1(_01357_),
    .A2(_01577_),
    .A3(\mem[56][9] ),
    .ZN(_02560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07615_ (.A1(_02559_),
    .A2(_02560_),
    .ZN(_02561_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07616_ (.A1(_02558_),
    .A2(_02561_),
    .ZN(_02562_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07617_ (.A1(_02555_),
    .A2(_02562_),
    .ZN(_02563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07618_ (.A1(_02563_),
    .A2(_01365_),
    .ZN(_02564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07619_ (.A1(_02548_),
    .A2(_02564_),
    .ZN(_02565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07620_ (.A1(_02532_),
    .A2(_02565_),
    .ZN(_02566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07621_ (.A1(_01585_),
    .A2(_01280_),
    .A3(\mem[4][9] ),
    .ZN(_02567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07622_ (.A1(_01372_),
    .A2(_01283_),
    .A3(\mem[3][9] ),
    .ZN(_02568_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07623_ (.A1(_02567_),
    .A2(_02568_),
    .ZN(_02569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07624_ (.A1(_01304_),
    .A2(_01878_),
    .A3(\mem[5][9] ),
    .ZN(_02570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07625_ (.A1(_01590_),
    .A2(\mem[6][9] ),
    .ZN(_02571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07626_ (.A1(_02570_),
    .A2(_02571_),
    .ZN(_02572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07627_ (.A1(_02569_),
    .A2(_02572_),
    .ZN(_02573_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07628_ (.A1(_02030_),
    .A2(_01594_),
    .A3(\mem[2][9] ),
    .ZN(_02574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07629_ (.A1(_02032_),
    .A2(_01377_),
    .A3(\mem[1][9] ),
    .ZN(_02575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07630_ (.A1(_02574_),
    .A2(_02575_),
    .ZN(_02576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07631_ (.A1(_01320_),
    .A2(\mem[7][9] ),
    .ZN(_02577_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07632_ (.A1(_01392_),
    .A2(_01324_),
    .A3(\mem[0][9] ),
    .ZN(_02578_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07633_ (.A1(_02577_),
    .A2(_02578_),
    .ZN(_02579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07634_ (.A1(_02576_),
    .A2(_02579_),
    .ZN(_02580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07635_ (.A1(_02573_),
    .A2(_02580_),
    .ZN(_02581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07636_ (.A1(_02581_),
    .A2(_01399_),
    .ZN(_02582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07637_ (.A1(_01333_),
    .A2(_01604_),
    .A3(\mem[12][9] ),
    .ZN(_02583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07638_ (.A1(_01404_),
    .A2(_01893_),
    .A3(\mem[11][9] ),
    .ZN(_02584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07639_ (.A1(_02583_),
    .A2(_02584_),
    .ZN(_02585_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07640_ (.A1(_01608_),
    .A2(_01352_),
    .A3(\mem[13][9] ),
    .ZN(_02586_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07641_ (.A1(_01610_),
    .A2(\mem[14][9] ),
    .ZN(_02587_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07642_ (.A1(_02586_),
    .A2(_02587_),
    .ZN(_02588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07643_ (.A1(_02585_),
    .A2(_02588_),
    .ZN(_02589_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07644_ (.A1(_02048_),
    .A2(_01614_),
    .A3(\mem[10][9] ),
    .ZN(_02590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07645_ (.A1(_01418_),
    .A2(_01439_),
    .A3(\mem[9][9] ),
    .ZN(_02591_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07646_ (.A1(_02590_),
    .A2(_02591_),
    .ZN(_02592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07647_ (.A1(_01355_),
    .A2(\mem[15][9] ),
    .ZN(_02593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07648_ (.A1(_02053_),
    .A2(_01359_),
    .A3(\mem[8][9] ),
    .ZN(_02594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07649_ (.A1(_02593_),
    .A2(_02594_),
    .ZN(_02595_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07650_ (.A1(_02592_),
    .A2(_02595_),
    .ZN(_02596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07651_ (.A1(_02589_),
    .A2(_02596_),
    .ZN(_02597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07652_ (.A1(_02597_),
    .A2(_01432_),
    .ZN(_02598_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07653_ (.A1(_02582_),
    .A2(_02598_),
    .ZN(_02599_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07654_ (.A1(_01625_),
    .A2(_01349_),
    .A3(\mem[20][9] ),
    .ZN(_02600_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07655_ (.A1(_01438_),
    .A2(_01911_),
    .A3(\mem[19][9] ),
    .ZN(_02601_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07656_ (.A1(_02600_),
    .A2(_02601_),
    .ZN(_02602_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07657_ (.A1(_01629_),
    .A2(_01487_),
    .A3(\mem[21][9] ),
    .ZN(_02603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07658_ (.A1(_01631_),
    .A2(\mem[22][9] ),
    .ZN(_02604_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07659_ (.A1(_02603_),
    .A2(_02604_),
    .ZN(_02605_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07660_ (.A1(_02602_),
    .A2(_02605_),
    .ZN(_02606_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07661_ (.A1(_02067_),
    .A2(_01635_),
    .A3(\mem[18][9] ),
    .ZN(_02607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07662_ (.A1(_02069_),
    .A2(_01919_),
    .A3(\mem[17][9] ),
    .ZN(_02608_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07663_ (.A1(_02607_),
    .A2(_02608_),
    .ZN(_02609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07664_ (.A1(_01172_),
    .A2(\mem[23][9] ),
    .ZN(_02610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07665_ (.A1(_02073_),
    .A2(_01494_),
    .A3(\mem[16][9] ),
    .ZN(_02611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07666_ (.A1(_02610_),
    .A2(_02611_),
    .ZN(_02612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07667_ (.A1(_02609_),
    .A2(_02612_),
    .ZN(_02613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07668_ (.A1(_02606_),
    .A2(_02613_),
    .ZN(_02614_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07669_ (.A1(_02614_),
    .A2(_01464_),
    .ZN(_02615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07670_ (.A1(_01408_),
    .A2(_01289_),
    .A3(\mem[28][9] ),
    .ZN(_02616_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07671_ (.A1(_01483_),
    .A2(_01929_),
    .A3(_01782_),
    .A4(\mem[27][9] ),
    .ZN(_02617_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07672_ (.A1(_02616_),
    .A2(_02617_),
    .ZN(_02618_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07673_ (.A1(_01055_),
    .A2(_01044_),
    .A3(_01474_),
    .A4(\mem[29][9] ),
    .ZN(_02619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07674_ (.A1(_01649_),
    .A2(_01786_),
    .A3(_01478_),
    .A4(\mem[30][9] ),
    .ZN(_02620_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07675_ (.A1(_02619_),
    .A2(_02620_),
    .ZN(_02621_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07676_ (.A1(_02618_),
    .A2(_02621_),
    .ZN(_02622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07677_ (.A1(_01476_),
    .A2(_01790_),
    .A3(_01470_),
    .A4(\mem[26][9] ),
    .ZN(_02623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07678_ (.A1(_01486_),
    .A2(_01937_),
    .A3(\mem[25][9] ),
    .ZN(_02624_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07679_ (.A1(_02623_),
    .A2(_02624_),
    .ZN(_02625_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07680_ (.A1(_01469_),
    .A2(_01477_),
    .A3(_02223_),
    .A4(\mem[31][9] ),
    .ZN(_02626_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07681_ (.A1(_01493_),
    .A2(_01657_),
    .A3(\mem[24][9] ),
    .ZN(_02627_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07682_ (.A1(_02626_),
    .A2(_02627_),
    .ZN(_02628_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07683_ (.A1(_02625_),
    .A2(_02628_),
    .ZN(_02629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07684_ (.A1(_02622_),
    .A2(_02629_),
    .ZN(_02630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07685_ (.A1(_02630_),
    .A2(_01499_),
    .ZN(_02631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07686_ (.A1(_02615_),
    .A2(_02631_),
    .ZN(_02632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07687_ (.A1(_02599_),
    .A2(_02632_),
    .ZN(_02633_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07688_ (.A1(_02566_),
    .A2(_02633_),
    .ZN(_00015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07689_ (.A1(_01503_),
    .A2(_01504_),
    .A3(\mem[36][10] ),
    .ZN(_02634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07690_ (.A1(_01279_),
    .A2(_01249_),
    .A3(\mem[35][10] ),
    .ZN(_02635_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07691_ (.A1(_02634_),
    .A2(_02635_),
    .ZN(_02636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07692_ (.A1(_01508_),
    .A2(_01269_),
    .A3(\mem[37][10] ),
    .ZN(_02637_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07693_ (.A1(_01510_),
    .A2(\mem[38][10] ),
    .ZN(_02638_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07694_ (.A1(_02637_),
    .A2(_02638_),
    .ZN(_02639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07695_ (.A1(_02636_),
    .A2(_02639_),
    .ZN(_02640_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07696_ (.A1(_01955_),
    .A2(_01264_),
    .A3(\mem[34][10] ),
    .ZN(_02641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07697_ (.A1(_01957_),
    .A2(_01810_),
    .A3(\mem[33][10] ),
    .ZN(_02642_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07698_ (.A1(_02641_),
    .A2(_02642_),
    .ZN(_02643_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07699_ (.A1(_01286_),
    .A2(\mem[39][10] ),
    .ZN(_02644_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07700_ (.A1(_01961_),
    .A2(_01450_),
    .A3(\mem[32][10] ),
    .ZN(_02645_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07701_ (.A1(_02644_),
    .A2(_02645_),
    .ZN(_02646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07702_ (.A1(_02643_),
    .A2(_02646_),
    .ZN(_02647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07703_ (.A1(_02640_),
    .A2(_02647_),
    .ZN(_02648_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07704_ (.A1(_02648_),
    .A2(_01261_),
    .ZN(_02649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07705_ (.A1(_01369_),
    .A2(_01523_),
    .A3(\mem[44][10] ),
    .ZN(_02650_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07706_ (.A1(_01383_),
    .A2(_01820_),
    .A3(\mem[43][10] ),
    .ZN(_02651_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07707_ (.A1(_02650_),
    .A2(_02651_),
    .ZN(_02652_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07708_ (.A1(_01435_),
    .A2(_01823_),
    .A3(\mem[45][10] ),
    .ZN(_02653_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07709_ (.A1(_01379_),
    .A2(\mem[46][10] ),
    .ZN(_02654_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07710_ (.A1(_02653_),
    .A2(_02654_),
    .ZN(_02655_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07711_ (.A1(_02652_),
    .A2(_02655_),
    .ZN(_02656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07712_ (.A1(_01974_),
    .A2(_01531_),
    .A3(\mem[42][10] ),
    .ZN(_02657_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07713_ (.A1(_01386_),
    .A2(_01829_),
    .A3(\mem[41][10] ),
    .ZN(_02658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07714_ (.A1(_02657_),
    .A2(_02658_),
    .ZN(_02659_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07715_ (.A1(_01535_),
    .A2(\mem[47][10] ),
    .ZN(_02660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07716_ (.A1(_01452_),
    .A2(_01537_),
    .A3(\mem[40][10] ),
    .ZN(_02661_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07717_ (.A1(_02660_),
    .A2(_02661_),
    .ZN(_02662_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07718_ (.A1(_02659_),
    .A2(_02662_),
    .ZN(_02663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07719_ (.A1(_02656_),
    .A2(_02663_),
    .ZN(_02664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07720_ (.A1(_02664_),
    .A2(_01294_),
    .ZN(_02665_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07721_ (.A1(_02649_),
    .A2(_02665_),
    .ZN(_02666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07722_ (.A1(_01241_),
    .A2(_01384_),
    .A3(\mem[52][10] ),
    .ZN(_02667_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07723_ (.A1(_01415_),
    .A2(_01273_),
    .A3(\mem[51][10] ),
    .ZN(_02668_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07724_ (.A1(_02667_),
    .A2(_02668_),
    .ZN(_02669_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07725_ (.A1(_01547_),
    .A2(_01337_),
    .A3(\mem[53][10] ),
    .ZN(_02670_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07726_ (.A1(_01411_),
    .A2(\mem[54][10] ),
    .ZN(_02671_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07727_ (.A1(_02670_),
    .A2(_02671_),
    .ZN(_02672_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07728_ (.A1(_02669_),
    .A2(_02672_),
    .ZN(_02673_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07729_ (.A1(_01992_),
    .A2(_01402_),
    .A3(\mem[50][10] ),
    .ZN(_02674_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07730_ (.A1(_01254_),
    .A2(_01405_),
    .A3(\mem[49][10] ),
    .ZN(_02675_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07731_ (.A1(_02674_),
    .A2(_02675_),
    .ZN(_02676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07732_ (.A1(_01555_),
    .A2(\mem[55][10] ),
    .ZN(_02677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07733_ (.A1(_01997_),
    .A2(_01557_),
    .A3(\mem[48][10] ),
    .ZN(_02678_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07734_ (.A1(_02677_),
    .A2(_02678_),
    .ZN(_02679_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07735_ (.A1(_02676_),
    .A2(_02679_),
    .ZN(_02680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07736_ (.A1(_02673_),
    .A2(_02680_),
    .ZN(_02681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07737_ (.A1(_02681_),
    .A2(_01331_),
    .ZN(_02682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07738_ (.A1(_01563_),
    .A2(_01416_),
    .A3(\mem[60][10] ),
    .ZN(_02683_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07739_ (.A1(_01449_),
    .A2(_01856_),
    .A3(\mem[59][10] ),
    .ZN(_02684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07740_ (.A1(_02683_),
    .A2(_02684_),
    .ZN(_02685_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07741_ (.A1(_01442_),
    .A2(_01453_),
    .A3(\mem[61][10] ),
    .ZN(_02686_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07742_ (.A1(_01445_),
    .A2(\mem[62][10] ),
    .ZN(_02687_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07743_ (.A1(_02686_),
    .A2(_02687_),
    .ZN(_02688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07744_ (.A1(_02685_),
    .A2(_02688_),
    .ZN(_02689_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07745_ (.A1(_02010_),
    .A2(_01571_),
    .A3(\mem[58][10] ),
    .ZN(_02690_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07746_ (.A1(_02012_),
    .A2(_01864_),
    .A3(\mem[57][10] ),
    .ZN(_02691_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07747_ (.A1(_02690_),
    .A2(_02691_),
    .ZN(_02692_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07748_ (.A1(_01575_),
    .A2(\mem[63][10] ),
    .ZN(_02693_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07749_ (.A1(_01458_),
    .A2(_01577_),
    .A3(\mem[56][10] ),
    .ZN(_02694_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07750_ (.A1(_02693_),
    .A2(_02694_),
    .ZN(_02695_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07751_ (.A1(_02692_),
    .A2(_02695_),
    .ZN(_02696_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07752_ (.A1(_02689_),
    .A2(_02696_),
    .ZN(_02697_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07753_ (.A1(_02697_),
    .A2(_01365_),
    .ZN(_02698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07754_ (.A1(_02682_),
    .A2(_02698_),
    .ZN(_02699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07755_ (.A1(_02666_),
    .A2(_02699_),
    .ZN(_02700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07756_ (.A1(_01585_),
    .A2(_01280_),
    .A3(\mem[4][10] ),
    .ZN(_02701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07757_ (.A1(_01312_),
    .A2(_01283_),
    .A3(\mem[3][10] ),
    .ZN(_02702_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07758_ (.A1(_02701_),
    .A2(_02702_),
    .ZN(_02703_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07759_ (.A1(_01304_),
    .A2(_01878_),
    .A3(\mem[5][10] ),
    .ZN(_02704_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07760_ (.A1(_01590_),
    .A2(\mem[6][10] ),
    .ZN(_02705_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07761_ (.A1(_02704_),
    .A2(_02705_),
    .ZN(_02706_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07762_ (.A1(_02703_),
    .A2(_02706_),
    .ZN(_02707_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07763_ (.A1(_02030_),
    .A2(_01594_),
    .A3(\mem[2][10] ),
    .ZN(_02708_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07764_ (.A1(_02032_),
    .A2(_01377_),
    .A3(\mem[1][10] ),
    .ZN(_02709_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07765_ (.A1(_02708_),
    .A2(_02709_),
    .ZN(_02710_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07766_ (.A1(_01320_),
    .A2(\mem[7][10] ),
    .ZN(_02711_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07767_ (.A1(_01323_),
    .A2(_01324_),
    .A3(\mem[0][10] ),
    .ZN(_02712_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07768_ (.A1(_02711_),
    .A2(_02712_),
    .ZN(_02713_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07769_ (.A1(_02710_),
    .A2(_02713_),
    .ZN(_02714_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07770_ (.A1(_02707_),
    .A2(_02714_),
    .ZN(_02715_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07771_ (.A1(_02715_),
    .A2(_01399_),
    .ZN(_02716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07772_ (.A1(_01333_),
    .A2(_01604_),
    .A3(\mem[12][10] ),
    .ZN(_02717_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07773_ (.A1(_01348_),
    .A2(_01893_),
    .A3(\mem[11][10] ),
    .ZN(_02718_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07774_ (.A1(_02717_),
    .A2(_02718_),
    .ZN(_02719_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07775_ (.A1(_01608_),
    .A2(_01352_),
    .A3(\mem[13][10] ),
    .ZN(_02720_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07776_ (.A1(_01610_),
    .A2(\mem[14][10] ),
    .ZN(_02721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07777_ (.A1(_02720_),
    .A2(_02721_),
    .ZN(_02722_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07778_ (.A1(_02719_),
    .A2(_02722_),
    .ZN(_02723_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07779_ (.A1(_02048_),
    .A2(_01614_),
    .A3(\mem[10][10] ),
    .ZN(_02724_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07780_ (.A1(_01351_),
    .A2(_01439_),
    .A3(\mem[9][10] ),
    .ZN(_02725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07781_ (.A1(_02724_),
    .A2(_02725_),
    .ZN(_02726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07782_ (.A1(_01355_),
    .A2(\mem[15][10] ),
    .ZN(_02727_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07783_ (.A1(_02053_),
    .A2(_01359_),
    .A3(\mem[8][10] ),
    .ZN(_02728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07784_ (.A1(_02727_),
    .A2(_02728_),
    .ZN(_02729_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07785_ (.A1(_02726_),
    .A2(_02729_),
    .ZN(_02730_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07786_ (.A1(_02723_),
    .A2(_02730_),
    .ZN(_02731_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07787_ (.A1(_02731_),
    .A2(_01432_),
    .ZN(_02732_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07788_ (.A1(_02716_),
    .A2(_02732_),
    .ZN(_02733_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07789_ (.A1(_01625_),
    .A2(_01349_),
    .A3(\mem[20][10] ),
    .ZN(_02734_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07790_ (.A1(_01057_),
    .A2(_01911_),
    .A3(\mem[19][10] ),
    .ZN(_02735_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07791_ (.A1(_02734_),
    .A2(_02735_),
    .ZN(_02736_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07792_ (.A1(_01629_),
    .A2(_01487_),
    .A3(\mem[21][10] ),
    .ZN(_02737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07793_ (.A1(_01631_),
    .A2(\mem[22][10] ),
    .ZN(_02738_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07794_ (.A1(_02737_),
    .A2(_02738_),
    .ZN(_02739_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07795_ (.A1(_02736_),
    .A2(_02739_),
    .ZN(_02740_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07796_ (.A1(_02067_),
    .A2(_01635_),
    .A3(\mem[18][10] ),
    .ZN(_02741_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07797_ (.A1(_02069_),
    .A2(_01919_),
    .A3(\mem[17][10] ),
    .ZN(_02742_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07798_ (.A1(_02741_),
    .A2(_02742_),
    .ZN(_02743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07799_ (.A1(_01172_),
    .A2(\mem[23][10] ),
    .ZN(_02744_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07800_ (.A1(_02073_),
    .A2(_01494_),
    .A3(\mem[16][10] ),
    .ZN(_02745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07801_ (.A1(_02744_),
    .A2(_02745_),
    .ZN(_02746_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07802_ (.A1(_02743_),
    .A2(_02746_),
    .ZN(_02747_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07803_ (.A1(_02740_),
    .A2(_02747_),
    .ZN(_02748_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07804_ (.A1(_02748_),
    .A2(_01464_),
    .ZN(_02749_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07805_ (.A1(_01408_),
    .A2(_01289_),
    .A3(\mem[28][10] ),
    .ZN(_02750_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07806_ (.A1(_01483_),
    .A2(_01929_),
    .A3(_01782_),
    .A4(\mem[27][10] ),
    .ZN(_02751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07807_ (.A1(_02750_),
    .A2(_02751_),
    .ZN(_02752_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07808_ (.A1(_01055_),
    .A2(_01044_),
    .A3(_01474_),
    .A4(\mem[29][10] ),
    .ZN(_02753_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07809_ (.A1(_01649_),
    .A2(_01786_),
    .A3(_01478_),
    .A4(\mem[30][10] ),
    .ZN(_02754_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07810_ (.A1(_02753_),
    .A2(_02754_),
    .ZN(_02755_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07811_ (.A1(_02752_),
    .A2(_02755_),
    .ZN(_02756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07812_ (.A1(_01476_),
    .A2(_01790_),
    .A3(_01470_),
    .A4(\mem[26][10] ),
    .ZN(_02757_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07813_ (.A1(_01424_),
    .A2(_01937_),
    .A3(\mem[25][10] ),
    .ZN(_02758_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07814_ (.A1(_02757_),
    .A2(_02758_),
    .ZN(_02759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07815_ (.A1(_01469_),
    .A2(_01477_),
    .A3(_02223_),
    .A4(\mem[31][10] ),
    .ZN(_02760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07816_ (.A1(_01049_),
    .A2(_01657_),
    .A3(\mem[24][10] ),
    .ZN(_02761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07817_ (.A1(_02760_),
    .A2(_02761_),
    .ZN(_02762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07818_ (.A1(_02759_),
    .A2(_02762_),
    .ZN(_02763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07819_ (.A1(_02756_),
    .A2(_02763_),
    .ZN(_02764_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07820_ (.A1(_02764_),
    .A2(_01499_),
    .ZN(_02765_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07821_ (.A1(_02749_),
    .A2(_02765_),
    .ZN(_02766_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07822_ (.A1(_02733_),
    .A2(_02766_),
    .ZN(_02767_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07823_ (.A1(_02700_),
    .A2(_02767_),
    .ZN(_00001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07824_ (.A1(_01503_),
    .A2(_01504_),
    .A3(\mem[36][11] ),
    .ZN(_02768_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07825_ (.A1(_01279_),
    .A2(_01249_),
    .A3(\mem[35][11] ),
    .ZN(_02769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07826_ (.A1(_02768_),
    .A2(_02769_),
    .ZN(_02770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07827_ (.A1(_01508_),
    .A2(_01269_),
    .A3(\mem[37][11] ),
    .ZN(_02771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07828_ (.A1(_01510_),
    .A2(\mem[38][11] ),
    .ZN(_02772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07829_ (.A1(_02771_),
    .A2(_02772_),
    .ZN(_02773_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07830_ (.A1(_02770_),
    .A2(_02773_),
    .ZN(_02774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07831_ (.A1(_01955_),
    .A2(_01264_),
    .A3(\mem[34][11] ),
    .ZN(_02775_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07832_ (.A1(_01957_),
    .A2(_01810_),
    .A3(\mem[33][11] ),
    .ZN(_02776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07833_ (.A1(_02775_),
    .A2(_02776_),
    .ZN(_02777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07834_ (.A1(_01286_),
    .A2(\mem[39][11] ),
    .ZN(_02778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07835_ (.A1(_01961_),
    .A2(_01450_),
    .A3(\mem[32][11] ),
    .ZN(_02779_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07836_ (.A1(_02778_),
    .A2(_02779_),
    .ZN(_02780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07837_ (.A1(_02777_),
    .A2(_02780_),
    .ZN(_02781_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07838_ (.A1(_02774_),
    .A2(_02781_),
    .ZN(_02782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07839_ (.A1(_02782_),
    .A2(_01127_),
    .ZN(_02783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07840_ (.A1(_01369_),
    .A2(_01523_),
    .A3(\mem[44][11] ),
    .ZN(_02784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07841_ (.A1(_01383_),
    .A2(_01820_),
    .A3(\mem[43][11] ),
    .ZN(_02785_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07842_ (.A1(_02784_),
    .A2(_02785_),
    .ZN(_02786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07843_ (.A1(_01435_),
    .A2(_01823_),
    .A3(\mem[45][11] ),
    .ZN(_02787_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07844_ (.A1(_01379_),
    .A2(\mem[46][11] ),
    .ZN(_02788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07845_ (.A1(_02787_),
    .A2(_02788_),
    .ZN(_02789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07846_ (.A1(_02786_),
    .A2(_02789_),
    .ZN(_02790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07847_ (.A1(_01974_),
    .A2(_01531_),
    .A3(\mem[42][11] ),
    .ZN(_02791_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07848_ (.A1(_01386_),
    .A2(_01829_),
    .A3(\mem[41][11] ),
    .ZN(_02792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07849_ (.A1(_02791_),
    .A2(_02792_),
    .ZN(_02793_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07850_ (.A1(_01535_),
    .A2(\mem[47][11] ),
    .ZN(_02794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07851_ (.A1(_01452_),
    .A2(_01537_),
    .A3(\mem[40][11] ),
    .ZN(_02795_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07852_ (.A1(_02794_),
    .A2(_02795_),
    .ZN(_02796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07853_ (.A1(_02793_),
    .A2(_02796_),
    .ZN(_02797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07854_ (.A1(_02790_),
    .A2(_02797_),
    .ZN(_02798_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07855_ (.A1(_02798_),
    .A2(_01149_),
    .ZN(_02799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07856_ (.A1(_02783_),
    .A2(_02799_),
    .ZN(_02800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07857_ (.A1(_01241_),
    .A2(_01384_),
    .A3(\mem[52][11] ),
    .ZN(_02801_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07858_ (.A1(_01415_),
    .A2(_01273_),
    .A3(\mem[51][11] ),
    .ZN(_02802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07859_ (.A1(_02801_),
    .A2(_02802_),
    .ZN(_02803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07860_ (.A1(_01547_),
    .A2(_01337_),
    .A3(\mem[53][11] ),
    .ZN(_02804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07861_ (.A1(_01411_),
    .A2(\mem[54][11] ),
    .ZN(_02805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07862_ (.A1(_02804_),
    .A2(_02805_),
    .ZN(_02806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07863_ (.A1(_02803_),
    .A2(_02806_),
    .ZN(_02807_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07864_ (.A1(_01992_),
    .A2(_01402_),
    .A3(\mem[50][11] ),
    .ZN(_02808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07865_ (.A1(_01254_),
    .A2(_01405_),
    .A3(\mem[49][11] ),
    .ZN(_02809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07866_ (.A1(_02808_),
    .A2(_02809_),
    .ZN(_02810_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07867_ (.A1(_01555_),
    .A2(\mem[55][11] ),
    .ZN(_02811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07868_ (.A1(_01997_),
    .A2(_01557_),
    .A3(\mem[48][11] ),
    .ZN(_02812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07869_ (.A1(_02811_),
    .A2(_02812_),
    .ZN(_02813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07870_ (.A1(_02810_),
    .A2(_02813_),
    .ZN(_02814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07871_ (.A1(_02807_),
    .A2(_02814_),
    .ZN(_02815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07872_ (.A1(_02815_),
    .A2(_01330_),
    .ZN(_02816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07873_ (.A1(_01563_),
    .A2(_01416_),
    .A3(\mem[60][11] ),
    .ZN(_02817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07874_ (.A1(_01449_),
    .A2(_01856_),
    .A3(\mem[59][11] ),
    .ZN(_02818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07875_ (.A1(_02817_),
    .A2(_02818_),
    .ZN(_02819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07876_ (.A1(_01442_),
    .A2(_01453_),
    .A3(\mem[61][11] ),
    .ZN(_02820_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07877_ (.A1(_01445_),
    .A2(\mem[62][11] ),
    .ZN(_02821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07878_ (.A1(_02820_),
    .A2(_02821_),
    .ZN(_02822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07879_ (.A1(_02819_),
    .A2(_02822_),
    .ZN(_02823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07880_ (.A1(_02010_),
    .A2(_01571_),
    .A3(\mem[58][11] ),
    .ZN(_02824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07881_ (.A1(_02012_),
    .A2(_01864_),
    .A3(\mem[57][11] ),
    .ZN(_02825_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07882_ (.A1(_02824_),
    .A2(_02825_),
    .ZN(_02826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07883_ (.A1(_01575_),
    .A2(\mem[63][11] ),
    .ZN(_02827_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07884_ (.A1(_01458_),
    .A2(_01577_),
    .A3(\mem[56][11] ),
    .ZN(_02828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07885_ (.A1(_02827_),
    .A2(_02828_),
    .ZN(_02829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07886_ (.A1(_02826_),
    .A2(_02829_),
    .ZN(_02830_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07887_ (.A1(_02823_),
    .A2(_02830_),
    .ZN(_02831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07888_ (.A1(_02831_),
    .A2(_01364_),
    .ZN(_02832_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07889_ (.A1(_02816_),
    .A2(_02832_),
    .ZN(_02833_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07890_ (.A1(_02800_),
    .A2(_02833_),
    .ZN(_02834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07891_ (.A1(_01585_),
    .A2(_01280_),
    .A3(\mem[4][11] ),
    .ZN(_02835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07892_ (.A1(_01312_),
    .A2(_01283_),
    .A3(\mem[3][11] ),
    .ZN(_02836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07893_ (.A1(_02835_),
    .A2(_02836_),
    .ZN(_02837_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07894_ (.A1(_01304_),
    .A2(_01878_),
    .A3(\mem[5][11] ),
    .ZN(_02838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07895_ (.A1(_01590_),
    .A2(\mem[6][11] ),
    .ZN(_02839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07896_ (.A1(_02838_),
    .A2(_02839_),
    .ZN(_02840_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07897_ (.A1(_02837_),
    .A2(_02840_),
    .ZN(_02841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07898_ (.A1(_02030_),
    .A2(_01594_),
    .A3(\mem[2][11] ),
    .ZN(_02842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07899_ (.A1(_02032_),
    .A2(_01377_),
    .A3(\mem[1][11] ),
    .ZN(_02843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07900_ (.A1(_02842_),
    .A2(_02843_),
    .ZN(_02844_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07901_ (.A1(_01320_),
    .A2(\mem[7][11] ),
    .ZN(_02845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07902_ (.A1(_01323_),
    .A2(_01324_),
    .A3(\mem[0][11] ),
    .ZN(_02846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07903_ (.A1(_02845_),
    .A2(_02846_),
    .ZN(_02847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07904_ (.A1(_02844_),
    .A2(_02847_),
    .ZN(_02848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07905_ (.A1(_02841_),
    .A2(_02848_),
    .ZN(_02849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07906_ (.A1(_02849_),
    .A2(_01398_),
    .ZN(_02850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07907_ (.A1(_01333_),
    .A2(_01604_),
    .A3(\mem[12][11] ),
    .ZN(_02851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07908_ (.A1(_01348_),
    .A2(_01893_),
    .A3(\mem[11][11] ),
    .ZN(_02852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07909_ (.A1(_02851_),
    .A2(_02852_),
    .ZN(_02853_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07910_ (.A1(_01608_),
    .A2(_01352_),
    .A3(\mem[13][11] ),
    .ZN(_02854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07911_ (.A1(_01610_),
    .A2(\mem[14][11] ),
    .ZN(_02855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07912_ (.A1(_02854_),
    .A2(_02855_),
    .ZN(_02856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07913_ (.A1(_02853_),
    .A2(_02856_),
    .ZN(_02857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07914_ (.A1(_02048_),
    .A2(_01614_),
    .A3(\mem[10][11] ),
    .ZN(_02858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07915_ (.A1(_01351_),
    .A2(_01439_),
    .A3(\mem[9][11] ),
    .ZN(_02859_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07916_ (.A1(_02858_),
    .A2(_02859_),
    .ZN(_02860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07917_ (.A1(_01355_),
    .A2(\mem[15][11] ),
    .ZN(_02861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07918_ (.A1(_02053_),
    .A2(_01359_),
    .A3(\mem[8][11] ),
    .ZN(_02862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07919_ (.A1(_02861_),
    .A2(_02862_),
    .ZN(_02863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07920_ (.A1(_02860_),
    .A2(_02863_),
    .ZN(_02864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07921_ (.A1(_02857_),
    .A2(_02864_),
    .ZN(_02865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07922_ (.A1(_02865_),
    .A2(_01431_),
    .ZN(_02866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07923_ (.A1(_02850_),
    .A2(_02866_),
    .ZN(_02867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07924_ (.A1(_01625_),
    .A2(_01349_),
    .A3(\mem[20][11] ),
    .ZN(_02868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07925_ (.A1(_01057_),
    .A2(_01911_),
    .A3(\mem[19][11] ),
    .ZN(_02869_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07926_ (.A1(_02868_),
    .A2(_02869_),
    .ZN(_02870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07927_ (.A1(_01629_),
    .A2(_01487_),
    .A3(\mem[21][11] ),
    .ZN(_02871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07928_ (.A1(_01631_),
    .A2(\mem[22][11] ),
    .ZN(_02872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07929_ (.A1(_02871_),
    .A2(_02872_),
    .ZN(_02873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07930_ (.A1(_02870_),
    .A2(_02873_),
    .ZN(_02874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07931_ (.A1(_02067_),
    .A2(_01635_),
    .A3(\mem[18][11] ),
    .ZN(_02875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07932_ (.A1(_02069_),
    .A2(_01919_),
    .A3(\mem[17][11] ),
    .ZN(_02876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07933_ (.A1(_02875_),
    .A2(_02876_),
    .ZN(_02877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07934_ (.A1(_01172_),
    .A2(\mem[23][11] ),
    .ZN(_02878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07935_ (.A1(_02073_),
    .A2(_01494_),
    .A3(\mem[16][11] ),
    .ZN(_02879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07936_ (.A1(_02878_),
    .A2(_02879_),
    .ZN(_02880_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07937_ (.A1(_02877_),
    .A2(_02880_),
    .ZN(_02881_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07938_ (.A1(_02874_),
    .A2(_02881_),
    .ZN(_02882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07939_ (.A1(_02882_),
    .A2(_01082_),
    .ZN(_02883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07940_ (.A1(_01408_),
    .A2(_01289_),
    .A3(\mem[28][11] ),
    .ZN(_02884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07941_ (.A1(_01483_),
    .A2(_01929_),
    .A3(_01782_),
    .A4(\mem[27][11] ),
    .ZN(_02885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07942_ (.A1(_02884_),
    .A2(_02885_),
    .ZN(_02886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07943_ (.A1(_01055_),
    .A2(_01044_),
    .A3(_01491_),
    .A4(\mem[29][11] ),
    .ZN(_02887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07944_ (.A1(_01649_),
    .A2(_01786_),
    .A3(_01047_),
    .A4(\mem[30][11] ),
    .ZN(_02888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07945_ (.A1(_02887_),
    .A2(_02888_),
    .ZN(_02889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07946_ (.A1(_02886_),
    .A2(_02889_),
    .ZN(_02890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07947_ (.A1(_01476_),
    .A2(_01790_),
    .A3(_01470_),
    .A4(\mem[26][11] ),
    .ZN(_02891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07948_ (.A1(_01424_),
    .A2(_01937_),
    .A3(\mem[25][11] ),
    .ZN(_02892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07949_ (.A1(_02891_),
    .A2(_02892_),
    .ZN(_02893_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07950_ (.A1(_01469_),
    .A2(_01477_),
    .A3(_02223_),
    .A4(\mem[31][11] ),
    .ZN(_02894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07951_ (.A1(_01049_),
    .A2(_01657_),
    .A3(\mem[24][11] ),
    .ZN(_02895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07952_ (.A1(_02894_),
    .A2(_02895_),
    .ZN(_02896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07953_ (.A1(_02893_),
    .A2(_02896_),
    .ZN(_02897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07954_ (.A1(_02890_),
    .A2(_02897_),
    .ZN(_02898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07955_ (.A1(_02898_),
    .A2(_01104_),
    .ZN(_02899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07956_ (.A1(_02883_),
    .A2(_02899_),
    .ZN(_02900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07957_ (.A1(_02867_),
    .A2(_02900_),
    .ZN(_02901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07958_ (.A1(_02834_),
    .A2(_02901_),
    .ZN(_00002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07959_ (.A1(_01263_),
    .A2(_01247_),
    .A3(\mem[36][12] ),
    .ZN(_02902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07960_ (.A1(_01279_),
    .A2(_01249_),
    .A3(\mem[35][12] ),
    .ZN(_02903_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07961_ (.A1(_02902_),
    .A2(_02903_),
    .ZN(_02904_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07962_ (.A1(_01401_),
    .A2(_01269_),
    .A3(\mem[37][12] ),
    .ZN(_02905_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07963_ (.A1(_01275_),
    .A2(\mem[38][12] ),
    .ZN(_02906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07964_ (.A1(_02905_),
    .A2(_02906_),
    .ZN(_02907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07965_ (.A1(_02904_),
    .A2(_02907_),
    .ZN(_02908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07966_ (.A1(_01955_),
    .A2(_01264_),
    .A3(\mem[34][12] ),
    .ZN(_02909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07967_ (.A1(_01957_),
    .A2(_01810_),
    .A3(\mem[33][12] ),
    .ZN(_02910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07968_ (.A1(_02909_),
    .A2(_02910_),
    .ZN(_02911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07969_ (.A1(_01286_),
    .A2(\mem[39][12] ),
    .ZN(_02912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07970_ (.A1(_01961_),
    .A2(_01450_),
    .A3(\mem[32][12] ),
    .ZN(_02913_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07971_ (.A1(_02912_),
    .A2(_02913_),
    .ZN(_02914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07972_ (.A1(_02911_),
    .A2(_02914_),
    .ZN(_02915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07973_ (.A1(_02908_),
    .A2(_02915_),
    .ZN(_02916_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07974_ (.A1(_02916_),
    .A2(_01127_),
    .ZN(_02917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07975_ (.A1(_01369_),
    .A2(_01370_),
    .A3(\mem[44][12] ),
    .ZN(_02918_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07976_ (.A1(_01383_),
    .A2(_01820_),
    .A3(\mem[43][12] ),
    .ZN(_02919_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07977_ (.A1(_02918_),
    .A2(_02919_),
    .ZN(_02920_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07978_ (.A1(_01435_),
    .A2(_01823_),
    .A3(\mem[45][12] ),
    .ZN(_02921_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07979_ (.A1(_01379_),
    .A2(\mem[46][12] ),
    .ZN(_02922_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07980_ (.A1(_02921_),
    .A2(_02922_),
    .ZN(_02923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07981_ (.A1(_02920_),
    .A2(_02923_),
    .ZN(_02924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07982_ (.A1(_01974_),
    .A2(_01298_),
    .A3(\mem[42][12] ),
    .ZN(_02925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07983_ (.A1(_01386_),
    .A2(_01829_),
    .A3(\mem[41][12] ),
    .ZN(_02926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07984_ (.A1(_02925_),
    .A2(_02926_),
    .ZN(_02927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07985_ (.A1(_01390_),
    .A2(\mem[47][12] ),
    .ZN(_02928_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07986_ (.A1(_01452_),
    .A2(_01393_),
    .A3(\mem[40][12] ),
    .ZN(_02929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07987_ (.A1(_02928_),
    .A2(_02929_),
    .ZN(_02930_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07988_ (.A1(_02927_),
    .A2(_02930_),
    .ZN(_02931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07989_ (.A1(_02924_),
    .A2(_02931_),
    .ZN(_02932_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07990_ (.A1(_02932_),
    .A2(_01149_),
    .ZN(_02933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07991_ (.A1(_02917_),
    .A2(_02933_),
    .ZN(_02934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07992_ (.A1(_01241_),
    .A2(_01384_),
    .A3(\mem[52][12] ),
    .ZN(_02935_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07993_ (.A1(_01415_),
    .A2(_01273_),
    .A3(\mem[51][12] ),
    .ZN(_02936_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07994_ (.A1(_02935_),
    .A2(_02936_),
    .ZN(_02937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07995_ (.A1(_01466_),
    .A2(_01337_),
    .A3(\mem[53][12] ),
    .ZN(_02938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07996_ (.A1(_01411_),
    .A2(\mem[54][12] ),
    .ZN(_02939_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07997_ (.A1(_02938_),
    .A2(_02939_),
    .ZN(_02940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07998_ (.A1(_02937_),
    .A2(_02940_),
    .ZN(_02941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07999_ (.A1(_01992_),
    .A2(_01402_),
    .A3(\mem[50][12] ),
    .ZN(_02942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08000_ (.A1(_01254_),
    .A2(_01405_),
    .A3(\mem[49][12] ),
    .ZN(_02943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08001_ (.A1(_02942_),
    .A2(_02943_),
    .ZN(_02944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08002_ (.A1(_01422_),
    .A2(\mem[55][12] ),
    .ZN(_02945_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08003_ (.A1(_01997_),
    .A2(_01425_),
    .A3(\mem[48][12] ),
    .ZN(_02946_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08004_ (.A1(_02945_),
    .A2(_02946_),
    .ZN(_02947_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08005_ (.A1(_02944_),
    .A2(_02947_),
    .ZN(_02948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08006_ (.A1(_02941_),
    .A2(_02948_),
    .ZN(_02949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08007_ (.A1(_02949_),
    .A2(_01330_),
    .ZN(_02950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08008_ (.A1(_01272_),
    .A2(_01416_),
    .A3(\mem[60][12] ),
    .ZN(_02951_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08009_ (.A1(_01449_),
    .A2(_01856_),
    .A3(\mem[59][12] ),
    .ZN(_02952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08010_ (.A1(_02951_),
    .A2(_02952_),
    .ZN(_02953_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08011_ (.A1(_01442_),
    .A2(_01453_),
    .A3(\mem[61][12] ),
    .ZN(_02954_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08012_ (.A1(_01445_),
    .A2(\mem[62][12] ),
    .ZN(_02955_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08013_ (.A1(_02954_),
    .A2(_02955_),
    .ZN(_02956_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08014_ (.A1(_02953_),
    .A2(_02956_),
    .ZN(_02957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08015_ (.A1(_02010_),
    .A2(_01256_),
    .A3(\mem[58][12] ),
    .ZN(_02958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08016_ (.A1(_02012_),
    .A2(_01864_),
    .A3(\mem[57][12] ),
    .ZN(_02959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08017_ (.A1(_02958_),
    .A2(_02959_),
    .ZN(_02960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08018_ (.A1(_01456_),
    .A2(\mem[63][12] ),
    .ZN(_02961_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08019_ (.A1(_01458_),
    .A2(_01459_),
    .A3(\mem[56][12] ),
    .ZN(_02962_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08020_ (.A1(_02961_),
    .A2(_02962_),
    .ZN(_02963_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08021_ (.A1(_02960_),
    .A2(_02963_),
    .ZN(_02964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08022_ (.A1(_02957_),
    .A2(_02964_),
    .ZN(_02965_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08023_ (.A1(_02965_),
    .A2(_01364_),
    .ZN(_02966_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08024_ (.A1(_02950_),
    .A2(_02966_),
    .ZN(_02967_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08025_ (.A1(_02934_),
    .A2(_02967_),
    .ZN(_02968_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08026_ (.A1(_01297_),
    .A2(_01280_),
    .A3(\mem[4][12] ),
    .ZN(_02969_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08027_ (.A1(_01312_),
    .A2(_01283_),
    .A3(\mem[3][12] ),
    .ZN(_02970_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08028_ (.A1(_02969_),
    .A2(_02970_),
    .ZN(_02971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08029_ (.A1(_01304_),
    .A2(_01878_),
    .A3(\mem[5][12] ),
    .ZN(_02972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08030_ (.A1(_01308_),
    .A2(\mem[6][12] ),
    .ZN(_02973_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08031_ (.A1(_02972_),
    .A2(_02973_),
    .ZN(_02974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08032_ (.A1(_02971_),
    .A2(_02974_),
    .ZN(_02975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08033_ (.A1(_02030_),
    .A2(_01314_),
    .A3(\mem[2][12] ),
    .ZN(_02976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08034_ (.A1(_02032_),
    .A2(_01377_),
    .A3(\mem[1][12] ),
    .ZN(_02977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08035_ (.A1(_02976_),
    .A2(_02977_),
    .ZN(_02978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08036_ (.A1(_01320_),
    .A2(\mem[7][12] ),
    .ZN(_02979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08037_ (.A1(_01323_),
    .A2(_01324_),
    .A3(\mem[0][12] ),
    .ZN(_02980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08038_ (.A1(_02979_),
    .A2(_02980_),
    .ZN(_02981_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08039_ (.A1(_02978_),
    .A2(_02981_),
    .ZN(_02982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08040_ (.A1(_02975_),
    .A2(_02982_),
    .ZN(_02983_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08041_ (.A1(_02983_),
    .A2(_01398_),
    .ZN(_02984_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08042_ (.A1(_01333_),
    .A2(_01334_),
    .A3(\mem[12][12] ),
    .ZN(_02985_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08043_ (.A1(_01348_),
    .A2(_01893_),
    .A3(\mem[11][12] ),
    .ZN(_02986_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08044_ (.A1(_02985_),
    .A2(_02986_),
    .ZN(_02987_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08045_ (.A1(_01340_),
    .A2(_01352_),
    .A3(\mem[13][12] ),
    .ZN(_02988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08046_ (.A1(_01344_),
    .A2(\mem[14][12] ),
    .ZN(_02989_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08047_ (.A1(_02988_),
    .A2(_02989_),
    .ZN(_02990_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08048_ (.A1(_02987_),
    .A2(_02990_),
    .ZN(_02991_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08049_ (.A1(_02048_),
    .A2(_01436_),
    .A3(\mem[10][12] ),
    .ZN(_02992_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08050_ (.A1(_01351_),
    .A2(_01439_),
    .A3(\mem[9][12] ),
    .ZN(_02993_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08051_ (.A1(_02992_),
    .A2(_02993_),
    .ZN(_02994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08052_ (.A1(_01355_),
    .A2(\mem[15][12] ),
    .ZN(_02995_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08053_ (.A1(_02053_),
    .A2(_01359_),
    .A3(\mem[8][12] ),
    .ZN(_02996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08054_ (.A1(_02995_),
    .A2(_02996_),
    .ZN(_02997_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08055_ (.A1(_02994_),
    .A2(_02997_),
    .ZN(_02998_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08056_ (.A1(_02991_),
    .A2(_02998_),
    .ZN(_02999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08057_ (.A1(_02999_),
    .A2(_01431_),
    .ZN(_03000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08058_ (.A1(_02984_),
    .A2(_03000_),
    .ZN(_03001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08059_ (.A1(_01376_),
    .A2(_01349_),
    .A3(\mem[20][12] ),
    .ZN(_03002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08060_ (.A1(_01057_),
    .A2(_01911_),
    .A3(\mem[19][12] ),
    .ZN(_03003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08061_ (.A1(_03002_),
    .A2(_03003_),
    .ZN(_03004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08062_ (.A1(_01067_),
    .A2(_01487_),
    .A3(\mem[21][12] ),
    .ZN(_03005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08063_ (.A1(_01161_),
    .A2(\mem[22][12] ),
    .ZN(_03006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08064_ (.A1(_03005_),
    .A2(_03006_),
    .ZN(_03007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08065_ (.A1(_03004_),
    .A2(_03007_),
    .ZN(_03008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08066_ (.A1(_02067_),
    .A2(_01467_),
    .A3(\mem[18][12] ),
    .ZN(_03009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08067_ (.A1(_02069_),
    .A2(_01919_),
    .A3(\mem[17][12] ),
    .ZN(_03010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08068_ (.A1(_03009_),
    .A2(_03010_),
    .ZN(_03011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08069_ (.A1(_01172_),
    .A2(\mem[23][12] ),
    .ZN(_03012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08070_ (.A1(_02073_),
    .A2(_01494_),
    .A3(\mem[16][12] ),
    .ZN(_03013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08071_ (.A1(_03012_),
    .A2(_03013_),
    .ZN(_03014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08072_ (.A1(_03011_),
    .A2(_03014_),
    .ZN(_03015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08073_ (.A1(_03008_),
    .A2(_03015_),
    .ZN(_03016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08074_ (.A1(_03016_),
    .A2(_01082_),
    .ZN(_03017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08075_ (.A1(_01408_),
    .A2(_01289_),
    .A3(\mem[28][12] ),
    .ZN(_03018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08076_ (.A1(_01483_),
    .A2(_01929_),
    .A3(_01782_),
    .A4(\mem[27][12] ),
    .ZN(_03019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08077_ (.A1(_03018_),
    .A2(_03019_),
    .ZN(_03020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08078_ (.A1(_01055_),
    .A2(_01044_),
    .A3(_01491_),
    .A4(\mem[29][12] ),
    .ZN(_03021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08079_ (.A1(_01041_),
    .A2(_01786_),
    .A3(_01047_),
    .A4(\mem[30][12] ),
    .ZN(_03022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08080_ (.A1(_03021_),
    .A2(_03022_),
    .ZN(_03023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08081_ (.A1(_03020_),
    .A2(_03023_),
    .ZN(_03024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08082_ (.A1(_01476_),
    .A2(_01790_),
    .A3(_01470_),
    .A4(\mem[26][12] ),
    .ZN(_03025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08083_ (.A1(_01424_),
    .A2(_01937_),
    .A3(\mem[25][12] ),
    .ZN(_03026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08084_ (.A1(_03025_),
    .A2(_03026_),
    .ZN(_03027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08085_ (.A1(_01469_),
    .A2(_01477_),
    .A3(_02223_),
    .A4(\mem[31][12] ),
    .ZN(_03028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08086_ (.A1(_01049_),
    .A2(_01482_),
    .A3(\mem[24][12] ),
    .ZN(_03029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08087_ (.A1(_03028_),
    .A2(_03029_),
    .ZN(_03030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08088_ (.A1(_03027_),
    .A2(_03030_),
    .ZN(_03031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08089_ (.A1(_03024_),
    .A2(_03031_),
    .ZN(_03032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08090_ (.A1(_03032_),
    .A2(_01104_),
    .ZN(_03033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08091_ (.A1(_03017_),
    .A2(_03033_),
    .ZN(_03034_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08092_ (.A1(_03001_),
    .A2(_03034_),
    .ZN(_03035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08093_ (.A1(_02968_),
    .A2(_03035_),
    .ZN(_00003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08094_ (.A1(_01263_),
    .A2(_01247_),
    .A3(\mem[36][13] ),
    .ZN(_03036_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08095_ (.A1(_01279_),
    .A2(_01249_),
    .A3(\mem[35][13] ),
    .ZN(_03037_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08096_ (.A1(_03036_),
    .A2(_03037_),
    .ZN(_03038_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08097_ (.A1(_01401_),
    .A2(_01269_),
    .A3(\mem[37][13] ),
    .ZN(_03039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08098_ (.A1(_01275_),
    .A2(\mem[38][13] ),
    .ZN(_03040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08099_ (.A1(_03039_),
    .A2(_03040_),
    .ZN(_03041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08100_ (.A1(_03038_),
    .A2(_03041_),
    .ZN(_03042_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08101_ (.A1(_01955_),
    .A2(_01264_),
    .A3(\mem[34][13] ),
    .ZN(_03043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08102_ (.A1(_01957_),
    .A2(_01810_),
    .A3(\mem[33][13] ),
    .ZN(_03044_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08103_ (.A1(_03043_),
    .A2(_03044_),
    .ZN(_03045_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08104_ (.A1(_01286_),
    .A2(\mem[39][13] ),
    .ZN(_03046_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08105_ (.A1(_01961_),
    .A2(_01450_),
    .A3(\mem[32][13] ),
    .ZN(_03047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08106_ (.A1(_03046_),
    .A2(_03047_),
    .ZN(_03048_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08107_ (.A1(_03045_),
    .A2(_03048_),
    .ZN(_03049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08108_ (.A1(_03042_),
    .A2(_03049_),
    .ZN(_03050_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08109_ (.A1(_03050_),
    .A2(_01127_),
    .ZN(_03051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08110_ (.A1(_01369_),
    .A2(_01370_),
    .A3(\mem[44][13] ),
    .ZN(_03052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08111_ (.A1(_01383_),
    .A2(_01820_),
    .A3(\mem[43][13] ),
    .ZN(_03053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08112_ (.A1(_03052_),
    .A2(_03053_),
    .ZN(_03054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08113_ (.A1(_01435_),
    .A2(_01823_),
    .A3(\mem[45][13] ),
    .ZN(_03055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08114_ (.A1(_01379_),
    .A2(\mem[46][13] ),
    .ZN(_03056_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08115_ (.A1(_03055_),
    .A2(_03056_),
    .ZN(_03057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08116_ (.A1(_03054_),
    .A2(_03057_),
    .ZN(_03058_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08117_ (.A1(_01974_),
    .A2(_01298_),
    .A3(\mem[42][13] ),
    .ZN(_03059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08118_ (.A1(_01386_),
    .A2(_01829_),
    .A3(\mem[41][13] ),
    .ZN(_03060_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08119_ (.A1(_03059_),
    .A2(_03060_),
    .ZN(_03061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08120_ (.A1(_01390_),
    .A2(\mem[47][13] ),
    .ZN(_03062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08121_ (.A1(_01452_),
    .A2(_01393_),
    .A3(\mem[40][13] ),
    .ZN(_03063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08122_ (.A1(_03062_),
    .A2(_03063_),
    .ZN(_03064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08123_ (.A1(_03061_),
    .A2(_03064_),
    .ZN(_03065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08124_ (.A1(_03058_),
    .A2(_03065_),
    .ZN(_03066_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08125_ (.A1(_03066_),
    .A2(_01149_),
    .ZN(_03067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08126_ (.A1(_03051_),
    .A2(_03067_),
    .ZN(_03068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08127_ (.A1(_01241_),
    .A2(_01384_),
    .A3(\mem[52][13] ),
    .ZN(_03069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08128_ (.A1(_01415_),
    .A2(_01273_),
    .A3(\mem[51][13] ),
    .ZN(_03070_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08129_ (.A1(_03069_),
    .A2(_03070_),
    .ZN(_03071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08130_ (.A1(_01466_),
    .A2(_01337_),
    .A3(\mem[53][13] ),
    .ZN(_03072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08131_ (.A1(_01411_),
    .A2(\mem[54][13] ),
    .ZN(_03073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08132_ (.A1(_03072_),
    .A2(_03073_),
    .ZN(_03074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08133_ (.A1(_03071_),
    .A2(_03074_),
    .ZN(_03075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08134_ (.A1(_01992_),
    .A2(_01402_),
    .A3(\mem[50][13] ),
    .ZN(_03076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08135_ (.A1(_01254_),
    .A2(_01405_),
    .A3(\mem[49][13] ),
    .ZN(_03077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08136_ (.A1(_03076_),
    .A2(_03077_),
    .ZN(_03078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08137_ (.A1(_01422_),
    .A2(\mem[55][13] ),
    .ZN(_03079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08138_ (.A1(_01997_),
    .A2(_01425_),
    .A3(\mem[48][13] ),
    .ZN(_03080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08139_ (.A1(_03079_),
    .A2(_03080_),
    .ZN(_03081_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08140_ (.A1(_03078_),
    .A2(_03081_),
    .ZN(_03082_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08141_ (.A1(_03075_),
    .A2(_03082_),
    .ZN(_03083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08142_ (.A1(_03083_),
    .A2(_01330_),
    .ZN(_03084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08143_ (.A1(_01272_),
    .A2(_01416_),
    .A3(\mem[60][13] ),
    .ZN(_03085_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08144_ (.A1(_01449_),
    .A2(_01856_),
    .A3(\mem[59][13] ),
    .ZN(_03086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08145_ (.A1(_03085_),
    .A2(_03086_),
    .ZN(_03087_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08146_ (.A1(_01442_),
    .A2(_01453_),
    .A3(\mem[61][13] ),
    .ZN(_03088_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08147_ (.A1(_01445_),
    .A2(\mem[62][13] ),
    .ZN(_03089_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08148_ (.A1(_03088_),
    .A2(_03089_),
    .ZN(_03090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08149_ (.A1(_03087_),
    .A2(_03090_),
    .ZN(_03091_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08150_ (.A1(_02010_),
    .A2(_01256_),
    .A3(\mem[58][13] ),
    .ZN(_03092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08151_ (.A1(_02012_),
    .A2(_01864_),
    .A3(\mem[57][13] ),
    .ZN(_03093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08152_ (.A1(_03092_),
    .A2(_03093_),
    .ZN(_03094_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08153_ (.A1(_01456_),
    .A2(\mem[63][13] ),
    .ZN(_03095_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08154_ (.A1(_01458_),
    .A2(_01459_),
    .A3(\mem[56][13] ),
    .ZN(_03096_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08155_ (.A1(_03095_),
    .A2(_03096_),
    .ZN(_03097_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08156_ (.A1(_03094_),
    .A2(_03097_),
    .ZN(_03098_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08157_ (.A1(_03091_),
    .A2(_03098_),
    .ZN(_03099_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08158_ (.A1(_03099_),
    .A2(_01364_),
    .ZN(_03100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08159_ (.A1(_03084_),
    .A2(_03100_),
    .ZN(_03101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08160_ (.A1(_03068_),
    .A2(_03101_),
    .ZN(_03102_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08161_ (.A1(_01297_),
    .A2(_01280_),
    .A3(\mem[4][13] ),
    .ZN(_03103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08162_ (.A1(_01312_),
    .A2(_01283_),
    .A3(\mem[3][13] ),
    .ZN(_03104_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08163_ (.A1(_03103_),
    .A2(_03104_),
    .ZN(_03105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08164_ (.A1(_01304_),
    .A2(_01878_),
    .A3(\mem[5][13] ),
    .ZN(_03106_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08165_ (.A1(_01308_),
    .A2(\mem[6][13] ),
    .ZN(_03107_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08166_ (.A1(_03106_),
    .A2(_03107_),
    .ZN(_03108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08167_ (.A1(_03105_),
    .A2(_03108_),
    .ZN(_03109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08168_ (.A1(_02030_),
    .A2(_01314_),
    .A3(\mem[2][13] ),
    .ZN(_03110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08169_ (.A1(_02032_),
    .A2(_01377_),
    .A3(\mem[1][13] ),
    .ZN(_03111_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08170_ (.A1(_03110_),
    .A2(_03111_),
    .ZN(_03112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08171_ (.A1(_01320_),
    .A2(\mem[7][13] ),
    .ZN(_03113_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08172_ (.A1(_01323_),
    .A2(_01324_),
    .A3(\mem[0][13] ),
    .ZN(_03114_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08173_ (.A1(_03113_),
    .A2(_03114_),
    .ZN(_03115_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08174_ (.A1(_03112_),
    .A2(_03115_),
    .ZN(_03116_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08175_ (.A1(_03109_),
    .A2(_03116_),
    .ZN(_03117_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08176_ (.A1(_03117_),
    .A2(_01398_),
    .ZN(_03118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08177_ (.A1(_01333_),
    .A2(_01334_),
    .A3(\mem[12][13] ),
    .ZN(_03119_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08178_ (.A1(_01348_),
    .A2(_01893_),
    .A3(\mem[11][13] ),
    .ZN(_03120_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08179_ (.A1(_03119_),
    .A2(_03120_),
    .ZN(_03121_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08180_ (.A1(_01340_),
    .A2(_01352_),
    .A3(\mem[13][13] ),
    .ZN(_03122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08181_ (.A1(_01344_),
    .A2(\mem[14][13] ),
    .ZN(_03123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08182_ (.A1(_03122_),
    .A2(_03123_),
    .ZN(_03124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08183_ (.A1(_03121_),
    .A2(_03124_),
    .ZN(_03125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08184_ (.A1(_02048_),
    .A2(_01436_),
    .A3(\mem[10][13] ),
    .ZN(_03126_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08185_ (.A1(_01351_),
    .A2(_01439_),
    .A3(\mem[9][13] ),
    .ZN(_03127_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08186_ (.A1(_03126_),
    .A2(_03127_),
    .ZN(_03128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08187_ (.A1(_01355_),
    .A2(\mem[15][13] ),
    .ZN(_03129_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08188_ (.A1(_02053_),
    .A2(_01359_),
    .A3(\mem[8][13] ),
    .ZN(_03130_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08189_ (.A1(_03129_),
    .A2(_03130_),
    .ZN(_03131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08190_ (.A1(_03128_),
    .A2(_03131_),
    .ZN(_03132_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08191_ (.A1(_03125_),
    .A2(_03132_),
    .ZN(_03133_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08192_ (.A1(_03133_),
    .A2(_01431_),
    .ZN(_03134_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08193_ (.A1(_03118_),
    .A2(_03134_),
    .ZN(_03135_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08194_ (.A1(_01376_),
    .A2(_01349_),
    .A3(\mem[20][13] ),
    .ZN(_03136_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08195_ (.A1(_01057_),
    .A2(_01911_),
    .A3(\mem[19][13] ),
    .ZN(_03137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08196_ (.A1(_03136_),
    .A2(_03137_),
    .ZN(_03138_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08197_ (.A1(_01067_),
    .A2(_01487_),
    .A3(\mem[21][13] ),
    .ZN(_03139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08198_ (.A1(_01161_),
    .A2(\mem[22][13] ),
    .ZN(_03140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08199_ (.A1(_03139_),
    .A2(_03140_),
    .ZN(_03141_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08200_ (.A1(_03138_),
    .A2(_03141_),
    .ZN(_03142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08201_ (.A1(_02067_),
    .A2(_01467_),
    .A3(\mem[18][13] ),
    .ZN(_03143_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08202_ (.A1(_02069_),
    .A2(_01919_),
    .A3(\mem[17][13] ),
    .ZN(_03144_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08203_ (.A1(_03143_),
    .A2(_03144_),
    .ZN(_03145_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08204_ (.A1(_01172_),
    .A2(\mem[23][13] ),
    .ZN(_03146_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08205_ (.A1(_02073_),
    .A2(_01494_),
    .A3(\mem[16][13] ),
    .ZN(_03147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08206_ (.A1(_03146_),
    .A2(_03147_),
    .ZN(_03148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08207_ (.A1(_03145_),
    .A2(_03148_),
    .ZN(_03149_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08208_ (.A1(_03142_),
    .A2(_03149_),
    .ZN(_03150_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08209_ (.A1(_03150_),
    .A2(_01082_),
    .ZN(_03151_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08210_ (.A1(_01408_),
    .A2(_01289_),
    .A3(\mem[28][13] ),
    .ZN(_03152_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08211_ (.A1(_01483_),
    .A2(_01929_),
    .A3(_01153_),
    .A4(\mem[27][13] ),
    .ZN(_03153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08212_ (.A1(_03152_),
    .A2(_03153_),
    .ZN(_03154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08213_ (.A1(_01055_),
    .A2(_01044_),
    .A3(_01491_),
    .A4(\mem[29][13] ),
    .ZN(_03155_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08214_ (.A1(_01041_),
    .A2(_01484_),
    .A3(_01047_),
    .A4(\mem[30][13] ),
    .ZN(_03156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08215_ (.A1(_03155_),
    .A2(_03156_),
    .ZN(_03157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08216_ (.A1(_03154_),
    .A2(_03157_),
    .ZN(_03158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08217_ (.A1(_01476_),
    .A2(_01065_),
    .A3(_01470_),
    .A4(\mem[26][13] ),
    .ZN(_03159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08218_ (.A1(_01424_),
    .A2(_01937_),
    .A3(\mem[25][13] ),
    .ZN(_03160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08219_ (.A1(_03159_),
    .A2(_03160_),
    .ZN(_03161_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08220_ (.A1(_01469_),
    .A2(_01477_),
    .A3(_02223_),
    .A4(\mem[31][13] ),
    .ZN(_03162_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08221_ (.A1(_01049_),
    .A2(_01482_),
    .A3(\mem[24][13] ),
    .ZN(_03163_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08222_ (.A1(_03162_),
    .A2(_03163_),
    .ZN(_03164_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08223_ (.A1(_03161_),
    .A2(_03164_),
    .ZN(_03165_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08224_ (.A1(_03158_),
    .A2(_03165_),
    .ZN(_03166_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08225_ (.A1(_03166_),
    .A2(_01104_),
    .ZN(_03167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08226_ (.A1(_03151_),
    .A2(_03167_),
    .ZN(_03168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08227_ (.A1(_03135_),
    .A2(_03168_),
    .ZN(_03169_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08228_ (.A1(_03102_),
    .A2(_03169_),
    .ZN(_00004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08229_ (.A1(_01263_),
    .A2(_01247_),
    .A3(\mem[36][14] ),
    .ZN(_03170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08230_ (.A1(_01279_),
    .A2(_01249_),
    .A3(\mem[35][14] ),
    .ZN(_03171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08231_ (.A1(_03170_),
    .A2(_03171_),
    .ZN(_03172_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08232_ (.A1(_01401_),
    .A2(_01269_),
    .A3(\mem[37][14] ),
    .ZN(_03173_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08233_ (.A1(_01275_),
    .A2(\mem[38][14] ),
    .ZN(_03174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08234_ (.A1(_03173_),
    .A2(_03174_),
    .ZN(_03175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08235_ (.A1(_03172_),
    .A2(_03175_),
    .ZN(_03176_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08236_ (.A1(_01955_),
    .A2(_01264_),
    .A3(\mem[34][14] ),
    .ZN(_03177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08237_ (.A1(_01957_),
    .A2(_01242_),
    .A3(\mem[33][14] ),
    .ZN(_03178_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08238_ (.A1(_03177_),
    .A2(_03178_),
    .ZN(_03179_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08239_ (.A1(_01286_),
    .A2(\mem[39][14] ),
    .ZN(_03180_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08240_ (.A1(_01961_),
    .A2(_01450_),
    .A3(\mem[32][14] ),
    .ZN(_03181_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08241_ (.A1(_03180_),
    .A2(_03181_),
    .ZN(_03182_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08242_ (.A1(_03179_),
    .A2(_03182_),
    .ZN(_03183_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08243_ (.A1(_03176_),
    .A2(_03183_),
    .ZN(_03184_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08244_ (.A1(_03184_),
    .A2(_01127_),
    .ZN(_03185_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08245_ (.A1(_01369_),
    .A2(_01370_),
    .A3(\mem[44][14] ),
    .ZN(_03186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08246_ (.A1(_01383_),
    .A2(_01373_),
    .A3(\mem[43][14] ),
    .ZN(_03187_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08247_ (.A1(_03186_),
    .A2(_03187_),
    .ZN(_03188_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08248_ (.A1(_01435_),
    .A2(_01387_),
    .A3(\mem[45][14] ),
    .ZN(_03189_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08249_ (.A1(_01379_),
    .A2(\mem[46][14] ),
    .ZN(_03190_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08250_ (.A1(_03189_),
    .A2(_03190_),
    .ZN(_03191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08251_ (.A1(_03188_),
    .A2(_03191_),
    .ZN(_03192_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08252_ (.A1(_01974_),
    .A2(_01298_),
    .A3(\mem[42][14] ),
    .ZN(_03193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08253_ (.A1(_01386_),
    .A2(_01301_),
    .A3(\mem[41][14] ),
    .ZN(_03194_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08254_ (.A1(_03193_),
    .A2(_03194_),
    .ZN(_03195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08255_ (.A1(_01390_),
    .A2(\mem[47][14] ),
    .ZN(_03196_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08256_ (.A1(_01452_),
    .A2(_01393_),
    .A3(\mem[40][14] ),
    .ZN(_03197_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08257_ (.A1(_03196_),
    .A2(_03197_),
    .ZN(_03198_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08258_ (.A1(_03195_),
    .A2(_03198_),
    .ZN(_03199_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08259_ (.A1(_03192_),
    .A2(_03199_),
    .ZN(_03200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08260_ (.A1(_03200_),
    .A2(_01149_),
    .ZN(_03201_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08261_ (.A1(_03185_),
    .A2(_03201_),
    .ZN(_03202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08262_ (.A1(_01241_),
    .A2(_01384_),
    .A3(\mem[52][14] ),
    .ZN(_03203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08263_ (.A1(_01415_),
    .A2(_01273_),
    .A3(\mem[51][14] ),
    .ZN(_03204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08264_ (.A1(_03203_),
    .A2(_03204_),
    .ZN(_03205_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08265_ (.A1(_01466_),
    .A2(_01337_),
    .A3(\mem[53][14] ),
    .ZN(_03206_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08266_ (.A1(_01411_),
    .A2(\mem[54][14] ),
    .ZN(_03207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08267_ (.A1(_03206_),
    .A2(_03207_),
    .ZN(_03208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08268_ (.A1(_03205_),
    .A2(_03208_),
    .ZN(_03209_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08269_ (.A1(_01992_),
    .A2(_01402_),
    .A3(\mem[50][14] ),
    .ZN(_03210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08270_ (.A1(_01254_),
    .A2(_01405_),
    .A3(\mem[49][14] ),
    .ZN(_03211_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08271_ (.A1(_03210_),
    .A2(_03211_),
    .ZN(_03212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08272_ (.A1(_01422_),
    .A2(\mem[55][14] ),
    .ZN(_03213_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08273_ (.A1(_01997_),
    .A2(_01425_),
    .A3(\mem[48][14] ),
    .ZN(_03214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08274_ (.A1(_03213_),
    .A2(_03214_),
    .ZN(_03215_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08275_ (.A1(_03212_),
    .A2(_03215_),
    .ZN(_03216_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08276_ (.A1(_03209_),
    .A2(_03216_),
    .ZN(_03217_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08277_ (.A1(_03217_),
    .A2(_01330_),
    .ZN(_03218_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08278_ (.A1(_01272_),
    .A2(_01416_),
    .A3(\mem[60][14] ),
    .ZN(_03219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08279_ (.A1(_01449_),
    .A2(_01419_),
    .A3(\mem[59][14] ),
    .ZN(_03220_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08280_ (.A1(_03219_),
    .A2(_03220_),
    .ZN(_03221_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08281_ (.A1(_01442_),
    .A2(_01453_),
    .A3(\mem[61][14] ),
    .ZN(_03222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08282_ (.A1(_01445_),
    .A2(\mem[62][14] ),
    .ZN(_03223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08283_ (.A1(_03222_),
    .A2(_03223_),
    .ZN(_03224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08284_ (.A1(_03221_),
    .A2(_03224_),
    .ZN(_03225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08285_ (.A1(_02010_),
    .A2(_01256_),
    .A3(\mem[58][14] ),
    .ZN(_03226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08286_ (.A1(_02012_),
    .A2(_01342_),
    .A3(\mem[57][14] ),
    .ZN(_03227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08287_ (.A1(_03226_),
    .A2(_03227_),
    .ZN(_03228_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08288_ (.A1(_01456_),
    .A2(\mem[63][14] ),
    .ZN(_03229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08289_ (.A1(_01458_),
    .A2(_01459_),
    .A3(\mem[56][14] ),
    .ZN(_03230_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08290_ (.A1(_03229_),
    .A2(_03230_),
    .ZN(_03231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08291_ (.A1(_03228_),
    .A2(_03231_),
    .ZN(_03232_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08292_ (.A1(_03225_),
    .A2(_03232_),
    .ZN(_03233_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08293_ (.A1(_03233_),
    .A2(_01364_),
    .ZN(_03234_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08294_ (.A1(_03218_),
    .A2(_03234_),
    .ZN(_03235_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08295_ (.A1(_03202_),
    .A2(_03235_),
    .ZN(_03236_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08296_ (.A1(_01297_),
    .A2(_01280_),
    .A3(\mem[4][14] ),
    .ZN(_03237_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08297_ (.A1(_01312_),
    .A2(_01283_),
    .A3(\mem[3][14] ),
    .ZN(_03238_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08298_ (.A1(_03237_),
    .A2(_03238_),
    .ZN(_03239_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08299_ (.A1(_01304_),
    .A2(_01317_),
    .A3(\mem[5][14] ),
    .ZN(_03240_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08300_ (.A1(_01308_),
    .A2(\mem[6][14] ),
    .ZN(_03241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08301_ (.A1(_03240_),
    .A2(_03241_),
    .ZN(_03242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08302_ (.A1(_03239_),
    .A2(_03242_),
    .ZN(_03243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08303_ (.A1(_02030_),
    .A2(_01314_),
    .A3(\mem[2][14] ),
    .ZN(_03244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08304_ (.A1(_02032_),
    .A2(_01377_),
    .A3(\mem[1][14] ),
    .ZN(_03245_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08305_ (.A1(_03244_),
    .A2(_03245_),
    .ZN(_03246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08306_ (.A1(_01320_),
    .A2(\mem[7][14] ),
    .ZN(_03247_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08307_ (.A1(_01323_),
    .A2(_01324_),
    .A3(\mem[0][14] ),
    .ZN(_03248_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08308_ (.A1(_03247_),
    .A2(_03248_),
    .ZN(_03249_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08309_ (.A1(_03246_),
    .A2(_03249_),
    .ZN(_03250_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08310_ (.A1(_03243_),
    .A2(_03250_),
    .ZN(_03251_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08311_ (.A1(_03251_),
    .A2(_01398_),
    .ZN(_03252_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08312_ (.A1(_01333_),
    .A2(_01334_),
    .A3(\mem[12][14] ),
    .ZN(_03253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08313_ (.A1(_01348_),
    .A2(_01306_),
    .A3(\mem[11][14] ),
    .ZN(_03254_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08314_ (.A1(_03253_),
    .A2(_03254_),
    .ZN(_03255_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08315_ (.A1(_01340_),
    .A2(_01352_),
    .A3(\mem[13][14] ),
    .ZN(_03256_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08316_ (.A1(_01344_),
    .A2(\mem[14][14] ),
    .ZN(_03257_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08317_ (.A1(_03256_),
    .A2(_03257_),
    .ZN(_03258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08318_ (.A1(_03255_),
    .A2(_03258_),
    .ZN(_03259_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08319_ (.A1(_02048_),
    .A2(_01436_),
    .A3(\mem[10][14] ),
    .ZN(_03260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08320_ (.A1(_01351_),
    .A2(_01439_),
    .A3(\mem[9][14] ),
    .ZN(_03261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08321_ (.A1(_03260_),
    .A2(_03261_),
    .ZN(_03262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08322_ (.A1(_01355_),
    .A2(\mem[15][14] ),
    .ZN(_03263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08323_ (.A1(_02053_),
    .A2(_01359_),
    .A3(\mem[8][14] ),
    .ZN(_03264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08324_ (.A1(_03263_),
    .A2(_03264_),
    .ZN(_03265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08325_ (.A1(_03262_),
    .A2(_03265_),
    .ZN(_03266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08326_ (.A1(_03259_),
    .A2(_03266_),
    .ZN(_03267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08327_ (.A1(_03267_),
    .A2(_01431_),
    .ZN(_03268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08328_ (.A1(_03252_),
    .A2(_03268_),
    .ZN(_03269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08329_ (.A1(_01376_),
    .A2(_01349_),
    .A3(\mem[20][14] ),
    .ZN(_03270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08330_ (.A1(_01057_),
    .A2(_01409_),
    .A3(\mem[19][14] ),
    .ZN(_03271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08331_ (.A1(_03270_),
    .A2(_03271_),
    .ZN(_03272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08332_ (.A1(_01067_),
    .A2(_01487_),
    .A3(\mem[21][14] ),
    .ZN(_03273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08333_ (.A1(_01161_),
    .A2(\mem[22][14] ),
    .ZN(_03274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08334_ (.A1(_03273_),
    .A2(_03274_),
    .ZN(_03275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08335_ (.A1(_03272_),
    .A2(_03275_),
    .ZN(_03276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08336_ (.A1(_02067_),
    .A2(_01467_),
    .A3(\mem[18][14] ),
    .ZN(_03277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08337_ (.A1(_02069_),
    .A2(_01443_),
    .A3(\mem[17][14] ),
    .ZN(_03278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08338_ (.A1(_03277_),
    .A2(_03278_),
    .ZN(_03279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08339_ (.A1(_01172_),
    .A2(\mem[23][14] ),
    .ZN(_03280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08340_ (.A1(_02073_),
    .A2(_01494_),
    .A3(\mem[16][14] ),
    .ZN(_03281_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08341_ (.A1(_03280_),
    .A2(_03281_),
    .ZN(_03282_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08342_ (.A1(_03279_),
    .A2(_03282_),
    .ZN(_03283_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08343_ (.A1(_03276_),
    .A2(_03283_),
    .ZN(_03284_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08344_ (.A1(_03284_),
    .A2(_01082_),
    .ZN(_03285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08345_ (.A1(_01408_),
    .A2(_01289_),
    .A3(\mem[28][14] ),
    .ZN(_03286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08346_ (.A1(_01483_),
    .A2(_01473_),
    .A3(_01153_),
    .A4(\mem[27][14] ),
    .ZN(_03287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08347_ (.A1(_03286_),
    .A2(_03287_),
    .ZN(_03288_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08348_ (.A1(_01055_),
    .A2(_01044_),
    .A3(_01491_),
    .A4(\mem[29][14] ),
    .ZN(_03289_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08349_ (.A1(_01041_),
    .A2(_01484_),
    .A3(_01047_),
    .A4(\mem[30][14] ),
    .ZN(_03290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08350_ (.A1(_03289_),
    .A2(_03290_),
    .ZN(_03291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08351_ (.A1(_03288_),
    .A2(_03291_),
    .ZN(_03292_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08352_ (.A1(_01476_),
    .A2(_01065_),
    .A3(_01470_),
    .A4(\mem[26][14] ),
    .ZN(_03293_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08353_ (.A1(_01424_),
    .A2(_01490_),
    .A3(\mem[25][14] ),
    .ZN(_03294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08354_ (.A1(_03293_),
    .A2(_03294_),
    .ZN(_03295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08355_ (.A1(_01469_),
    .A2(_01477_),
    .A3(_02223_),
    .A4(\mem[31][14] ),
    .ZN(_03296_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08356_ (.A1(_01049_),
    .A2(_01482_),
    .A3(\mem[24][14] ),
    .ZN(_03297_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08357_ (.A1(_03296_),
    .A2(_03297_),
    .ZN(_03298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08358_ (.A1(_03295_),
    .A2(_03298_),
    .ZN(_03299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08359_ (.A1(_03292_),
    .A2(_03299_),
    .ZN(_03300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08360_ (.A1(_03300_),
    .A2(_01104_),
    .ZN(_03301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08361_ (.A1(_03285_),
    .A2(_03301_),
    .ZN(_03302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08362_ (.A1(_03269_),
    .A2(_03302_),
    .ZN(_03303_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08363_ (.A1(_03236_),
    .A2(_03303_),
    .ZN(_00005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08364_ (.A1(_01263_),
    .A2(_01247_),
    .A3(\mem[36][15] ),
    .ZN(_03304_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08365_ (.A1(_01279_),
    .A2(_01249_),
    .A3(\mem[35][15] ),
    .ZN(_03305_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08366_ (.A1(_03304_),
    .A2(_03305_),
    .ZN(_03306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08367_ (.A1(_01401_),
    .A2(_01269_),
    .A3(\mem[37][15] ),
    .ZN(_03307_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08368_ (.A1(_01275_),
    .A2(\mem[38][15] ),
    .ZN(_03308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08369_ (.A1(_03307_),
    .A2(_03308_),
    .ZN(_03309_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08370_ (.A1(_03306_),
    .A2(_03309_),
    .ZN(_03310_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08371_ (.A1(_01237_),
    .A2(_01264_),
    .A3(\mem[34][15] ),
    .ZN(_03311_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08372_ (.A1(_01282_),
    .A2(_01242_),
    .A3(\mem[33][15] ),
    .ZN(_03312_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08373_ (.A1(_03311_),
    .A2(_03312_),
    .ZN(_03313_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08374_ (.A1(_01286_),
    .A2(\mem[39][15] ),
    .ZN(_03314_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08375_ (.A1(_01418_),
    .A2(_01450_),
    .A3(\mem[32][15] ),
    .ZN(_03315_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08376_ (.A1(_03314_),
    .A2(_03315_),
    .ZN(_03316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08377_ (.A1(_03313_),
    .A2(_03316_),
    .ZN(_03317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08378_ (.A1(_03310_),
    .A2(_03317_),
    .ZN(_03318_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08379_ (.A1(_03318_),
    .A2(_01127_),
    .ZN(_03319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08380_ (.A1(_01369_),
    .A2(_01370_),
    .A3(\mem[44][15] ),
    .ZN(_03320_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08381_ (.A1(_01383_),
    .A2(_01373_),
    .A3(\mem[43][15] ),
    .ZN(_03321_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08382_ (.A1(_03320_),
    .A2(_03321_),
    .ZN(_03322_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08383_ (.A1(_01435_),
    .A2(_01387_),
    .A3(\mem[45][15] ),
    .ZN(_03323_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08384_ (.A1(_01379_),
    .A2(\mem[46][15] ),
    .ZN(_03324_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08385_ (.A1(_03323_),
    .A2(_03324_),
    .ZN(_03325_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08386_ (.A1(_03322_),
    .A2(_03325_),
    .ZN(_03326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08387_ (.A1(_01268_),
    .A2(_01298_),
    .A3(\mem[42][15] ),
    .ZN(_03327_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08388_ (.A1(_01386_),
    .A2(_01301_),
    .A3(\mem[41][15] ),
    .ZN(_03328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08389_ (.A1(_03327_),
    .A2(_03328_),
    .ZN(_03329_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08390_ (.A1(_01390_),
    .A2(\mem[47][15] ),
    .ZN(_03330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08391_ (.A1(_01452_),
    .A2(_01393_),
    .A3(\mem[40][15] ),
    .ZN(_03331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08392_ (.A1(_03330_),
    .A2(_03331_),
    .ZN(_03332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08393_ (.A1(_03329_),
    .A2(_03332_),
    .ZN(_03333_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08394_ (.A1(_03326_),
    .A2(_03333_),
    .ZN(_03334_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08395_ (.A1(_03334_),
    .A2(_01149_),
    .ZN(_03335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08396_ (.A1(_03319_),
    .A2(_03335_),
    .ZN(_03336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08397_ (.A1(_01241_),
    .A2(_01384_),
    .A3(\mem[52][15] ),
    .ZN(_03337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08398_ (.A1(_01415_),
    .A2(_01273_),
    .A3(\mem[51][15] ),
    .ZN(_03338_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08399_ (.A1(_03337_),
    .A2(_03338_),
    .ZN(_03339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08400_ (.A1(_01466_),
    .A2(_01337_),
    .A3(\mem[53][15] ),
    .ZN(_03340_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08401_ (.A1(_01411_),
    .A2(\mem[54][15] ),
    .ZN(_03341_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08402_ (.A1(_03340_),
    .A2(_03341_),
    .ZN(_03342_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08403_ (.A1(_03339_),
    .A2(_03342_),
    .ZN(_03343_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08404_ (.A1(_01300_),
    .A2(_01402_),
    .A3(\mem[50][15] ),
    .ZN(_03344_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08405_ (.A1(_01254_),
    .A2(_01405_),
    .A3(\mem[49][15] ),
    .ZN(_03345_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08406_ (.A1(_03344_),
    .A2(_03345_),
    .ZN(_03346_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08407_ (.A1(_01422_),
    .A2(\mem[55][15] ),
    .ZN(_03347_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08408_ (.A1(_01486_),
    .A2(_01425_),
    .A3(\mem[48][15] ),
    .ZN(_03348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08409_ (.A1(_03347_),
    .A2(_03348_),
    .ZN(_03349_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08410_ (.A1(_03346_),
    .A2(_03349_),
    .ZN(_03350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08411_ (.A1(_03343_),
    .A2(_03350_),
    .ZN(_03351_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08412_ (.A1(_03351_),
    .A2(_01330_),
    .ZN(_03352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08413_ (.A1(_01272_),
    .A2(_01416_),
    .A3(\mem[60][15] ),
    .ZN(_03353_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08414_ (.A1(_01449_),
    .A2(_01419_),
    .A3(\mem[59][15] ),
    .ZN(_03354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08415_ (.A1(_03353_),
    .A2(_03354_),
    .ZN(_03355_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08416_ (.A1(_01442_),
    .A2(_01453_),
    .A3(\mem[61][15] ),
    .ZN(_03356_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08417_ (.A1(_01445_),
    .A2(\mem[62][15] ),
    .ZN(_03357_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08418_ (.A1(_03356_),
    .A2(_03357_),
    .ZN(_03358_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08419_ (.A1(_03355_),
    .A2(_03358_),
    .ZN(_03359_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08420_ (.A1(_01336_),
    .A2(_01256_),
    .A3(\mem[58][15] ),
    .ZN(_03360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08421_ (.A1(_01288_),
    .A2(_01342_),
    .A3(\mem[57][15] ),
    .ZN(_03361_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08422_ (.A1(_03360_),
    .A2(_03361_),
    .ZN(_03362_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08423_ (.A1(_01456_),
    .A2(\mem[63][15] ),
    .ZN(_03363_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08424_ (.A1(_01458_),
    .A2(_01459_),
    .A3(\mem[56][15] ),
    .ZN(_03364_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08425_ (.A1(_03363_),
    .A2(_03364_),
    .ZN(_03365_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08426_ (.A1(_03362_),
    .A2(_03365_),
    .ZN(_03366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08427_ (.A1(_03359_),
    .A2(_03366_),
    .ZN(_03367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08428_ (.A1(_03367_),
    .A2(_01364_),
    .ZN(_03368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08429_ (.A1(_03352_),
    .A2(_03368_),
    .ZN(_03369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08430_ (.A1(_03336_),
    .A2(_03369_),
    .ZN(_03370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08431_ (.A1(_01297_),
    .A2(_01280_),
    .A3(\mem[4][15] ),
    .ZN(_03371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08432_ (.A1(_01312_),
    .A2(_01283_),
    .A3(\mem[3][15] ),
    .ZN(_03372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08433_ (.A1(_03371_),
    .A2(_03372_),
    .ZN(_03373_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08434_ (.A1(_01304_),
    .A2(_01317_),
    .A3(\mem[5][15] ),
    .ZN(_03374_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08435_ (.A1(_01308_),
    .A2(\mem[6][15] ),
    .ZN(_03375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08436_ (.A1(_03374_),
    .A2(_03375_),
    .ZN(_03376_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08437_ (.A1(_03373_),
    .A2(_03376_),
    .ZN(_03377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08438_ (.A1(_01372_),
    .A2(_01314_),
    .A3(\mem[2][15] ),
    .ZN(_03378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08439_ (.A1(_01316_),
    .A2(_01377_),
    .A3(\mem[1][15] ),
    .ZN(_03379_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08440_ (.A1(_03378_),
    .A2(_03379_),
    .ZN(_03380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08441_ (.A1(_01320_),
    .A2(\mem[7][15] ),
    .ZN(_03381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08442_ (.A1(_01323_),
    .A2(_01324_),
    .A3(\mem[0][15] ),
    .ZN(_03382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08443_ (.A1(_03381_),
    .A2(_03382_),
    .ZN(_03383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08444_ (.A1(_03380_),
    .A2(_03383_),
    .ZN(_03384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08445_ (.A1(_03377_),
    .A2(_03384_),
    .ZN(_03385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08446_ (.A1(_03385_),
    .A2(_01398_),
    .ZN(_03386_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08447_ (.A1(_01333_),
    .A2(_01334_),
    .A3(\mem[12][15] ),
    .ZN(_03387_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08448_ (.A1(_01348_),
    .A2(_01306_),
    .A3(\mem[11][15] ),
    .ZN(_03388_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08449_ (.A1(_03387_),
    .A2(_03388_),
    .ZN(_03389_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08450_ (.A1(_01340_),
    .A2(_01352_),
    .A3(\mem[13][15] ),
    .ZN(_03390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08451_ (.A1(_01344_),
    .A2(\mem[14][15] ),
    .ZN(_03391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08452_ (.A1(_03390_),
    .A2(_03391_),
    .ZN(_03392_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08453_ (.A1(_03389_),
    .A2(_03392_),
    .ZN(_03393_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08454_ (.A1(_01404_),
    .A2(_01436_),
    .A3(\mem[10][15] ),
    .ZN(_03394_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08455_ (.A1(_01351_),
    .A2(_01439_),
    .A3(\mem[9][15] ),
    .ZN(_03395_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08456_ (.A1(_03394_),
    .A2(_03395_),
    .ZN(_03396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08457_ (.A1(_01355_),
    .A2(\mem[15][15] ),
    .ZN(_03397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08458_ (.A1(_01357_),
    .A2(_01359_),
    .A3(\mem[8][15] ),
    .ZN(_03398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08459_ (.A1(_03397_),
    .A2(_03398_),
    .ZN(_03399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08460_ (.A1(_03396_),
    .A2(_03399_),
    .ZN(_03400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08461_ (.A1(_03393_),
    .A2(_03400_),
    .ZN(_03401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08462_ (.A1(_03401_),
    .A2(_01431_),
    .ZN(_03402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08463_ (.A1(_03386_),
    .A2(_03402_),
    .ZN(_03403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08464_ (.A1(_01376_),
    .A2(_01349_),
    .A3(\mem[20][15] ),
    .ZN(_03404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08465_ (.A1(_01057_),
    .A2(_01409_),
    .A3(\mem[19][15] ),
    .ZN(_03405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08466_ (.A1(_03404_),
    .A2(_03405_),
    .ZN(_03406_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08467_ (.A1(_01067_),
    .A2(_01487_),
    .A3(\mem[21][15] ),
    .ZN(_03407_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08468_ (.A1(_01161_),
    .A2(\mem[22][15] ),
    .ZN(_03408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08469_ (.A1(_03407_),
    .A2(_03408_),
    .ZN(_03409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08470_ (.A1(_03406_),
    .A2(_03409_),
    .ZN(_03410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08471_ (.A1(_01438_),
    .A2(_01467_),
    .A3(\mem[18][15] ),
    .ZN(_03411_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08472_ (.A1(_01392_),
    .A2(_01443_),
    .A3(\mem[17][15] ),
    .ZN(_03412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08473_ (.A1(_03411_),
    .A2(_03412_),
    .ZN(_03413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08474_ (.A1(_01172_),
    .A2(\mem[23][15] ),
    .ZN(_03414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08475_ (.A1(_01493_),
    .A2(_01494_),
    .A3(\mem[16][15] ),
    .ZN(_03415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08476_ (.A1(_03414_),
    .A2(_03415_),
    .ZN(_03416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08477_ (.A1(_03413_),
    .A2(_03416_),
    .ZN(_03417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08478_ (.A1(_03410_),
    .A2(_03417_),
    .ZN(_03418_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08479_ (.A1(_03418_),
    .A2(_01082_),
    .ZN(_03419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08480_ (.A1(_01408_),
    .A2(_01289_),
    .A3(\mem[28][15] ),
    .ZN(_03420_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08481_ (.A1(_01483_),
    .A2(_01473_),
    .A3(_01153_),
    .A4(\mem[27][15] ),
    .ZN(_03421_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08482_ (.A1(_03420_),
    .A2(_03421_),
    .ZN(_03422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08483_ (.A1(_01055_),
    .A2(_01044_),
    .A3(_01491_),
    .A4(\mem[29][15] ),
    .ZN(_03423_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08484_ (.A1(_01041_),
    .A2(_01484_),
    .A3(_01047_),
    .A4(\mem[30][15] ),
    .ZN(_03424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08485_ (.A1(_03423_),
    .A2(_03424_),
    .ZN(_03425_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08486_ (.A1(_03422_),
    .A2(_03425_),
    .ZN(_03426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08487_ (.A1(_01476_),
    .A2(_01065_),
    .A3(_01470_),
    .A4(\mem[26][15] ),
    .ZN(_03427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08488_ (.A1(_01424_),
    .A2(_01490_),
    .A3(\mem[25][15] ),
    .ZN(_03428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08489_ (.A1(_03427_),
    .A2(_03428_),
    .ZN(_03429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08490_ (.A1(_01469_),
    .A2(_01477_),
    .A3(_02223_),
    .A4(\mem[31][15] ),
    .ZN(_03430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08491_ (.A1(_01049_),
    .A2(_01482_),
    .A3(\mem[24][15] ),
    .ZN(_03431_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08492_ (.A1(_03430_),
    .A2(_03431_),
    .ZN(_03432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08493_ (.A1(_03429_),
    .A2(_03432_),
    .ZN(_03433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08494_ (.A1(_03426_),
    .A2(_03433_),
    .ZN(_03434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08495_ (.A1(_03434_),
    .A2(_01104_),
    .ZN(_03435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08496_ (.A1(_03419_),
    .A2(_03435_),
    .ZN(_03436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08497_ (.A1(_03403_),
    .A2(_03436_),
    .ZN(_03437_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08498_ (.A1(_03370_),
    .A2(_03437_),
    .ZN(_00006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _08499_ (.I(net100),
    .ZN(_03438_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08500_ (.I(_03438_),
    .Z(_03439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08501_ (.I(net91),
    .ZN(_03440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08502_ (.A1(net59),
    .A2(_01313_),
    .A3(_03440_),
    .ZN(_03441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08503_ (.A1(net60),
    .A2(_01398_),
    .ZN(_03442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08504_ (.I(net61),
    .Z(_03443_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08505_ (.I(net61),
    .Z(_03444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08506_ (.A1(_03444_),
    .A2(\mem[7][13] ),
    .ZN(_03445_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08507_ (.A1(_03439_),
    .A2(net62),
    .B(_03445_),
    .ZN(_00016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08508_ (.I(net84),
    .ZN(_03446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08509_ (.I(_03446_),
    .Z(_03447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08510_ (.A1(_03444_),
    .A2(\mem[7][14] ),
    .ZN(_03448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08511_ (.A1(_03447_),
    .A2(net62),
    .B(_03448_),
    .ZN(_00017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08512_ (.I(net55),
    .ZN(_03449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08513_ (.I(_03449_),
    .Z(_03450_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08514_ (.A1(_03444_),
    .A2(\mem[7][15] ),
    .ZN(_03451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08515_ (.A1(_03450_),
    .A2(net62),
    .B(_03451_),
    .ZN(_00018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08516_ (.I(net82),
    .ZN(_03452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08517_ (.I(_03452_),
    .Z(_03453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08518_ (.A1(net87),
    .A2(_03440_),
    .ZN(_03454_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08519_ (.A1(_01266_),
    .A2(_01043_),
    .ZN(_03455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _08520_ (.I(_03455_),
    .ZN(_03456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08521_ (.A1(net88),
    .A2(_03456_),
    .ZN(_03457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08522_ (.I(_03457_),
    .Z(_03458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08523_ (.I(_03457_),
    .Z(_03459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08524_ (.A1(_03459_),
    .A2(\mem[59][0] ),
    .ZN(_03460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08525_ (.A1(_03453_),
    .A2(_03458_),
    .B(_03460_),
    .ZN(_00019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08526_ (.I(net43),
    .ZN(_03461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08527_ (.I(_03461_),
    .Z(_03462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08528_ (.A1(_03459_),
    .A2(\mem[59][1] ),
    .ZN(_03463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08529_ (.A1(_03462_),
    .A2(_03458_),
    .B(_03463_),
    .ZN(_00020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08530_ (.I(net80),
    .ZN(_03464_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08531_ (.I(_03464_),
    .Z(_03465_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08532_ (.A1(_03459_),
    .A2(\mem[59][2] ),
    .ZN(_03466_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08533_ (.A1(_03465_),
    .A2(_03458_),
    .B(_03466_),
    .ZN(_00021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08534_ (.I(net52),
    .ZN(_03467_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08535_ (.I(_03467_),
    .Z(_03468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08536_ (.A1(_03459_),
    .A2(\mem[59][3] ),
    .ZN(_03469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08537_ (.A1(_03468_),
    .A2(_03458_),
    .B(_03469_),
    .ZN(_00022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08538_ (.I(net46),
    .ZN(_03470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08539_ (.I(_03470_),
    .Z(_03471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08540_ (.I(_03457_),
    .Z(_03472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08541_ (.A1(_03472_),
    .A2(\mem[59][4] ),
    .ZN(_03473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08542_ (.A1(_03471_),
    .A2(_03458_),
    .B(_03473_),
    .ZN(_00023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08543_ (.I(net49),
    .ZN(_03474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08544_ (.I(_03474_),
    .Z(_03475_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08545_ (.A1(_03472_),
    .A2(\mem[59][5] ),
    .ZN(_03476_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08546_ (.A1(_03475_),
    .A2(_03458_),
    .B(_03476_),
    .ZN(_00024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08547_ (.I(net65),
    .ZN(_03477_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08548_ (.I(_03477_),
    .Z(_03478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08549_ (.A1(_03472_),
    .A2(\mem[59][6] ),
    .ZN(_03479_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08550_ (.A1(_03478_),
    .A2(_03458_),
    .B(_03479_),
    .ZN(_00025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08551_ (.I(net95),
    .ZN(_03480_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08552_ (.I(_03480_),
    .Z(_03481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08553_ (.A1(_03472_),
    .A2(\mem[59][7] ),
    .ZN(_03482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08554_ (.A1(_03481_),
    .A2(_03458_),
    .B(_03482_),
    .ZN(_00026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _08555_ (.I(net106),
    .ZN(_03483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08556_ (.I(_03483_),
    .Z(_03484_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08557_ (.A1(_03472_),
    .A2(\mem[59][8] ),
    .ZN(_03485_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08558_ (.A1(_03484_),
    .A2(_03458_),
    .B(_03485_),
    .ZN(_00027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_8 _08559_ (.I(net114),
    .ZN(_03486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08560_ (.I(_03486_),
    .Z(_03487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08561_ (.A1(_03472_),
    .A2(\mem[59][9] ),
    .ZN(_03488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08562_ (.A1(_03487_),
    .A2(_03458_),
    .B(_03488_),
    .ZN(_00028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08563_ (.I(net112),
    .ZN(_03489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08564_ (.I(_03489_),
    .Z(_03490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08565_ (.A1(_03472_),
    .A2(\mem[59][10] ),
    .ZN(_03491_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08566_ (.A1(_03490_),
    .A2(_03459_),
    .B(_03491_),
    .ZN(_00029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08567_ (.I(net104),
    .ZN(_03492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08568_ (.I(_03492_),
    .Z(_03493_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08569_ (.A1(_03472_),
    .A2(\mem[59][11] ),
    .ZN(_03494_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08570_ (.A1(_03493_),
    .A2(_03459_),
    .B(_03494_),
    .ZN(_00030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08571_ (.I(net102),
    .ZN(_03495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08572_ (.I(_03495_),
    .Z(_03496_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08573_ (.A1(_03472_),
    .A2(\mem[59][12] ),
    .ZN(_03497_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08574_ (.A1(_03496_),
    .A2(_03459_),
    .B(_03497_),
    .ZN(_00031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08575_ (.A1(_03472_),
    .A2(\mem[59][13] ),
    .ZN(_03498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08576_ (.A1(_03439_),
    .A2(_03459_),
    .B(_03498_),
    .ZN(_00032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08577_ (.A1(_03457_),
    .A2(\mem[59][14] ),
    .ZN(_03499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08578_ (.A1(_03447_),
    .A2(_03459_),
    .B(_03499_),
    .ZN(_00033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08579_ (.A1(_03457_),
    .A2(\mem[59][15] ),
    .ZN(_03500_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08580_ (.A1(_03450_),
    .A2(_03459_),
    .B(_03500_),
    .ZN(_00034_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08581_ (.A1(net40),
    .A2(_01364_),
    .ZN(_03501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08582_ (.I(_03501_),
    .Z(_03502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08583_ (.I(_03501_),
    .Z(_03503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08584_ (.A1(_03503_),
    .A2(\mem[63][0] ),
    .ZN(_03504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08585_ (.A1(_03453_),
    .A2(_03502_),
    .B(_03504_),
    .ZN(_00035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08586_ (.A1(_03503_),
    .A2(\mem[63][1] ),
    .ZN(_03505_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08587_ (.A1(_03462_),
    .A2(_03502_),
    .B(_03505_),
    .ZN(_00036_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08588_ (.A1(_03503_),
    .A2(\mem[63][2] ),
    .ZN(_03506_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08589_ (.A1(_03465_),
    .A2(_03502_),
    .B(_03506_),
    .ZN(_00037_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08590_ (.A1(_03503_),
    .A2(\mem[63][3] ),
    .ZN(_03507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08591_ (.A1(_03468_),
    .A2(_03502_),
    .B(_03507_),
    .ZN(_00038_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08592_ (.I(_03501_),
    .Z(_03508_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08593_ (.A1(_03508_),
    .A2(\mem[63][4] ),
    .ZN(_03509_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08594_ (.A1(_03471_),
    .A2(_03502_),
    .B(_03509_),
    .ZN(_00039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08595_ (.A1(_03508_),
    .A2(\mem[63][5] ),
    .ZN(_03510_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08596_ (.A1(_03475_),
    .A2(_03502_),
    .B(_03510_),
    .ZN(_00040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08597_ (.A1(_03508_),
    .A2(\mem[63][6] ),
    .ZN(_03511_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08598_ (.A1(_03478_),
    .A2(_03502_),
    .B(_03511_),
    .ZN(_00041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08599_ (.A1(_03508_),
    .A2(\mem[63][7] ),
    .ZN(_03512_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08600_ (.A1(_03481_),
    .A2(_03502_),
    .B(_03512_),
    .ZN(_00042_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08601_ (.A1(_03508_),
    .A2(\mem[63][8] ),
    .ZN(_03513_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08602_ (.A1(_03484_),
    .A2(_03502_),
    .B(_03513_),
    .ZN(_00043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08603_ (.A1(_03508_),
    .A2(\mem[63][9] ),
    .ZN(_03514_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08604_ (.A1(_03487_),
    .A2(_03502_),
    .B(_03514_),
    .ZN(_00044_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08605_ (.A1(_03508_),
    .A2(\mem[63][10] ),
    .ZN(_03515_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08606_ (.A1(_03490_),
    .A2(_03503_),
    .B(_03515_),
    .ZN(_00045_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08607_ (.A1(_03508_),
    .A2(\mem[63][11] ),
    .ZN(_03516_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08608_ (.A1(_03493_),
    .A2(_03503_),
    .B(_03516_),
    .ZN(_00046_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08609_ (.A1(_03508_),
    .A2(\mem[63][12] ),
    .ZN(_03517_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08610_ (.A1(_03496_),
    .A2(_03503_),
    .B(_03517_),
    .ZN(_00047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08611_ (.A1(_03508_),
    .A2(\mem[63][13] ),
    .ZN(_03518_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08612_ (.A1(_03439_),
    .A2(_03503_),
    .B(_03518_),
    .ZN(_00048_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08613_ (.A1(_03501_),
    .A2(\mem[63][14] ),
    .ZN(_03519_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08614_ (.A1(_03447_),
    .A2(_03503_),
    .B(_03519_),
    .ZN(_00049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08615_ (.A1(_03501_),
    .A2(\mem[63][15] ),
    .ZN(_03520_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08616_ (.A1(_03450_),
    .A2(_03503_),
    .B(_03520_),
    .ZN(_00050_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08617_ (.A1(_01398_),
    .A2(net91),
    .ZN(_03521_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _08618_ (.I(net124),
    .ZN(_03522_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08619_ (.A1(_03522_),
    .A2(_01162_),
    .ZN(_03523_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08620_ (.I(_03523_),
    .Z(_03524_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08621_ (.I(_03523_),
    .Z(_03525_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08622_ (.A1(_03525_),
    .A2(\mem[6][0] ),
    .ZN(_03526_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08623_ (.A1(_03453_),
    .A2(_03524_),
    .B(_03526_),
    .ZN(_00051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08624_ (.A1(_03525_),
    .A2(\mem[6][1] ),
    .ZN(_03527_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08625_ (.A1(_03462_),
    .A2(_03524_),
    .B(_03527_),
    .ZN(_00052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08626_ (.A1(_03525_),
    .A2(\mem[6][2] ),
    .ZN(_03528_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08627_ (.A1(_03465_),
    .A2(_03524_),
    .B(_03528_),
    .ZN(_00053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08628_ (.A1(_03525_),
    .A2(\mem[6][3] ),
    .ZN(_03529_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08629_ (.A1(_03468_),
    .A2(_03524_),
    .B(_03529_),
    .ZN(_00054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08630_ (.I(_03523_),
    .Z(_03530_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08631_ (.A1(_03530_),
    .A2(\mem[6][4] ),
    .ZN(_03531_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08632_ (.A1(_03471_),
    .A2(_03524_),
    .B(_03531_),
    .ZN(_00055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08633_ (.A1(_03530_),
    .A2(\mem[6][5] ),
    .ZN(_03532_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08634_ (.A1(_03475_),
    .A2(_03524_),
    .B(_03532_),
    .ZN(_00056_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08635_ (.A1(_03530_),
    .A2(\mem[6][6] ),
    .ZN(_03533_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08636_ (.A1(_03478_),
    .A2(_03524_),
    .B(_03533_),
    .ZN(_00057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08637_ (.A1(_03530_),
    .A2(\mem[6][7] ),
    .ZN(_03534_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08638_ (.A1(_03481_),
    .A2(_03524_),
    .B(_03534_),
    .ZN(_00058_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08639_ (.A1(_03530_),
    .A2(\mem[6][8] ),
    .ZN(_03535_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08640_ (.A1(_03484_),
    .A2(_03524_),
    .B(_03535_),
    .ZN(_00059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08641_ (.A1(_03530_),
    .A2(\mem[6][9] ),
    .ZN(_03536_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08642_ (.A1(_03487_),
    .A2(_03524_),
    .B(_03536_),
    .ZN(_00060_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08643_ (.A1(_03530_),
    .A2(\mem[6][10] ),
    .ZN(_03537_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08644_ (.A1(_03490_),
    .A2(_03525_),
    .B(_03537_),
    .ZN(_00061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08645_ (.A1(_03530_),
    .A2(\mem[6][11] ),
    .ZN(_03538_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08646_ (.A1(_03493_),
    .A2(_03525_),
    .B(_03538_),
    .ZN(_00062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08647_ (.A1(_03530_),
    .A2(\mem[6][12] ),
    .ZN(_03539_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08648_ (.A1(_03496_),
    .A2(_03525_),
    .B(_03539_),
    .ZN(_00063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08649_ (.A1(_03530_),
    .A2(\mem[6][13] ),
    .ZN(_03540_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08650_ (.A1(_03439_),
    .A2(_03525_),
    .B(_03540_),
    .ZN(_00064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08651_ (.A1(_03523_),
    .A2(\mem[6][14] ),
    .ZN(_03541_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08652_ (.A1(_03447_),
    .A2(_03525_),
    .B(_03541_),
    .ZN(_00065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08653_ (.A1(_03523_),
    .A2(\mem[6][15] ),
    .ZN(_03542_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08654_ (.A1(_03450_),
    .A2(_03525_),
    .B(_03542_),
    .ZN(_00066_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08655_ (.A1(_03455_),
    .A2(_03440_),
    .ZN(_03543_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08656_ (.A1(_03543_),
    .A2(_01082_),
    .ZN(_03544_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08657_ (.I(_03544_),
    .Z(_03545_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08658_ (.I(_03544_),
    .Z(_03546_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08659_ (.A1(_03546_),
    .A2(\mem[19][0] ),
    .ZN(_03547_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08660_ (.A1(_03453_),
    .A2(_03545_),
    .B(_03547_),
    .ZN(_00067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08661_ (.A1(_03546_),
    .A2(\mem[19][1] ),
    .ZN(_03548_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08662_ (.A1(_03462_),
    .A2(_03545_),
    .B(_03548_),
    .ZN(_00068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08663_ (.A1(_03546_),
    .A2(\mem[19][2] ),
    .ZN(_03549_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08664_ (.A1(_03465_),
    .A2(_03545_),
    .B(_03549_),
    .ZN(_00069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08665_ (.A1(_03546_),
    .A2(\mem[19][3] ),
    .ZN(_03550_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08666_ (.A1(_03468_),
    .A2(_03545_),
    .B(_03550_),
    .ZN(_00070_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08667_ (.I(_03544_),
    .Z(_03551_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08668_ (.A1(_03551_),
    .A2(\mem[19][4] ),
    .ZN(_03552_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08669_ (.A1(_03471_),
    .A2(_03545_),
    .B(_03552_),
    .ZN(_00071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08670_ (.A1(_03551_),
    .A2(\mem[19][5] ),
    .ZN(_03553_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08671_ (.A1(_03475_),
    .A2(_03545_),
    .B(_03553_),
    .ZN(_00072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08672_ (.A1(_03551_),
    .A2(\mem[19][6] ),
    .ZN(_03554_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08673_ (.A1(_03478_),
    .A2(_03545_),
    .B(_03554_),
    .ZN(_00073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08674_ (.A1(_03551_),
    .A2(\mem[19][7] ),
    .ZN(_03555_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08675_ (.A1(_03481_),
    .A2(_03545_),
    .B(_03555_),
    .ZN(_00074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08676_ (.A1(_03551_),
    .A2(\mem[19][8] ),
    .ZN(_03556_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08677_ (.A1(_03484_),
    .A2(_03545_),
    .B(_03556_),
    .ZN(_00075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08678_ (.A1(_03551_),
    .A2(\mem[19][9] ),
    .ZN(_03557_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08679_ (.A1(_03487_),
    .A2(_03545_),
    .B(_03557_),
    .ZN(_00076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08680_ (.A1(_03551_),
    .A2(\mem[19][10] ),
    .ZN(_03558_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08681_ (.A1(_03490_),
    .A2(_03546_),
    .B(_03558_),
    .ZN(_00077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08682_ (.A1(_03551_),
    .A2(\mem[19][11] ),
    .ZN(_03559_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08683_ (.A1(_03493_),
    .A2(_03546_),
    .B(_03559_),
    .ZN(_00078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08684_ (.A1(_03551_),
    .A2(\mem[19][12] ),
    .ZN(_03560_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08685_ (.A1(_03496_),
    .A2(_03546_),
    .B(_03560_),
    .ZN(_00079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08686_ (.A1(_03551_),
    .A2(\mem[19][13] ),
    .ZN(_03561_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08687_ (.A1(_03439_),
    .A2(_03546_),
    .B(_03561_),
    .ZN(_00080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08688_ (.A1(_03544_),
    .A2(\mem[19][14] ),
    .ZN(_03562_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08689_ (.A1(_03447_),
    .A2(_03546_),
    .B(_03562_),
    .ZN(_00081_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08690_ (.A1(_03544_),
    .A2(\mem[19][15] ),
    .ZN(_03563_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08691_ (.A1(_03450_),
    .A2(_03546_),
    .B(_03563_),
    .ZN(_00082_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08692_ (.A1(net118),
    .A2(_03440_),
    .ZN(_03564_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08693_ (.A1(_01066_),
    .A2(_01341_),
    .ZN(_03565_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _08694_ (.I(_03565_),
    .ZN(_03566_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08695_ (.A1(net119),
    .A2(_03566_),
    .ZN(_03567_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08696_ (.I(_03567_),
    .Z(_03568_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08697_ (.I(_03567_),
    .Z(_03569_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08698_ (.A1(_03569_),
    .A2(\mem[29][0] ),
    .ZN(_03570_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08699_ (.A1(_03453_),
    .A2(_03568_),
    .B(_03570_),
    .ZN(_00083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08700_ (.A1(_03569_),
    .A2(\mem[29][1] ),
    .ZN(_03571_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08701_ (.A1(_03462_),
    .A2(_03568_),
    .B(_03571_),
    .ZN(_00084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08702_ (.A1(_03569_),
    .A2(\mem[29][2] ),
    .ZN(_03572_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08703_ (.A1(_03465_),
    .A2(_03568_),
    .B(_03572_),
    .ZN(_00085_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08704_ (.A1(_03569_),
    .A2(\mem[29][3] ),
    .ZN(_03573_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08705_ (.A1(_03468_),
    .A2(_03568_),
    .B(_03573_),
    .ZN(_00086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08706_ (.I(_03567_),
    .Z(_03574_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08707_ (.A1(_03574_),
    .A2(\mem[29][4] ),
    .ZN(_03575_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08708_ (.A1(_03471_),
    .A2(_03568_),
    .B(_03575_),
    .ZN(_00087_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08709_ (.A1(_03574_),
    .A2(\mem[29][5] ),
    .ZN(_03576_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08710_ (.A1(_03475_),
    .A2(_03568_),
    .B(_03576_),
    .ZN(_00088_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08711_ (.A1(_03574_),
    .A2(\mem[29][6] ),
    .ZN(_03577_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08712_ (.A1(_03478_),
    .A2(_03568_),
    .B(_03577_),
    .ZN(_00089_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08713_ (.A1(_03574_),
    .A2(\mem[29][7] ),
    .ZN(_03578_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08714_ (.A1(_03481_),
    .A2(_03568_),
    .B(_03578_),
    .ZN(_00090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08715_ (.A1(_03574_),
    .A2(\mem[29][8] ),
    .ZN(_03579_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08716_ (.A1(_03484_),
    .A2(_03568_),
    .B(_03579_),
    .ZN(_00091_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08717_ (.A1(_03574_),
    .A2(\mem[29][9] ),
    .ZN(_03580_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08718_ (.A1(_03487_),
    .A2(_03568_),
    .B(_03580_),
    .ZN(_00092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08719_ (.A1(_03574_),
    .A2(\mem[29][10] ),
    .ZN(_03581_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08720_ (.A1(_03490_),
    .A2(_03569_),
    .B(_03581_),
    .ZN(_00093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08721_ (.A1(_03574_),
    .A2(\mem[29][11] ),
    .ZN(_03582_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08722_ (.A1(_03493_),
    .A2(_03569_),
    .B(_03582_),
    .ZN(_00094_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08723_ (.A1(_03574_),
    .A2(\mem[29][12] ),
    .ZN(_03583_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08724_ (.A1(_03496_),
    .A2(_03569_),
    .B(_03583_),
    .ZN(_00095_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08725_ (.A1(_03574_),
    .A2(\mem[29][13] ),
    .ZN(_03584_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08726_ (.A1(_03439_),
    .A2(_03569_),
    .B(_03584_),
    .ZN(_00096_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08727_ (.A1(_03567_),
    .A2(\mem[29][14] ),
    .ZN(_03585_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08728_ (.A1(_03447_),
    .A2(_03569_),
    .B(_03585_),
    .ZN(_00097_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08729_ (.A1(_03567_),
    .A2(\mem[29][15] ),
    .ZN(_03586_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08730_ (.A1(_03450_),
    .A2(_03569_),
    .B(_03586_),
    .ZN(_00098_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08731_ (.A1(net126),
    .A2(_01040_),
    .A3(net91),
    .ZN(_03587_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _08732_ (.I(net127),
    .ZN(_03588_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08733_ (.A1(_03588_),
    .A2(_01431_),
    .ZN(_03589_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08734_ (.I(_03589_),
    .Z(_03590_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08735_ (.I(_03589_),
    .Z(_03591_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08736_ (.A1(_03591_),
    .A2(\mem[8][0] ),
    .ZN(_03592_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08737_ (.A1(_03453_),
    .A2(_03590_),
    .B(_03592_),
    .ZN(_00099_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08738_ (.A1(_03591_),
    .A2(\mem[8][1] ),
    .ZN(_03593_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08739_ (.A1(_03462_),
    .A2(_03590_),
    .B(_03593_),
    .ZN(_00100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08740_ (.A1(_03591_),
    .A2(\mem[8][2] ),
    .ZN(_03594_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08741_ (.A1(_03465_),
    .A2(_03590_),
    .B(_03594_),
    .ZN(_00101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08742_ (.A1(_03591_),
    .A2(\mem[8][3] ),
    .ZN(_03595_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08743_ (.A1(_03468_),
    .A2(_03590_),
    .B(_03595_),
    .ZN(_00102_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08744_ (.I(_03589_),
    .Z(_03596_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08745_ (.A1(_03596_),
    .A2(\mem[8][4] ),
    .ZN(_03597_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08746_ (.A1(_03471_),
    .A2(_03590_),
    .B(_03597_),
    .ZN(_00103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08747_ (.A1(_03596_),
    .A2(\mem[8][5] ),
    .ZN(_03598_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08748_ (.A1(_03475_),
    .A2(_03590_),
    .B(_03598_),
    .ZN(_00104_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08749_ (.A1(_03596_),
    .A2(\mem[8][6] ),
    .ZN(_03599_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08750_ (.A1(_03478_),
    .A2(_03590_),
    .B(_03599_),
    .ZN(_00105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08751_ (.A1(_03596_),
    .A2(\mem[8][7] ),
    .ZN(_03600_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08752_ (.A1(_03481_),
    .A2(_03590_),
    .B(_03600_),
    .ZN(_00106_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08753_ (.A1(_03596_),
    .A2(\mem[8][8] ),
    .ZN(_03601_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08754_ (.A1(_03484_),
    .A2(_03590_),
    .B(_03601_),
    .ZN(_00107_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08755_ (.A1(_03596_),
    .A2(\mem[8][9] ),
    .ZN(_03602_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08756_ (.A1(_03487_),
    .A2(_03590_),
    .B(_03602_),
    .ZN(_00108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08757_ (.A1(_03596_),
    .A2(\mem[8][10] ),
    .ZN(_03603_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08758_ (.A1(_03490_),
    .A2(_03591_),
    .B(_03603_),
    .ZN(_00109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08759_ (.A1(_03596_),
    .A2(\mem[8][11] ),
    .ZN(_03604_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08760_ (.A1(_03493_),
    .A2(_03591_),
    .B(_03604_),
    .ZN(_00110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08761_ (.A1(_03596_),
    .A2(\mem[8][12] ),
    .ZN(_03605_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08762_ (.A1(_03496_),
    .A2(_03591_),
    .B(_03605_),
    .ZN(_00111_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08763_ (.A1(_03596_),
    .A2(\mem[8][13] ),
    .ZN(_03606_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08764_ (.A1(_03439_),
    .A2(_03591_),
    .B(_03606_),
    .ZN(_00112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08765_ (.A1(_03589_),
    .A2(\mem[8][14] ),
    .ZN(_03607_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08766_ (.A1(_03447_),
    .A2(_03591_),
    .B(_03607_),
    .ZN(_00113_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08767_ (.A1(_03589_),
    .A2(\mem[8][15] ),
    .ZN(_03608_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08768_ (.A1(_03450_),
    .A2(_03591_),
    .B(_03608_),
    .ZN(_00114_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08769_ (.A1(_03588_),
    .A2(_01398_),
    .ZN(_03609_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08770_ (.I(_03609_),
    .Z(_03610_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08771_ (.I(_03609_),
    .Z(_03611_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08772_ (.A1(_03611_),
    .A2(\mem[0][0] ),
    .ZN(_03612_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08773_ (.A1(_03453_),
    .A2(_03610_),
    .B(_03612_),
    .ZN(_00115_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08774_ (.A1(_03611_),
    .A2(\mem[0][1] ),
    .ZN(_03613_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08775_ (.A1(_03462_),
    .A2(_03610_),
    .B(_03613_),
    .ZN(_00116_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08776_ (.A1(_03611_),
    .A2(\mem[0][2] ),
    .ZN(_03614_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08777_ (.A1(_03465_),
    .A2(_03610_),
    .B(_03614_),
    .ZN(_00117_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08778_ (.A1(_03611_),
    .A2(\mem[0][3] ),
    .ZN(_03615_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08779_ (.A1(_03468_),
    .A2(_03610_),
    .B(_03615_),
    .ZN(_00118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08780_ (.I(_03609_),
    .Z(_03616_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08781_ (.A1(_03616_),
    .A2(\mem[0][4] ),
    .ZN(_03617_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08782_ (.A1(_03471_),
    .A2(_03610_),
    .B(_03617_),
    .ZN(_00119_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08783_ (.A1(_03616_),
    .A2(\mem[0][5] ),
    .ZN(_03618_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08784_ (.A1(_03475_),
    .A2(_03610_),
    .B(_03618_),
    .ZN(_00120_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08785_ (.A1(_03616_),
    .A2(\mem[0][6] ),
    .ZN(_03619_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08786_ (.A1(_03478_),
    .A2(_03610_),
    .B(_03619_),
    .ZN(_00121_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08787_ (.A1(_03616_),
    .A2(\mem[0][7] ),
    .ZN(_03620_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08788_ (.A1(_03481_),
    .A2(_03610_),
    .B(_03620_),
    .ZN(_00122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08789_ (.A1(_03616_),
    .A2(\mem[0][8] ),
    .ZN(_03621_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08790_ (.A1(_03484_),
    .A2(_03610_),
    .B(_03621_),
    .ZN(_00123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08791_ (.A1(_03616_),
    .A2(\mem[0][9] ),
    .ZN(_03622_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08792_ (.A1(_03487_),
    .A2(_03610_),
    .B(_03622_),
    .ZN(_00124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08793_ (.A1(_03616_),
    .A2(\mem[0][10] ),
    .ZN(_03623_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08794_ (.A1(_03490_),
    .A2(_03611_),
    .B(_03623_),
    .ZN(_00125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08795_ (.A1(_03616_),
    .A2(\mem[0][11] ),
    .ZN(_03624_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08796_ (.A1(_03493_),
    .A2(_03611_),
    .B(_03624_),
    .ZN(_00126_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08797_ (.A1(_03616_),
    .A2(\mem[0][12] ),
    .ZN(_03625_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08798_ (.A1(_03496_),
    .A2(_03611_),
    .B(_03625_),
    .ZN(_00127_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08799_ (.A1(_03616_),
    .A2(\mem[0][13] ),
    .ZN(_03626_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08800_ (.A1(_03439_),
    .A2(_03611_),
    .B(_03626_),
    .ZN(_00128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08801_ (.A1(_03609_),
    .A2(\mem[0][14] ),
    .ZN(_03627_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08802_ (.A1(_03447_),
    .A2(_03611_),
    .B(_03627_),
    .ZN(_00129_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08803_ (.A1(_03609_),
    .A2(\mem[0][15] ),
    .ZN(_03628_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08804_ (.A1(_03450_),
    .A2(_03611_),
    .B(_03628_),
    .ZN(_00130_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08805_ (.A1(_01430_),
    .A2(net91),
    .ZN(_03629_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _08806_ (.I(_03629_),
    .ZN(_03630_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08807_ (.A1(_01266_),
    .A2(_01358_),
    .ZN(_03631_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _08808_ (.I(_03631_),
    .ZN(_03632_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08809_ (.A1(_03630_),
    .A2(_03632_),
    .ZN(_03633_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08810_ (.I(_03633_),
    .Z(_03634_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08811_ (.I(_03633_),
    .Z(_03635_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08812_ (.A1(_03635_),
    .A2(\mem[10][0] ),
    .ZN(_03636_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08813_ (.A1(_03453_),
    .A2(_03634_),
    .B(_03636_),
    .ZN(_00131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08814_ (.A1(_03635_),
    .A2(\mem[10][1] ),
    .ZN(_03637_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08815_ (.A1(_03462_),
    .A2(_03634_),
    .B(_03637_),
    .ZN(_00132_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08816_ (.A1(_03635_),
    .A2(\mem[10][2] ),
    .ZN(_03638_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08817_ (.A1(_03465_),
    .A2(_03634_),
    .B(_03638_),
    .ZN(_00133_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08818_ (.A1(_03635_),
    .A2(\mem[10][3] ),
    .ZN(_03639_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08819_ (.A1(_03468_),
    .A2(_03634_),
    .B(_03639_),
    .ZN(_00134_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08820_ (.I(_03633_),
    .Z(_03640_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08821_ (.A1(_03640_),
    .A2(\mem[10][4] ),
    .ZN(_03641_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08822_ (.A1(_03471_),
    .A2(_03634_),
    .B(_03641_),
    .ZN(_00135_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08823_ (.A1(_03640_),
    .A2(\mem[10][5] ),
    .ZN(_03642_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08824_ (.A1(_03475_),
    .A2(_03634_),
    .B(_03642_),
    .ZN(_00136_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08825_ (.A1(_03640_),
    .A2(\mem[10][6] ),
    .ZN(_03643_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08826_ (.A1(_03478_),
    .A2(_03634_),
    .B(_03643_),
    .ZN(_00137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08827_ (.A1(_03640_),
    .A2(\mem[10][7] ),
    .ZN(_03644_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08828_ (.A1(_03481_),
    .A2(_03634_),
    .B(_03644_),
    .ZN(_00138_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08829_ (.A1(_03640_),
    .A2(\mem[10][8] ),
    .ZN(_03645_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08830_ (.A1(_03484_),
    .A2(_03634_),
    .B(_03645_),
    .ZN(_00139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08831_ (.A1(_03640_),
    .A2(\mem[10][9] ),
    .ZN(_03646_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08832_ (.A1(_03487_),
    .A2(_03634_),
    .B(_03646_),
    .ZN(_00140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08833_ (.A1(_03640_),
    .A2(\mem[10][10] ),
    .ZN(_03647_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08834_ (.A1(_03490_),
    .A2(_03635_),
    .B(_03647_),
    .ZN(_00141_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08835_ (.A1(_03640_),
    .A2(\mem[10][11] ),
    .ZN(_03648_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08836_ (.A1(_03493_),
    .A2(_03635_),
    .B(_03648_),
    .ZN(_00142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08837_ (.A1(_03640_),
    .A2(\mem[10][12] ),
    .ZN(_03649_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08838_ (.A1(_03496_),
    .A2(_03635_),
    .B(_03649_),
    .ZN(_00143_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08839_ (.A1(_03640_),
    .A2(\mem[10][13] ),
    .ZN(_03650_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08840_ (.A1(_03439_),
    .A2(_03635_),
    .B(_03650_),
    .ZN(_00144_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08841_ (.A1(_03633_),
    .A2(\mem[10][14] ),
    .ZN(_03651_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08842_ (.A1(_03447_),
    .A2(_03635_),
    .B(_03651_),
    .ZN(_00145_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08843_ (.A1(_03633_),
    .A2(\mem[10][15] ),
    .ZN(_03652_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08844_ (.A1(_03450_),
    .A2(_03635_),
    .B(_03652_),
    .ZN(_00146_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08845_ (.A1(_03543_),
    .A2(_01431_),
    .ZN(_03653_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08846_ (.I(_03653_),
    .Z(_03654_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08847_ (.I(_03653_),
    .Z(_03655_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08848_ (.A1(_03655_),
    .A2(\mem[11][0] ),
    .ZN(_03656_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08849_ (.A1(_03453_),
    .A2(_03654_),
    .B(_03656_),
    .ZN(_00147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08850_ (.A1(_03655_),
    .A2(\mem[11][1] ),
    .ZN(_03657_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08851_ (.A1(_03462_),
    .A2(_03654_),
    .B(_03657_),
    .ZN(_00148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08852_ (.A1(_03655_),
    .A2(\mem[11][2] ),
    .ZN(_03658_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08853_ (.A1(_03465_),
    .A2(_03654_),
    .B(_03658_),
    .ZN(_00149_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08854_ (.A1(_03655_),
    .A2(\mem[11][3] ),
    .ZN(_03659_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08855_ (.A1(_03468_),
    .A2(_03654_),
    .B(_03659_),
    .ZN(_00150_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08856_ (.I(_03653_),
    .Z(_03660_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08857_ (.A1(_03660_),
    .A2(\mem[11][4] ),
    .ZN(_03661_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08858_ (.A1(_03471_),
    .A2(_03654_),
    .B(_03661_),
    .ZN(_00151_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08859_ (.A1(_03660_),
    .A2(\mem[11][5] ),
    .ZN(_03662_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08860_ (.A1(_03475_),
    .A2(_03654_),
    .B(_03662_),
    .ZN(_00152_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08861_ (.A1(_03660_),
    .A2(\mem[11][6] ),
    .ZN(_03663_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08862_ (.A1(_03478_),
    .A2(_03654_),
    .B(_03663_),
    .ZN(_00153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08863_ (.A1(_03660_),
    .A2(\mem[11][7] ),
    .ZN(_03664_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08864_ (.A1(_03481_),
    .A2(_03654_),
    .B(_03664_),
    .ZN(_00154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08865_ (.A1(_03660_),
    .A2(\mem[11][8] ),
    .ZN(_03665_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08866_ (.A1(_03484_),
    .A2(_03654_),
    .B(_03665_),
    .ZN(_00155_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08867_ (.A1(_03660_),
    .A2(\mem[11][9] ),
    .ZN(_03666_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08868_ (.A1(_03487_),
    .A2(_03654_),
    .B(_03666_),
    .ZN(_00156_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08869_ (.A1(_03660_),
    .A2(\mem[11][10] ),
    .ZN(_03667_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08870_ (.A1(_03490_),
    .A2(_03655_),
    .B(_03667_),
    .ZN(_00157_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08871_ (.A1(_03660_),
    .A2(\mem[11][11] ),
    .ZN(_03668_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08872_ (.A1(_03493_),
    .A2(_03655_),
    .B(_03668_),
    .ZN(_00158_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08873_ (.A1(_03660_),
    .A2(\mem[11][12] ),
    .ZN(_03669_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08874_ (.A1(_03496_),
    .A2(_03655_),
    .B(_03669_),
    .ZN(_00159_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08875_ (.A1(_03660_),
    .A2(\mem[11][13] ),
    .ZN(_03670_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08876_ (.A1(_03439_),
    .A2(_03655_),
    .B(_03670_),
    .ZN(_00160_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08877_ (.A1(_03653_),
    .A2(\mem[11][14] ),
    .ZN(_03671_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08878_ (.A1(_03447_),
    .A2(_03655_),
    .B(_03671_),
    .ZN(_00161_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08879_ (.A1(_03653_),
    .A2(\mem[11][15] ),
    .ZN(_03672_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08880_ (.A1(_03450_),
    .A2(_03655_),
    .B(_03672_),
    .ZN(_00162_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08881_ (.A1(_03630_),
    .A2(net41),
    .ZN(_03673_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08882_ (.I(_03673_),
    .Z(_03674_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08883_ (.I(_03673_),
    .Z(_03675_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08884_ (.A1(_03675_),
    .A2(\mem[12][0] ),
    .ZN(_03676_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08885_ (.A1(_03453_),
    .A2(_03674_),
    .B(_03676_),
    .ZN(_00163_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08886_ (.A1(_03675_),
    .A2(\mem[12][1] ),
    .ZN(_03677_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08887_ (.A1(_03462_),
    .A2(_03674_),
    .B(_03677_),
    .ZN(_00164_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08888_ (.A1(_03675_),
    .A2(\mem[12][2] ),
    .ZN(_03678_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08889_ (.A1(_03465_),
    .A2(_03674_),
    .B(_03678_),
    .ZN(_00165_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08890_ (.A1(_03675_),
    .A2(\mem[12][3] ),
    .ZN(_03679_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08891_ (.A1(_03468_),
    .A2(_03674_),
    .B(_03679_),
    .ZN(_00166_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08892_ (.I(_03673_),
    .Z(_03680_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08893_ (.A1(_03680_),
    .A2(\mem[12][4] ),
    .ZN(_03681_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08894_ (.A1(_03471_),
    .A2(_03674_),
    .B(_03681_),
    .ZN(_00167_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08895_ (.A1(_03680_),
    .A2(\mem[12][5] ),
    .ZN(_03682_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08896_ (.A1(_03475_),
    .A2(_03674_),
    .B(_03682_),
    .ZN(_00168_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08897_ (.A1(_03680_),
    .A2(\mem[12][6] ),
    .ZN(_03683_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08898_ (.A1(_03478_),
    .A2(_03674_),
    .B(_03683_),
    .ZN(_00169_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08899_ (.A1(_03680_),
    .A2(\mem[12][7] ),
    .ZN(_03684_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08900_ (.A1(_03481_),
    .A2(_03674_),
    .B(_03684_),
    .ZN(_00170_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08901_ (.A1(_03680_),
    .A2(\mem[12][8] ),
    .ZN(_03685_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08902_ (.A1(_03484_),
    .A2(_03674_),
    .B(_03685_),
    .ZN(_00171_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08903_ (.A1(_03680_),
    .A2(\mem[12][9] ),
    .ZN(_03686_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08904_ (.A1(_03487_),
    .A2(_03674_),
    .B(_03686_),
    .ZN(_00172_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08905_ (.A1(_03680_),
    .A2(\mem[12][10] ),
    .ZN(_03687_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08906_ (.A1(_03490_),
    .A2(_03675_),
    .B(_03687_),
    .ZN(_00173_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08907_ (.A1(_03680_),
    .A2(\mem[12][11] ),
    .ZN(_03688_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08908_ (.A1(_03493_),
    .A2(_03675_),
    .B(_03688_),
    .ZN(_00174_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08909_ (.A1(_03680_),
    .A2(\mem[12][12] ),
    .ZN(_03689_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08910_ (.A1(_03496_),
    .A2(_03675_),
    .B(_03689_),
    .ZN(_00175_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08911_ (.I(_03438_),
    .Z(_03690_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08912_ (.A1(_03680_),
    .A2(\mem[12][13] ),
    .ZN(_03691_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08913_ (.A1(_03690_),
    .A2(_03675_),
    .B(_03691_),
    .ZN(_00176_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08914_ (.I(_03446_),
    .Z(_03692_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08915_ (.A1(_03673_),
    .A2(\mem[12][14] ),
    .ZN(_03693_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08916_ (.A1(_03692_),
    .A2(_03675_),
    .B(_03693_),
    .ZN(_00177_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08917_ (.I(_03449_),
    .Z(_03694_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(_03673_),
    .A2(\mem[12][15] ),
    .ZN(_03695_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08919_ (.A1(_03694_),
    .A2(_03675_),
    .B(_03695_),
    .ZN(_00178_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08920_ (.I(_03452_),
    .Z(_03696_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08921_ (.A1(_03630_),
    .A2(_03566_),
    .ZN(_03697_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08922_ (.I(_03697_),
    .Z(_03698_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08923_ (.I(_03697_),
    .Z(_03699_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08924_ (.A1(_03699_),
    .A2(\mem[13][0] ),
    .ZN(_03700_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08925_ (.A1(_03696_),
    .A2(_03698_),
    .B(_03700_),
    .ZN(_00179_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08926_ (.I(_03461_),
    .Z(_03701_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08927_ (.A1(_03699_),
    .A2(\mem[13][1] ),
    .ZN(_03702_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08928_ (.A1(_03701_),
    .A2(_03698_),
    .B(_03702_),
    .ZN(_00180_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08929_ (.I(_03464_),
    .Z(_03703_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08930_ (.A1(_03699_),
    .A2(\mem[13][2] ),
    .ZN(_03704_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08931_ (.A1(_03703_),
    .A2(_03698_),
    .B(_03704_),
    .ZN(_00181_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08932_ (.I(_03467_),
    .Z(_03705_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08933_ (.A1(_03699_),
    .A2(\mem[13][3] ),
    .ZN(_03706_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08934_ (.A1(_03705_),
    .A2(_03698_),
    .B(_03706_),
    .ZN(_00182_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08935_ (.I(_03470_),
    .Z(_03707_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08936_ (.I(_03697_),
    .Z(_03708_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08937_ (.A1(_03708_),
    .A2(\mem[13][4] ),
    .ZN(_03709_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08938_ (.A1(_03707_),
    .A2(_03698_),
    .B(_03709_),
    .ZN(_00183_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08939_ (.I(_03474_),
    .Z(_03710_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08940_ (.A1(_03708_),
    .A2(\mem[13][5] ),
    .ZN(_03711_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08941_ (.A1(_03710_),
    .A2(_03698_),
    .B(_03711_),
    .ZN(_00184_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08942_ (.I(_03477_),
    .Z(_03712_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08943_ (.A1(_03708_),
    .A2(\mem[13][6] ),
    .ZN(_03713_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08944_ (.A1(_03712_),
    .A2(_03698_),
    .B(_03713_),
    .ZN(_00185_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08945_ (.I(_03480_),
    .Z(_03714_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08946_ (.A1(_03708_),
    .A2(\mem[13][7] ),
    .ZN(_03715_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08947_ (.A1(_03714_),
    .A2(_03698_),
    .B(_03715_),
    .ZN(_00186_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08948_ (.I(_03483_),
    .Z(_03716_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08949_ (.A1(_03708_),
    .A2(\mem[13][8] ),
    .ZN(_03717_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08950_ (.A1(_03716_),
    .A2(_03698_),
    .B(_03717_),
    .ZN(_00187_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08951_ (.I(_03486_),
    .Z(_03718_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08952_ (.A1(_03708_),
    .A2(\mem[13][9] ),
    .ZN(_03719_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08953_ (.A1(_03718_),
    .A2(_03698_),
    .B(_03719_),
    .ZN(_00188_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08954_ (.I(_03489_),
    .Z(_03720_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08955_ (.A1(_03708_),
    .A2(\mem[13][10] ),
    .ZN(_03721_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08956_ (.A1(_03720_),
    .A2(_03699_),
    .B(_03721_),
    .ZN(_00189_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08957_ (.I(_03492_),
    .Z(_03722_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08958_ (.A1(_03708_),
    .A2(\mem[13][11] ),
    .ZN(_03723_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08959_ (.A1(_03722_),
    .A2(_03699_),
    .B(_03723_),
    .ZN(_00190_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08960_ (.I(_03495_),
    .Z(_03724_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08961_ (.A1(_03708_),
    .A2(\mem[13][12] ),
    .ZN(_03725_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08962_ (.A1(_03724_),
    .A2(_03699_),
    .B(_03725_),
    .ZN(_00191_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08963_ (.A1(_03708_),
    .A2(\mem[13][13] ),
    .ZN(_03726_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08964_ (.A1(_03690_),
    .A2(_03699_),
    .B(_03726_),
    .ZN(_00192_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08965_ (.A1(_03697_),
    .A2(\mem[13][14] ),
    .ZN(_03727_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08966_ (.A1(_03692_),
    .A2(_03699_),
    .B(_03727_),
    .ZN(_00193_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08967_ (.A1(_03697_),
    .A2(\mem[13][15] ),
    .ZN(_03728_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08968_ (.A1(_03694_),
    .A2(_03699_),
    .B(_03728_),
    .ZN(_00194_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08969_ (.A1(_03630_),
    .A2(_01162_),
    .ZN(_03729_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08970_ (.I(_03729_),
    .Z(_03730_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08971_ (.I(_03729_),
    .Z(_03731_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08972_ (.A1(_03731_),
    .A2(\mem[14][0] ),
    .ZN(_03732_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08973_ (.A1(_03696_),
    .A2(_03730_),
    .B(_03732_),
    .ZN(_00195_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08974_ (.A1(_03731_),
    .A2(\mem[14][1] ),
    .ZN(_03733_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08975_ (.A1(_03701_),
    .A2(_03730_),
    .B(_03733_),
    .ZN(_00196_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08976_ (.A1(_03731_),
    .A2(\mem[14][2] ),
    .ZN(_03734_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08977_ (.A1(_03703_),
    .A2(_03730_),
    .B(_03734_),
    .ZN(_00197_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08978_ (.A1(_03731_),
    .A2(\mem[14][3] ),
    .ZN(_03735_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08979_ (.A1(_03705_),
    .A2(_03730_),
    .B(_03735_),
    .ZN(_00198_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08980_ (.I(_03729_),
    .Z(_03736_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08981_ (.A1(_03736_),
    .A2(\mem[14][4] ),
    .ZN(_03737_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08982_ (.A1(_03707_),
    .A2(_03730_),
    .B(_03737_),
    .ZN(_00199_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08983_ (.A1(_03736_),
    .A2(\mem[14][5] ),
    .ZN(_03738_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08984_ (.A1(_03710_),
    .A2(_03730_),
    .B(_03738_),
    .ZN(_00200_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08985_ (.A1(_03736_),
    .A2(\mem[14][6] ),
    .ZN(_03739_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08986_ (.A1(_03712_),
    .A2(_03730_),
    .B(_03739_),
    .ZN(_00201_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08987_ (.A1(_03736_),
    .A2(\mem[14][7] ),
    .ZN(_03740_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08988_ (.A1(_03714_),
    .A2(_03730_),
    .B(_03740_),
    .ZN(_00202_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08989_ (.A1(_03736_),
    .A2(\mem[14][8] ),
    .ZN(_03741_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08990_ (.A1(_03716_),
    .A2(_03730_),
    .B(_03741_),
    .ZN(_00203_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08991_ (.A1(_03736_),
    .A2(\mem[14][9] ),
    .ZN(_03742_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08992_ (.A1(_03718_),
    .A2(_03730_),
    .B(_03742_),
    .ZN(_00204_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08993_ (.A1(_03736_),
    .A2(\mem[14][10] ),
    .ZN(_03743_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08994_ (.A1(_03720_),
    .A2(_03731_),
    .B(_03743_),
    .ZN(_00205_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08995_ (.A1(_03736_),
    .A2(\mem[14][11] ),
    .ZN(_03744_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08996_ (.A1(_03722_),
    .A2(_03731_),
    .B(_03744_),
    .ZN(_00206_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08997_ (.A1(_03736_),
    .A2(\mem[14][12] ),
    .ZN(_03745_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08998_ (.A1(_03724_),
    .A2(_03731_),
    .B(_03745_),
    .ZN(_00207_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08999_ (.A1(_03736_),
    .A2(\mem[14][13] ),
    .ZN(_03746_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09000_ (.A1(_03690_),
    .A2(_03731_),
    .B(_03746_),
    .ZN(_00208_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09001_ (.A1(_03729_),
    .A2(\mem[14][14] ),
    .ZN(_03747_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09002_ (.A1(_03692_),
    .A2(_03731_),
    .B(_03747_),
    .ZN(_00209_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09003_ (.A1(_03729_),
    .A2(\mem[14][15] ),
    .ZN(_03748_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09004_ (.A1(_03694_),
    .A2(_03731_),
    .B(_03748_),
    .ZN(_00210_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09005_ (.A1(net40),
    .A2(_01431_),
    .ZN(_03749_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09006_ (.I(_03749_),
    .Z(_03750_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09007_ (.I(_03749_),
    .Z(_03751_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09008_ (.A1(_03751_),
    .A2(\mem[15][0] ),
    .ZN(_03752_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09009_ (.A1(_03696_),
    .A2(_03750_),
    .B(_03752_),
    .ZN(_00211_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09010_ (.A1(_03751_),
    .A2(\mem[15][1] ),
    .ZN(_03753_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09011_ (.A1(_03701_),
    .A2(_03750_),
    .B(_03753_),
    .ZN(_00212_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09012_ (.A1(_03751_),
    .A2(\mem[15][2] ),
    .ZN(_03754_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09013_ (.A1(_03703_),
    .A2(_03750_),
    .B(_03754_),
    .ZN(_00213_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09014_ (.A1(_03751_),
    .A2(\mem[15][3] ),
    .ZN(_03755_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09015_ (.A1(_03705_),
    .A2(_03750_),
    .B(_03755_),
    .ZN(_00214_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09016_ (.I(_03749_),
    .Z(_03756_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09017_ (.A1(_03756_),
    .A2(\mem[15][4] ),
    .ZN(_03757_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09018_ (.A1(_03707_),
    .A2(_03750_),
    .B(_03757_),
    .ZN(_00215_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09019_ (.A1(_03756_),
    .A2(\mem[15][5] ),
    .ZN(_03758_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09020_ (.A1(_03710_),
    .A2(_03750_),
    .B(_03758_),
    .ZN(_00216_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09021_ (.A1(_03756_),
    .A2(\mem[15][6] ),
    .ZN(_03759_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09022_ (.A1(_03712_),
    .A2(_03750_),
    .B(_03759_),
    .ZN(_00217_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09023_ (.A1(_03756_),
    .A2(\mem[15][7] ),
    .ZN(_03760_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09024_ (.A1(_03714_),
    .A2(_03750_),
    .B(_03760_),
    .ZN(_00218_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09025_ (.A1(_03756_),
    .A2(\mem[15][8] ),
    .ZN(_03761_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09026_ (.A1(_03716_),
    .A2(_03750_),
    .B(_03761_),
    .ZN(_00219_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09027_ (.A1(_03756_),
    .A2(\mem[15][9] ),
    .ZN(_03762_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09028_ (.A1(_03718_),
    .A2(_03750_),
    .B(_03762_),
    .ZN(_00220_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09029_ (.A1(_03756_),
    .A2(\mem[15][10] ),
    .ZN(_03763_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09030_ (.A1(_03720_),
    .A2(_03751_),
    .B(_03763_),
    .ZN(_00221_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09031_ (.A1(_03756_),
    .A2(\mem[15][11] ),
    .ZN(_03764_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09032_ (.A1(_03722_),
    .A2(_03751_),
    .B(_03764_),
    .ZN(_00222_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09033_ (.A1(_03756_),
    .A2(\mem[15][12] ),
    .ZN(_03765_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09034_ (.A1(_03724_),
    .A2(_03751_),
    .B(_03765_),
    .ZN(_00223_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09035_ (.A1(_03756_),
    .A2(\mem[15][13] ),
    .ZN(_03766_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09036_ (.A1(_03690_),
    .A2(_03751_),
    .B(_03766_),
    .ZN(_00224_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09037_ (.A1(_03749_),
    .A2(\mem[15][14] ),
    .ZN(_03767_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09038_ (.A1(_03692_),
    .A2(_03751_),
    .B(_03767_),
    .ZN(_00225_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09039_ (.A1(_03749_),
    .A2(\mem[15][15] ),
    .ZN(_03768_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09040_ (.A1(_03694_),
    .A2(_03751_),
    .B(_03768_),
    .ZN(_00226_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09041_ (.A1(_03588_),
    .A2(_01082_),
    .ZN(_03769_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09042_ (.I(_03769_),
    .Z(_03770_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09043_ (.I(_03769_),
    .Z(_03771_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09044_ (.A1(_03771_),
    .A2(\mem[16][0] ),
    .ZN(_03772_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09045_ (.A1(_03696_),
    .A2(_03770_),
    .B(_03772_),
    .ZN(_00227_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09046_ (.A1(_03771_),
    .A2(\mem[16][1] ),
    .ZN(_03773_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09047_ (.A1(_03701_),
    .A2(_03770_),
    .B(_03773_),
    .ZN(_00228_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09048_ (.A1(_03771_),
    .A2(\mem[16][2] ),
    .ZN(_03774_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09049_ (.A1(_03703_),
    .A2(_03770_),
    .B(_03774_),
    .ZN(_00229_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09050_ (.A1(_03771_),
    .A2(\mem[16][3] ),
    .ZN(_03775_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09051_ (.A1(_03705_),
    .A2(_03770_),
    .B(_03775_),
    .ZN(_00230_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09052_ (.I(_03769_),
    .Z(_03776_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09053_ (.A1(_03776_),
    .A2(\mem[16][4] ),
    .ZN(_03777_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09054_ (.A1(_03707_),
    .A2(_03770_),
    .B(_03777_),
    .ZN(_00231_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09055_ (.A1(_03776_),
    .A2(\mem[16][5] ),
    .ZN(_03778_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09056_ (.A1(_03710_),
    .A2(_03770_),
    .B(_03778_),
    .ZN(_00232_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09057_ (.A1(_03776_),
    .A2(\mem[16][6] ),
    .ZN(_03779_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09058_ (.A1(_03712_),
    .A2(_03770_),
    .B(_03779_),
    .ZN(_00233_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09059_ (.A1(_03776_),
    .A2(\mem[16][7] ),
    .ZN(_03780_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09060_ (.A1(_03714_),
    .A2(_03770_),
    .B(_03780_),
    .ZN(_00234_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09061_ (.A1(_03776_),
    .A2(\mem[16][8] ),
    .ZN(_03781_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09062_ (.A1(_03716_),
    .A2(_03770_),
    .B(_03781_),
    .ZN(_00235_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09063_ (.A1(_03776_),
    .A2(\mem[16][9] ),
    .ZN(_03782_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09064_ (.A1(_03718_),
    .A2(_03770_),
    .B(_03782_),
    .ZN(_00236_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09065_ (.A1(_03776_),
    .A2(\mem[16][10] ),
    .ZN(_03783_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09066_ (.A1(_03720_),
    .A2(_03771_),
    .B(_03783_),
    .ZN(_00237_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09067_ (.A1(_03776_),
    .A2(\mem[16][11] ),
    .ZN(_03784_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09068_ (.A1(_03722_),
    .A2(_03771_),
    .B(_03784_),
    .ZN(_00238_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09069_ (.A1(_03776_),
    .A2(\mem[16][12] ),
    .ZN(_03785_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09070_ (.A1(_03724_),
    .A2(_03771_),
    .B(_03785_),
    .ZN(_00239_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09071_ (.A1(_03776_),
    .A2(\mem[16][13] ),
    .ZN(_03786_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09072_ (.A1(_03690_),
    .A2(_03771_),
    .B(_03786_),
    .ZN(_00240_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09073_ (.A1(_03769_),
    .A2(\mem[16][14] ),
    .ZN(_03787_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09074_ (.A1(_03692_),
    .A2(_03771_),
    .B(_03787_),
    .ZN(_00241_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09075_ (.A1(_03769_),
    .A2(\mem[16][15] ),
    .ZN(_03788_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09076_ (.A1(_03694_),
    .A2(_03771_),
    .B(_03788_),
    .ZN(_00242_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09077_ (.A1(_01048_),
    .A2(_01043_),
    .A3(net91),
    .ZN(_03789_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _09078_ (.I(net92),
    .ZN(_03790_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09079_ (.A1(net93),
    .A2(_01082_),
    .ZN(_03791_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09080_ (.I(_03791_),
    .Z(_03792_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09081_ (.I(_03791_),
    .Z(_03793_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09082_ (.A1(_03793_),
    .A2(\mem[17][0] ),
    .ZN(_03794_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09083_ (.A1(_03696_),
    .A2(_03792_),
    .B(_03794_),
    .ZN(_00243_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09084_ (.A1(_03793_),
    .A2(\mem[17][1] ),
    .ZN(_03795_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09085_ (.A1(_03701_),
    .A2(_03792_),
    .B(_03795_),
    .ZN(_00244_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09086_ (.A1(_03793_),
    .A2(\mem[17][2] ),
    .ZN(_03796_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09087_ (.A1(_03703_),
    .A2(_03792_),
    .B(_03796_),
    .ZN(_00245_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09088_ (.A1(_03793_),
    .A2(\mem[17][3] ),
    .ZN(_03797_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09089_ (.A1(_03705_),
    .A2(_03792_),
    .B(_03797_),
    .ZN(_00246_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09090_ (.I(_03791_),
    .Z(_03798_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09091_ (.A1(_03798_),
    .A2(\mem[17][4] ),
    .ZN(_03799_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09092_ (.A1(_03707_),
    .A2(_03792_),
    .B(_03799_),
    .ZN(_00247_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09093_ (.A1(_03798_),
    .A2(\mem[17][5] ),
    .ZN(_03800_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09094_ (.A1(_03710_),
    .A2(_03792_),
    .B(_03800_),
    .ZN(_00248_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09095_ (.A1(_03798_),
    .A2(\mem[17][6] ),
    .ZN(_03801_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09096_ (.A1(_03712_),
    .A2(_03792_),
    .B(_03801_),
    .ZN(_00249_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09097_ (.A1(_03798_),
    .A2(\mem[17][7] ),
    .ZN(_03802_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09098_ (.A1(_03714_),
    .A2(_03792_),
    .B(_03802_),
    .ZN(_00250_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09099_ (.A1(_03798_),
    .A2(\mem[17][8] ),
    .ZN(_03803_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09100_ (.A1(_03716_),
    .A2(_03792_),
    .B(_03803_),
    .ZN(_00251_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09101_ (.A1(_03798_),
    .A2(\mem[17][9] ),
    .ZN(_03804_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09102_ (.A1(_03718_),
    .A2(_03792_),
    .B(_03804_),
    .ZN(_00252_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09103_ (.A1(_03798_),
    .A2(\mem[17][10] ),
    .ZN(_03805_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09104_ (.A1(_03720_),
    .A2(_03793_),
    .B(_03805_),
    .ZN(_00253_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09105_ (.A1(_03798_),
    .A2(\mem[17][11] ),
    .ZN(_03806_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09106_ (.A1(_03722_),
    .A2(_03793_),
    .B(_03806_),
    .ZN(_00254_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09107_ (.A1(_03798_),
    .A2(\mem[17][12] ),
    .ZN(_03807_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09108_ (.A1(_03724_),
    .A2(_03793_),
    .B(_03807_),
    .ZN(_00255_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09109_ (.A1(_03798_),
    .A2(\mem[17][13] ),
    .ZN(_03808_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09110_ (.A1(_03690_),
    .A2(_03793_),
    .B(_03808_),
    .ZN(_00256_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09111_ (.A1(_03791_),
    .A2(\mem[17][14] ),
    .ZN(_03809_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09112_ (.A1(_03692_),
    .A2(_03793_),
    .B(_03809_),
    .ZN(_00257_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09113_ (.A1(_03791_),
    .A2(\mem[17][15] ),
    .ZN(_03810_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09114_ (.A1(_03694_),
    .A2(_03793_),
    .B(_03810_),
    .ZN(_00258_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09115_ (.A1(net137),
    .A2(_03440_),
    .ZN(_03811_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09116_ (.A1(_03811_),
    .A2(_03632_),
    .ZN(_03812_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09117_ (.I(_03812_),
    .Z(_03813_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09118_ (.I(_03812_),
    .Z(_03814_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09119_ (.A1(_03814_),
    .A2(\mem[18][0] ),
    .ZN(_03815_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09120_ (.A1(_03696_),
    .A2(_03813_),
    .B(_03815_),
    .ZN(_00259_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09121_ (.A1(_03814_),
    .A2(\mem[18][1] ),
    .ZN(_03816_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09122_ (.A1(_03701_),
    .A2(_03813_),
    .B(_03816_),
    .ZN(_00260_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09123_ (.A1(_03814_),
    .A2(\mem[18][2] ),
    .ZN(_03817_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09124_ (.A1(_03703_),
    .A2(_03813_),
    .B(_03817_),
    .ZN(_00261_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09125_ (.A1(_03814_),
    .A2(\mem[18][3] ),
    .ZN(_03818_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09126_ (.A1(_03705_),
    .A2(_03813_),
    .B(_03818_),
    .ZN(_00262_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09127_ (.I(_03812_),
    .Z(_03819_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09128_ (.A1(_03819_),
    .A2(\mem[18][4] ),
    .ZN(_03820_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09129_ (.A1(_03707_),
    .A2(_03813_),
    .B(_03820_),
    .ZN(_00263_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09130_ (.A1(_03819_),
    .A2(\mem[18][5] ),
    .ZN(_03821_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09131_ (.A1(_03710_),
    .A2(_03813_),
    .B(_03821_),
    .ZN(_00264_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09132_ (.A1(_03819_),
    .A2(\mem[18][6] ),
    .ZN(_03822_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09133_ (.A1(_03712_),
    .A2(_03813_),
    .B(_03822_),
    .ZN(_00265_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09134_ (.A1(_03819_),
    .A2(\mem[18][7] ),
    .ZN(_03823_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09135_ (.A1(_03714_),
    .A2(_03813_),
    .B(_03823_),
    .ZN(_00266_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09136_ (.A1(_03819_),
    .A2(\mem[18][8] ),
    .ZN(_03824_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09137_ (.A1(_03716_),
    .A2(_03813_),
    .B(_03824_),
    .ZN(_00267_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09138_ (.A1(_03819_),
    .A2(\mem[18][9] ),
    .ZN(_03825_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09139_ (.A1(_03718_),
    .A2(_03813_),
    .B(_03825_),
    .ZN(_00268_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09140_ (.A1(_03819_),
    .A2(\mem[18][10] ),
    .ZN(_03826_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09141_ (.A1(_03720_),
    .A2(_03814_),
    .B(_03826_),
    .ZN(_00269_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09142_ (.A1(_03819_),
    .A2(\mem[18][11] ),
    .ZN(_03827_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09143_ (.A1(_03722_),
    .A2(_03814_),
    .B(_03827_),
    .ZN(_00270_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09144_ (.A1(_03819_),
    .A2(\mem[18][12] ),
    .ZN(_03828_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09145_ (.A1(_03724_),
    .A2(_03814_),
    .B(_03828_),
    .ZN(_00271_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09146_ (.A1(_03819_),
    .A2(\mem[18][13] ),
    .ZN(_03829_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09147_ (.A1(_03690_),
    .A2(_03814_),
    .B(_03829_),
    .ZN(_00272_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09148_ (.A1(_03812_),
    .A2(\mem[18][14] ),
    .ZN(_03830_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09149_ (.A1(_03692_),
    .A2(_03814_),
    .B(_03830_),
    .ZN(_00273_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09150_ (.A1(_03812_),
    .A2(\mem[18][15] ),
    .ZN(_03831_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09151_ (.A1(_03694_),
    .A2(_03814_),
    .B(_03831_),
    .ZN(_00274_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09152_ (.A1(net93),
    .A2(_01398_),
    .ZN(_03832_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09153_ (.I(_03832_),
    .Z(_03833_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09154_ (.I(_03832_),
    .Z(_03834_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09155_ (.A1(_03834_),
    .A2(\mem[1][0] ),
    .ZN(_03835_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09156_ (.A1(_03696_),
    .A2(_03833_),
    .B(_03835_),
    .ZN(_00275_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09157_ (.A1(_03834_),
    .A2(\mem[1][1] ),
    .ZN(_03836_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09158_ (.A1(_03701_),
    .A2(_03833_),
    .B(_03836_),
    .ZN(_00276_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09159_ (.A1(_03834_),
    .A2(\mem[1][2] ),
    .ZN(_03837_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09160_ (.A1(_03703_),
    .A2(_03833_),
    .B(_03837_),
    .ZN(_00277_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09161_ (.A1(_03834_),
    .A2(\mem[1][3] ),
    .ZN(_03838_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09162_ (.A1(_03705_),
    .A2(_03833_),
    .B(_03838_),
    .ZN(_00278_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09163_ (.I(_03832_),
    .Z(_03839_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09164_ (.A1(_03839_),
    .A2(\mem[1][4] ),
    .ZN(_03840_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09165_ (.A1(_03707_),
    .A2(_03833_),
    .B(_03840_),
    .ZN(_00279_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09166_ (.A1(_03839_),
    .A2(\mem[1][5] ),
    .ZN(_03841_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09167_ (.A1(_03710_),
    .A2(_03833_),
    .B(_03841_),
    .ZN(_00280_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09168_ (.A1(_03839_),
    .A2(\mem[1][6] ),
    .ZN(_03842_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09169_ (.A1(_03712_),
    .A2(_03833_),
    .B(_03842_),
    .ZN(_00281_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09170_ (.A1(_03839_),
    .A2(\mem[1][7] ),
    .ZN(_03843_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09171_ (.A1(_03714_),
    .A2(_03833_),
    .B(_03843_),
    .ZN(_00282_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09172_ (.A1(_03839_),
    .A2(\mem[1][8] ),
    .ZN(_03844_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09173_ (.A1(_03716_),
    .A2(_03833_),
    .B(_03844_),
    .ZN(_00283_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09174_ (.A1(_03839_),
    .A2(\mem[1][9] ),
    .ZN(_03845_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09175_ (.A1(_03718_),
    .A2(_03833_),
    .B(_03845_),
    .ZN(_00284_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09176_ (.A1(_03839_),
    .A2(\mem[1][10] ),
    .ZN(_03846_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09177_ (.A1(_03720_),
    .A2(_03834_),
    .B(_03846_),
    .ZN(_00285_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09178_ (.A1(_03839_),
    .A2(\mem[1][11] ),
    .ZN(_03847_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09179_ (.A1(_03722_),
    .A2(_03834_),
    .B(_03847_),
    .ZN(_00286_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09180_ (.A1(_03839_),
    .A2(\mem[1][12] ),
    .ZN(_03848_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09181_ (.A1(_03724_),
    .A2(_03834_),
    .B(_03848_),
    .ZN(_00287_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09182_ (.A1(_03839_),
    .A2(\mem[1][13] ),
    .ZN(_03849_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09183_ (.A1(_03690_),
    .A2(_03834_),
    .B(_03849_),
    .ZN(_00288_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09184_ (.A1(_03832_),
    .A2(\mem[1][14] ),
    .ZN(_03850_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09185_ (.A1(_03692_),
    .A2(_03834_),
    .B(_03850_),
    .ZN(_00289_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09186_ (.A1(_03832_),
    .A2(\mem[1][15] ),
    .ZN(_03851_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09187_ (.A1(_03694_),
    .A2(_03834_),
    .B(_03851_),
    .ZN(_00290_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09188_ (.A1(_03811_),
    .A2(net41),
    .ZN(_03852_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09189_ (.I(_03852_),
    .Z(_03853_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09190_ (.I(_03852_),
    .Z(_03854_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09191_ (.A1(_03854_),
    .A2(\mem[20][0] ),
    .ZN(_03855_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09192_ (.A1(_03696_),
    .A2(_03853_),
    .B(_03855_),
    .ZN(_00291_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09193_ (.A1(_03854_),
    .A2(\mem[20][1] ),
    .ZN(_03856_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09194_ (.A1(_03701_),
    .A2(_03853_),
    .B(_03856_),
    .ZN(_00292_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09195_ (.A1(_03854_),
    .A2(\mem[20][2] ),
    .ZN(_03857_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09196_ (.A1(_03703_),
    .A2(_03853_),
    .B(_03857_),
    .ZN(_00293_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09197_ (.A1(_03854_),
    .A2(\mem[20][3] ),
    .ZN(_03858_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09198_ (.A1(_03705_),
    .A2(_03853_),
    .B(_03858_),
    .ZN(_00294_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09199_ (.I(_03852_),
    .Z(_03859_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09200_ (.A1(_03859_),
    .A2(\mem[20][4] ),
    .ZN(_03860_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09201_ (.A1(_03707_),
    .A2(_03853_),
    .B(_03860_),
    .ZN(_00295_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09202_ (.A1(_03859_),
    .A2(\mem[20][5] ),
    .ZN(_03861_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09203_ (.A1(_03710_),
    .A2(_03853_),
    .B(_03861_),
    .ZN(_00296_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09204_ (.A1(_03859_),
    .A2(\mem[20][6] ),
    .ZN(_03862_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09205_ (.A1(_03712_),
    .A2(_03853_),
    .B(_03862_),
    .ZN(_00297_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09206_ (.A1(_03859_),
    .A2(\mem[20][7] ),
    .ZN(_03863_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09207_ (.A1(_03714_),
    .A2(_03853_),
    .B(_03863_),
    .ZN(_00298_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09208_ (.A1(_03859_),
    .A2(\mem[20][8] ),
    .ZN(_03864_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09209_ (.A1(_03716_),
    .A2(_03853_),
    .B(_03864_),
    .ZN(_00299_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09210_ (.A1(_03859_),
    .A2(\mem[20][9] ),
    .ZN(_03865_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09211_ (.A1(_03718_),
    .A2(_03853_),
    .B(_03865_),
    .ZN(_00300_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09212_ (.A1(_03859_),
    .A2(\mem[20][10] ),
    .ZN(_03866_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09213_ (.A1(_03720_),
    .A2(_03854_),
    .B(_03866_),
    .ZN(_00301_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09214_ (.A1(_03859_),
    .A2(\mem[20][11] ),
    .ZN(_03867_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09215_ (.A1(_03722_),
    .A2(_03854_),
    .B(_03867_),
    .ZN(_00302_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09216_ (.A1(_03859_),
    .A2(\mem[20][12] ),
    .ZN(_03868_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09217_ (.A1(_03724_),
    .A2(_03854_),
    .B(_03868_),
    .ZN(_00303_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09218_ (.A1(_03859_),
    .A2(\mem[20][13] ),
    .ZN(_03869_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09219_ (.A1(_03690_),
    .A2(_03854_),
    .B(_03869_),
    .ZN(_00304_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09220_ (.A1(_03852_),
    .A2(\mem[20][14] ),
    .ZN(_03870_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09221_ (.A1(_03692_),
    .A2(_03854_),
    .B(_03870_),
    .ZN(_00305_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09222_ (.A1(_03852_),
    .A2(\mem[20][15] ),
    .ZN(_03871_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09223_ (.A1(_03694_),
    .A2(_03854_),
    .B(_03871_),
    .ZN(_00306_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09224_ (.A1(_03811_),
    .A2(_03566_),
    .ZN(_03872_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09225_ (.I(_03872_),
    .Z(_03873_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09226_ (.I(_03872_),
    .Z(_03874_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09227_ (.A1(_03874_),
    .A2(\mem[21][0] ),
    .ZN(_03875_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09228_ (.A1(_03696_),
    .A2(_03873_),
    .B(_03875_),
    .ZN(_00307_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09229_ (.A1(_03874_),
    .A2(\mem[21][1] ),
    .ZN(_03876_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09230_ (.A1(_03701_),
    .A2(_03873_),
    .B(_03876_),
    .ZN(_00308_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09231_ (.A1(_03874_),
    .A2(\mem[21][2] ),
    .ZN(_03877_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09232_ (.A1(_03703_),
    .A2(_03873_),
    .B(_03877_),
    .ZN(_00309_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09233_ (.A1(_03874_),
    .A2(\mem[21][3] ),
    .ZN(_03878_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09234_ (.A1(_03705_),
    .A2(_03873_),
    .B(_03878_),
    .ZN(_00310_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09235_ (.I(_03872_),
    .Z(_03879_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09236_ (.A1(_03879_),
    .A2(\mem[21][4] ),
    .ZN(_03880_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09237_ (.A1(_03707_),
    .A2(_03873_),
    .B(_03880_),
    .ZN(_00311_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09238_ (.A1(_03879_),
    .A2(\mem[21][5] ),
    .ZN(_03881_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09239_ (.A1(_03710_),
    .A2(_03873_),
    .B(_03881_),
    .ZN(_00312_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09240_ (.A1(_03879_),
    .A2(\mem[21][6] ),
    .ZN(_03882_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09241_ (.A1(_03712_),
    .A2(_03873_),
    .B(_03882_),
    .ZN(_00313_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09242_ (.A1(_03879_),
    .A2(\mem[21][7] ),
    .ZN(_03883_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09243_ (.A1(_03714_),
    .A2(_03873_),
    .B(_03883_),
    .ZN(_00314_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09244_ (.A1(_03879_),
    .A2(\mem[21][8] ),
    .ZN(_03884_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09245_ (.A1(_03716_),
    .A2(_03873_),
    .B(_03884_),
    .ZN(_00315_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09246_ (.A1(_03879_),
    .A2(\mem[21][9] ),
    .ZN(_03885_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09247_ (.A1(_03718_),
    .A2(_03873_),
    .B(_03885_),
    .ZN(_00316_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09248_ (.A1(_03879_),
    .A2(\mem[21][10] ),
    .ZN(_03886_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09249_ (.A1(_03720_),
    .A2(_03874_),
    .B(_03886_),
    .ZN(_00317_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09250_ (.A1(_03879_),
    .A2(\mem[21][11] ),
    .ZN(_03887_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09251_ (.A1(_03722_),
    .A2(_03874_),
    .B(_03887_),
    .ZN(_00318_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09252_ (.A1(_03879_),
    .A2(\mem[21][12] ),
    .ZN(_03888_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09253_ (.A1(_03724_),
    .A2(_03874_),
    .B(_03888_),
    .ZN(_00319_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09254_ (.A1(_03879_),
    .A2(\mem[21][13] ),
    .ZN(_03889_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09255_ (.A1(_03690_),
    .A2(_03874_),
    .B(_03889_),
    .ZN(_00320_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09256_ (.A1(_03872_),
    .A2(\mem[21][14] ),
    .ZN(_03890_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09257_ (.A1(_03692_),
    .A2(_03874_),
    .B(_03890_),
    .ZN(_00321_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09258_ (.A1(_03872_),
    .A2(\mem[21][15] ),
    .ZN(_03891_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09259_ (.A1(_03694_),
    .A2(_03874_),
    .B(_03891_),
    .ZN(_00322_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09260_ (.A1(_03811_),
    .A2(_01162_),
    .ZN(_03892_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09261_ (.I(_03892_),
    .Z(_03893_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09262_ (.I(_03892_),
    .Z(_03894_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09263_ (.A1(_03894_),
    .A2(\mem[22][0] ),
    .ZN(_03895_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09264_ (.A1(_03696_),
    .A2(_03893_),
    .B(_03895_),
    .ZN(_00323_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09265_ (.A1(_03894_),
    .A2(\mem[22][1] ),
    .ZN(_03896_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09266_ (.A1(_03701_),
    .A2(_03893_),
    .B(_03896_),
    .ZN(_00324_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09267_ (.A1(_03894_),
    .A2(\mem[22][2] ),
    .ZN(_03897_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09268_ (.A1(_03703_),
    .A2(_03893_),
    .B(_03897_),
    .ZN(_00325_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09269_ (.A1(_03894_),
    .A2(\mem[22][3] ),
    .ZN(_03898_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09270_ (.A1(_03705_),
    .A2(_03893_),
    .B(_03898_),
    .ZN(_00326_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09271_ (.I(_03892_),
    .Z(_03899_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09272_ (.A1(_03899_),
    .A2(\mem[22][4] ),
    .ZN(_03900_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09273_ (.A1(_03707_),
    .A2(_03893_),
    .B(_03900_),
    .ZN(_00327_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09274_ (.A1(_03899_),
    .A2(\mem[22][5] ),
    .ZN(_03901_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09275_ (.A1(_03710_),
    .A2(_03893_),
    .B(_03901_),
    .ZN(_00328_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09276_ (.A1(_03899_),
    .A2(\mem[22][6] ),
    .ZN(_03902_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09277_ (.A1(_03712_),
    .A2(_03893_),
    .B(_03902_),
    .ZN(_00329_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09278_ (.A1(_03899_),
    .A2(\mem[22][7] ),
    .ZN(_03903_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09279_ (.A1(_03714_),
    .A2(_03893_),
    .B(_03903_),
    .ZN(_00330_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09280_ (.A1(_03899_),
    .A2(\mem[22][8] ),
    .ZN(_03904_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09281_ (.A1(_03716_),
    .A2(_03893_),
    .B(_03904_),
    .ZN(_00331_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09282_ (.A1(_03899_),
    .A2(\mem[22][9] ),
    .ZN(_03905_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09283_ (.A1(_03718_),
    .A2(_03893_),
    .B(_03905_),
    .ZN(_00332_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09284_ (.A1(_03899_),
    .A2(\mem[22][10] ),
    .ZN(_03906_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09285_ (.A1(_03720_),
    .A2(_03894_),
    .B(_03906_),
    .ZN(_00333_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09286_ (.A1(_03899_),
    .A2(\mem[22][11] ),
    .ZN(_03907_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09287_ (.A1(_03722_),
    .A2(_03894_),
    .B(_03907_),
    .ZN(_00334_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09288_ (.A1(_03899_),
    .A2(\mem[22][12] ),
    .ZN(_03908_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09289_ (.A1(_03724_),
    .A2(_03894_),
    .B(_03908_),
    .ZN(_00335_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09290_ (.I(_03438_),
    .Z(_03909_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09291_ (.A1(_03899_),
    .A2(\mem[22][13] ),
    .ZN(_03910_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09292_ (.A1(_03909_),
    .A2(_03894_),
    .B(_03910_),
    .ZN(_00336_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09293_ (.I(_03446_),
    .Z(_03911_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09294_ (.A1(_03892_),
    .A2(\mem[22][14] ),
    .ZN(_03912_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09295_ (.A1(_03911_),
    .A2(_03894_),
    .B(_03912_),
    .ZN(_00337_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09296_ (.I(_03449_),
    .Z(_03913_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09297_ (.A1(_03892_),
    .A2(\mem[22][15] ),
    .ZN(_03914_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09298_ (.A1(_03913_),
    .A2(_03894_),
    .B(_03914_),
    .ZN(_00338_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09299_ (.I(_03452_),
    .Z(_03915_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09300_ (.A1(net40),
    .A2(_01081_),
    .ZN(_03916_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09301_ (.I(_03916_),
    .Z(_03917_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09302_ (.I(_03916_),
    .Z(_03918_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09303_ (.A1(_03918_),
    .A2(\mem[23][0] ),
    .ZN(_03919_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09304_ (.A1(_03915_),
    .A2(_03917_),
    .B(_03919_),
    .ZN(_00339_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09305_ (.I(_03461_),
    .Z(_03920_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09306_ (.A1(_03918_),
    .A2(\mem[23][1] ),
    .ZN(_03921_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09307_ (.A1(_03920_),
    .A2(_03917_),
    .B(_03921_),
    .ZN(_00340_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09308_ (.I(_03464_),
    .Z(_03922_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09309_ (.A1(_03918_),
    .A2(\mem[23][2] ),
    .ZN(_03923_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09310_ (.A1(_03922_),
    .A2(_03917_),
    .B(_03923_),
    .ZN(_00341_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09311_ (.I(_03467_),
    .Z(_03924_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09312_ (.A1(_03918_),
    .A2(\mem[23][3] ),
    .ZN(_03925_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09313_ (.A1(_03924_),
    .A2(_03917_),
    .B(_03925_),
    .ZN(_00342_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09314_ (.I(_03470_),
    .Z(_03926_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09315_ (.I(_03916_),
    .Z(_03927_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09316_ (.A1(_03927_),
    .A2(\mem[23][4] ),
    .ZN(_03928_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09317_ (.A1(_03926_),
    .A2(_03917_),
    .B(_03928_),
    .ZN(_00343_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09318_ (.I(_03474_),
    .Z(_03929_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09319_ (.A1(_03927_),
    .A2(\mem[23][5] ),
    .ZN(_03930_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09320_ (.A1(_03929_),
    .A2(_03917_),
    .B(_03930_),
    .ZN(_00344_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09321_ (.I(_03477_),
    .Z(_03931_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09322_ (.A1(_03927_),
    .A2(\mem[23][6] ),
    .ZN(_03932_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09323_ (.A1(_03931_),
    .A2(_03917_),
    .B(_03932_),
    .ZN(_00345_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09324_ (.I(_03480_),
    .Z(_03933_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09325_ (.A1(_03927_),
    .A2(\mem[23][7] ),
    .ZN(_03934_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09326_ (.A1(_03933_),
    .A2(_03917_),
    .B(_03934_),
    .ZN(_00346_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09327_ (.I(_03483_),
    .Z(_03935_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09328_ (.A1(_03927_),
    .A2(\mem[23][8] ),
    .ZN(_03936_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09329_ (.A1(_03935_),
    .A2(_03917_),
    .B(_03936_),
    .ZN(_00347_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09330_ (.I(_03486_),
    .Z(_03937_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09331_ (.A1(_03927_),
    .A2(\mem[23][9] ),
    .ZN(_03938_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09332_ (.A1(_03937_),
    .A2(_03917_),
    .B(_03938_),
    .ZN(_00348_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09333_ (.I(_03489_),
    .Z(_03939_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09334_ (.A1(_03927_),
    .A2(\mem[23][10] ),
    .ZN(_03940_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09335_ (.A1(_03939_),
    .A2(_03918_),
    .B(_03940_),
    .ZN(_00349_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09336_ (.I(_03492_),
    .Z(_03941_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09337_ (.A1(_03927_),
    .A2(\mem[23][11] ),
    .ZN(_03942_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09338_ (.A1(_03941_),
    .A2(_03918_),
    .B(_03942_),
    .ZN(_00350_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09339_ (.I(_03495_),
    .Z(_03943_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09340_ (.A1(_03927_),
    .A2(\mem[23][12] ),
    .ZN(_03944_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09341_ (.A1(_03943_),
    .A2(_03918_),
    .B(_03944_),
    .ZN(_00351_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09342_ (.A1(_03927_),
    .A2(\mem[23][13] ),
    .ZN(_03945_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09343_ (.A1(_03909_),
    .A2(_03918_),
    .B(_03945_),
    .ZN(_00352_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09344_ (.A1(_03916_),
    .A2(\mem[23][14] ),
    .ZN(_03946_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09345_ (.A1(_03911_),
    .A2(_03918_),
    .B(_03946_),
    .ZN(_00353_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09346_ (.A1(_03916_),
    .A2(\mem[23][15] ),
    .ZN(_03947_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09347_ (.A1(_03913_),
    .A2(_03918_),
    .B(_03947_),
    .ZN(_00354_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09348_ (.A1(_03588_),
    .A2(_01104_),
    .ZN(_03948_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09349_ (.I(_03948_),
    .Z(_03949_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09350_ (.I(_03948_),
    .Z(_03950_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09351_ (.A1(_03950_),
    .A2(\mem[24][0] ),
    .ZN(_03951_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09352_ (.A1(_03915_),
    .A2(_03949_),
    .B(_03951_),
    .ZN(_00355_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09353_ (.A1(_03950_),
    .A2(\mem[24][1] ),
    .ZN(_03952_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09354_ (.A1(_03920_),
    .A2(_03949_),
    .B(_03952_),
    .ZN(_00356_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09355_ (.A1(_03950_),
    .A2(\mem[24][2] ),
    .ZN(_03953_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09356_ (.A1(_03922_),
    .A2(_03949_),
    .B(_03953_),
    .ZN(_00357_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09357_ (.A1(_03950_),
    .A2(\mem[24][3] ),
    .ZN(_03954_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09358_ (.A1(_03924_),
    .A2(_03949_),
    .B(_03954_),
    .ZN(_00358_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09359_ (.I(_03948_),
    .Z(_03955_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09360_ (.A1(_03955_),
    .A2(\mem[24][4] ),
    .ZN(_03956_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09361_ (.A1(_03926_),
    .A2(_03949_),
    .B(_03956_),
    .ZN(_00359_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09362_ (.A1(_03955_),
    .A2(\mem[24][5] ),
    .ZN(_03957_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09363_ (.A1(_03929_),
    .A2(_03949_),
    .B(_03957_),
    .ZN(_00360_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09364_ (.A1(_03955_),
    .A2(\mem[24][6] ),
    .ZN(_03958_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09365_ (.A1(_03931_),
    .A2(_03949_),
    .B(_03958_),
    .ZN(_00361_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09366_ (.A1(_03955_),
    .A2(\mem[24][7] ),
    .ZN(_03959_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09367_ (.A1(_03933_),
    .A2(_03949_),
    .B(_03959_),
    .ZN(_00362_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09368_ (.A1(_03955_),
    .A2(\mem[24][8] ),
    .ZN(_03960_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09369_ (.A1(_03935_),
    .A2(_03949_),
    .B(_03960_),
    .ZN(_00363_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09370_ (.A1(_03955_),
    .A2(\mem[24][9] ),
    .ZN(_03961_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09371_ (.A1(_03937_),
    .A2(_03949_),
    .B(_03961_),
    .ZN(_00364_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09372_ (.A1(_03955_),
    .A2(\mem[24][10] ),
    .ZN(_03962_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09373_ (.A1(_03939_),
    .A2(_03950_),
    .B(_03962_),
    .ZN(_00365_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09374_ (.A1(_03955_),
    .A2(\mem[24][11] ),
    .ZN(_03963_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09375_ (.A1(_03941_),
    .A2(_03950_),
    .B(_03963_),
    .ZN(_00366_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09376_ (.A1(_03955_),
    .A2(\mem[24][12] ),
    .ZN(_03964_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09377_ (.A1(_03943_),
    .A2(_03950_),
    .B(_03964_),
    .ZN(_00367_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09378_ (.A1(_03955_),
    .A2(\mem[24][13] ),
    .ZN(_03965_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09379_ (.A1(_03909_),
    .A2(_03950_),
    .B(_03965_),
    .ZN(_00368_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09380_ (.A1(_03948_),
    .A2(\mem[24][14] ),
    .ZN(_03966_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09381_ (.A1(_03911_),
    .A2(_03950_),
    .B(_03966_),
    .ZN(_00369_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09382_ (.A1(_03948_),
    .A2(\mem[24][15] ),
    .ZN(_03967_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09383_ (.A1(_03913_),
    .A2(_03950_),
    .B(_03967_),
    .ZN(_00370_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09384_ (.A1(net93),
    .A2(_01104_),
    .ZN(_03968_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09385_ (.I(_03968_),
    .Z(_03969_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09386_ (.I(_03968_),
    .Z(_03970_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09387_ (.A1(_03970_),
    .A2(\mem[25][0] ),
    .ZN(_03971_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09388_ (.A1(_03915_),
    .A2(_03969_),
    .B(_03971_),
    .ZN(_00371_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09389_ (.A1(_03970_),
    .A2(\mem[25][1] ),
    .ZN(_03972_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09390_ (.A1(_03920_),
    .A2(_03969_),
    .B(_03972_),
    .ZN(_00372_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09391_ (.A1(_03970_),
    .A2(\mem[25][2] ),
    .ZN(_03973_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09392_ (.A1(_03922_),
    .A2(_03969_),
    .B(_03973_),
    .ZN(_00373_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09393_ (.A1(_03970_),
    .A2(\mem[25][3] ),
    .ZN(_03974_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09394_ (.A1(_03924_),
    .A2(_03969_),
    .B(_03974_),
    .ZN(_00374_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09395_ (.I(_03968_),
    .Z(_03975_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09396_ (.A1(_03975_),
    .A2(\mem[25][4] ),
    .ZN(_03976_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09397_ (.A1(_03926_),
    .A2(_03969_),
    .B(_03976_),
    .ZN(_00375_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09398_ (.A1(_03975_),
    .A2(\mem[25][5] ),
    .ZN(_03977_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09399_ (.A1(_03929_),
    .A2(_03969_),
    .B(_03977_),
    .ZN(_00376_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09400_ (.A1(_03975_),
    .A2(\mem[25][6] ),
    .ZN(_03978_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09401_ (.A1(_03931_),
    .A2(_03969_),
    .B(_03978_),
    .ZN(_00377_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09402_ (.A1(_03975_),
    .A2(\mem[25][7] ),
    .ZN(_03979_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09403_ (.A1(_03933_),
    .A2(_03969_),
    .B(_03979_),
    .ZN(_00378_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09404_ (.A1(_03975_),
    .A2(\mem[25][8] ),
    .ZN(_03980_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09405_ (.A1(_03935_),
    .A2(_03969_),
    .B(_03980_),
    .ZN(_00379_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09406_ (.A1(_03975_),
    .A2(\mem[25][9] ),
    .ZN(_03981_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09407_ (.A1(_03937_),
    .A2(_03969_),
    .B(_03981_),
    .ZN(_00380_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09408_ (.A1(_03975_),
    .A2(\mem[25][10] ),
    .ZN(_03982_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09409_ (.A1(_03939_),
    .A2(_03970_),
    .B(_03982_),
    .ZN(_00381_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09410_ (.A1(_03975_),
    .A2(\mem[25][11] ),
    .ZN(_03983_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09411_ (.A1(_03941_),
    .A2(_03970_),
    .B(_03983_),
    .ZN(_00382_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09412_ (.A1(_03975_),
    .A2(\mem[25][12] ),
    .ZN(_03984_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09413_ (.A1(_03943_),
    .A2(_03970_),
    .B(_03984_),
    .ZN(_00383_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09414_ (.A1(_03975_),
    .A2(\mem[25][13] ),
    .ZN(_03985_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09415_ (.A1(_03909_),
    .A2(_03970_),
    .B(_03985_),
    .ZN(_00384_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09416_ (.A1(_03968_),
    .A2(\mem[25][14] ),
    .ZN(_03986_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09417_ (.A1(_03911_),
    .A2(_03970_),
    .B(_03986_),
    .ZN(_00385_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09418_ (.A1(_03968_),
    .A2(\mem[25][15] ),
    .ZN(_03987_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09419_ (.A1(_03913_),
    .A2(_03970_),
    .B(_03987_),
    .ZN(_00386_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09420_ (.A1(net119),
    .A2(_03632_),
    .ZN(_03988_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09421_ (.I(_03988_),
    .Z(_03989_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09422_ (.I(_03988_),
    .Z(_03990_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09423_ (.A1(_03990_),
    .A2(\mem[26][0] ),
    .ZN(_03991_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09424_ (.A1(_03915_),
    .A2(_03989_),
    .B(_03991_),
    .ZN(_00387_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09425_ (.A1(_03990_),
    .A2(\mem[26][1] ),
    .ZN(_03992_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09426_ (.A1(_03920_),
    .A2(_03989_),
    .B(_03992_),
    .ZN(_00388_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09427_ (.A1(_03990_),
    .A2(\mem[26][2] ),
    .ZN(_03993_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09428_ (.A1(_03922_),
    .A2(_03989_),
    .B(_03993_),
    .ZN(_00389_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09429_ (.A1(_03990_),
    .A2(\mem[26][3] ),
    .ZN(_03994_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09430_ (.A1(_03924_),
    .A2(_03989_),
    .B(_03994_),
    .ZN(_00390_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09431_ (.I(_03988_),
    .Z(_03995_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09432_ (.A1(_03995_),
    .A2(\mem[26][4] ),
    .ZN(_03996_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09433_ (.A1(_03926_),
    .A2(_03989_),
    .B(_03996_),
    .ZN(_00391_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09434_ (.A1(_03995_),
    .A2(\mem[26][5] ),
    .ZN(_03997_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09435_ (.A1(_03929_),
    .A2(_03989_),
    .B(_03997_),
    .ZN(_00392_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09436_ (.A1(_03995_),
    .A2(\mem[26][6] ),
    .ZN(_03998_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09437_ (.A1(_03931_),
    .A2(_03989_),
    .B(_03998_),
    .ZN(_00393_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09438_ (.A1(_03995_),
    .A2(\mem[26][7] ),
    .ZN(_03999_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09439_ (.A1(_03933_),
    .A2(_03989_),
    .B(_03999_),
    .ZN(_00394_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09440_ (.A1(_03995_),
    .A2(\mem[26][8] ),
    .ZN(_04000_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09441_ (.A1(_03935_),
    .A2(_03989_),
    .B(_04000_),
    .ZN(_00395_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09442_ (.A1(_03995_),
    .A2(\mem[26][9] ),
    .ZN(_04001_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09443_ (.A1(_03937_),
    .A2(_03989_),
    .B(_04001_),
    .ZN(_00396_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09444_ (.A1(_03995_),
    .A2(\mem[26][10] ),
    .ZN(_04002_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09445_ (.A1(_03939_),
    .A2(_03990_),
    .B(_04002_),
    .ZN(_00397_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09446_ (.A1(_03995_),
    .A2(\mem[26][11] ),
    .ZN(_04003_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09447_ (.A1(_03941_),
    .A2(_03990_),
    .B(_04003_),
    .ZN(_00398_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09448_ (.A1(_03995_),
    .A2(\mem[26][12] ),
    .ZN(_04004_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09449_ (.A1(_03943_),
    .A2(_03990_),
    .B(_04004_),
    .ZN(_00399_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09450_ (.A1(_03995_),
    .A2(\mem[26][13] ),
    .ZN(_04005_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09451_ (.A1(_03909_),
    .A2(_03990_),
    .B(_04005_),
    .ZN(_00400_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09452_ (.A1(_03988_),
    .A2(\mem[26][14] ),
    .ZN(_04006_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09453_ (.A1(_03911_),
    .A2(_03990_),
    .B(_04006_),
    .ZN(_00401_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09454_ (.A1(_03988_),
    .A2(\mem[26][15] ),
    .ZN(_04007_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09455_ (.A1(_03913_),
    .A2(_03990_),
    .B(_04007_),
    .ZN(_00402_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09456_ (.A1(_03543_),
    .A2(_01104_),
    .ZN(_04008_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09457_ (.I(_04008_),
    .Z(_04009_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09458_ (.I(_04008_),
    .Z(_04010_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09459_ (.A1(_04010_),
    .A2(\mem[27][0] ),
    .ZN(_04011_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09460_ (.A1(_03915_),
    .A2(_04009_),
    .B(_04011_),
    .ZN(_00403_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09461_ (.A1(_04010_),
    .A2(\mem[27][1] ),
    .ZN(_04012_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09462_ (.A1(_03920_),
    .A2(_04009_),
    .B(_04012_),
    .ZN(_00404_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09463_ (.A1(_04010_),
    .A2(\mem[27][2] ),
    .ZN(_04013_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09464_ (.A1(_03922_),
    .A2(_04009_),
    .B(_04013_),
    .ZN(_00405_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09465_ (.A1(_04010_),
    .A2(\mem[27][3] ),
    .ZN(_04014_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09466_ (.A1(_03924_),
    .A2(_04009_),
    .B(_04014_),
    .ZN(_00406_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09467_ (.I(_04008_),
    .Z(_04015_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09468_ (.A1(_04015_),
    .A2(\mem[27][4] ),
    .ZN(_04016_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09469_ (.A1(_03926_),
    .A2(_04009_),
    .B(_04016_),
    .ZN(_00407_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09470_ (.A1(_04015_),
    .A2(\mem[27][5] ),
    .ZN(_04017_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09471_ (.A1(_03929_),
    .A2(_04009_),
    .B(_04017_),
    .ZN(_00408_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09472_ (.A1(_04015_),
    .A2(\mem[27][6] ),
    .ZN(_04018_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09473_ (.A1(_03931_),
    .A2(_04009_),
    .B(_04018_),
    .ZN(_00409_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09474_ (.A1(_04015_),
    .A2(\mem[27][7] ),
    .ZN(_04019_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09475_ (.A1(_03933_),
    .A2(_04009_),
    .B(_04019_),
    .ZN(_00410_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09476_ (.A1(_04015_),
    .A2(\mem[27][8] ),
    .ZN(_04020_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09477_ (.A1(_03935_),
    .A2(_04009_),
    .B(_04020_),
    .ZN(_00411_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09478_ (.A1(_04015_),
    .A2(\mem[27][9] ),
    .ZN(_04021_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09479_ (.A1(_03937_),
    .A2(_04009_),
    .B(_04021_),
    .ZN(_00412_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09480_ (.A1(_04015_),
    .A2(\mem[27][10] ),
    .ZN(_04022_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09481_ (.A1(_03939_),
    .A2(_04010_),
    .B(_04022_),
    .ZN(_00413_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09482_ (.A1(_04015_),
    .A2(\mem[27][11] ),
    .ZN(_04023_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09483_ (.A1(_03941_),
    .A2(_04010_),
    .B(_04023_),
    .ZN(_00414_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09484_ (.A1(_04015_),
    .A2(\mem[27][12] ),
    .ZN(_04024_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09485_ (.A1(_03943_),
    .A2(_04010_),
    .B(_04024_),
    .ZN(_00415_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09486_ (.A1(_04015_),
    .A2(\mem[27][13] ),
    .ZN(_04025_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09487_ (.A1(_03909_),
    .A2(_04010_),
    .B(_04025_),
    .ZN(_00416_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09488_ (.A1(_04008_),
    .A2(\mem[27][14] ),
    .ZN(_04026_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09489_ (.A1(_03911_),
    .A2(_04010_),
    .B(_04026_),
    .ZN(_00417_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09490_ (.A1(_04008_),
    .A2(\mem[27][15] ),
    .ZN(_04027_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09491_ (.A1(_03913_),
    .A2(_04010_),
    .B(_04027_),
    .ZN(_00418_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09492_ (.A1(net119),
    .A2(net132),
    .ZN(_04028_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09493_ (.I(_04028_),
    .Z(_04029_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09494_ (.I(_04028_),
    .Z(_04030_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09495_ (.A1(_04030_),
    .A2(\mem[28][0] ),
    .ZN(_04031_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09496_ (.A1(_03915_),
    .A2(_04029_),
    .B(_04031_),
    .ZN(_00419_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09497_ (.A1(_04030_),
    .A2(\mem[28][1] ),
    .ZN(_04032_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09498_ (.A1(_03920_),
    .A2(_04029_),
    .B(_04032_),
    .ZN(_00420_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09499_ (.A1(_04030_),
    .A2(\mem[28][2] ),
    .ZN(_04033_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09500_ (.A1(_03922_),
    .A2(_04029_),
    .B(_04033_),
    .ZN(_00421_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09501_ (.A1(_04030_),
    .A2(\mem[28][3] ),
    .ZN(_04034_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09502_ (.A1(_03924_),
    .A2(_04029_),
    .B(_04034_),
    .ZN(_00422_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09503_ (.I(_04028_),
    .Z(_04035_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09504_ (.A1(_04035_),
    .A2(\mem[28][4] ),
    .ZN(_04036_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09505_ (.A1(_03926_),
    .A2(_04029_),
    .B(_04036_),
    .ZN(_00423_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09506_ (.A1(_04035_),
    .A2(\mem[28][5] ),
    .ZN(_04037_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09507_ (.A1(_03929_),
    .A2(_04029_),
    .B(_04037_),
    .ZN(_00424_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09508_ (.A1(_04035_),
    .A2(\mem[28][6] ),
    .ZN(_04038_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09509_ (.A1(_03931_),
    .A2(_04029_),
    .B(_04038_),
    .ZN(_00425_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09510_ (.A1(_04035_),
    .A2(\mem[28][7] ),
    .ZN(_04039_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09511_ (.A1(_03933_),
    .A2(_04029_),
    .B(_04039_),
    .ZN(_00426_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09512_ (.A1(_04035_),
    .A2(\mem[28][8] ),
    .ZN(_04040_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09513_ (.A1(_03935_),
    .A2(_04029_),
    .B(_04040_),
    .ZN(_00427_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09514_ (.A1(_04035_),
    .A2(\mem[28][9] ),
    .ZN(_04041_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09515_ (.A1(_03937_),
    .A2(_04029_),
    .B(_04041_),
    .ZN(_00428_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09516_ (.A1(_04035_),
    .A2(\mem[28][10] ),
    .ZN(_04042_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09517_ (.A1(_03939_),
    .A2(_04030_),
    .B(_04042_),
    .ZN(_00429_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09518_ (.A1(_04035_),
    .A2(\mem[28][11] ),
    .ZN(_04043_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09519_ (.A1(_03941_),
    .A2(_04030_),
    .B(_04043_),
    .ZN(_00430_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09520_ (.A1(_04035_),
    .A2(\mem[28][12] ),
    .ZN(_04044_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09521_ (.A1(_03943_),
    .A2(_04030_),
    .B(_04044_),
    .ZN(_00431_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09522_ (.A1(_04035_),
    .A2(\mem[28][13] ),
    .ZN(_04045_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09523_ (.A1(_03909_),
    .A2(_04030_),
    .B(_04045_),
    .ZN(_00432_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09524_ (.A1(_04028_),
    .A2(\mem[28][14] ),
    .ZN(_04046_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09525_ (.A1(_03911_),
    .A2(_04030_),
    .B(_04046_),
    .ZN(_00433_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09526_ (.A1(_04028_),
    .A2(\mem[28][15] ),
    .ZN(_04047_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09527_ (.A1(_03913_),
    .A2(_04030_),
    .B(_04047_),
    .ZN(_00434_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09528_ (.A1(_03522_),
    .A2(_03632_),
    .ZN(_04048_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09529_ (.I(_04048_),
    .Z(_04049_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09530_ (.I(_04048_),
    .Z(_04050_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09531_ (.A1(_04050_),
    .A2(\mem[2][0] ),
    .ZN(_04051_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09532_ (.A1(_03915_),
    .A2(_04049_),
    .B(_04051_),
    .ZN(_00435_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09533_ (.A1(_04050_),
    .A2(\mem[2][1] ),
    .ZN(_04052_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09534_ (.A1(_03920_),
    .A2(_04049_),
    .B(_04052_),
    .ZN(_00436_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09535_ (.A1(_04050_),
    .A2(\mem[2][2] ),
    .ZN(_04053_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09536_ (.A1(_03922_),
    .A2(_04049_),
    .B(_04053_),
    .ZN(_00437_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09537_ (.A1(_04050_),
    .A2(\mem[2][3] ),
    .ZN(_04054_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09538_ (.A1(_03924_),
    .A2(_04049_),
    .B(_04054_),
    .ZN(_00438_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09539_ (.I(_04048_),
    .Z(_04055_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09540_ (.A1(_04055_),
    .A2(\mem[2][4] ),
    .ZN(_04056_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09541_ (.A1(_03926_),
    .A2(_04049_),
    .B(_04056_),
    .ZN(_00439_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09542_ (.A1(_04055_),
    .A2(\mem[2][5] ),
    .ZN(_04057_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09543_ (.A1(_03929_),
    .A2(_04049_),
    .B(_04057_),
    .ZN(_00440_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09544_ (.A1(_04055_),
    .A2(\mem[2][6] ),
    .ZN(_04058_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09545_ (.A1(_03931_),
    .A2(_04049_),
    .B(_04058_),
    .ZN(_00441_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09546_ (.A1(_04055_),
    .A2(\mem[2][7] ),
    .ZN(_04059_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09547_ (.A1(_03933_),
    .A2(_04049_),
    .B(_04059_),
    .ZN(_00442_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09548_ (.A1(_04055_),
    .A2(\mem[2][8] ),
    .ZN(_04060_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09549_ (.A1(_03935_),
    .A2(_04049_),
    .B(_04060_),
    .ZN(_00443_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09550_ (.A1(_04055_),
    .A2(\mem[2][9] ),
    .ZN(_04061_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09551_ (.A1(_03937_),
    .A2(_04049_),
    .B(_04061_),
    .ZN(_00444_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09552_ (.A1(_04055_),
    .A2(\mem[2][10] ),
    .ZN(_04062_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09553_ (.A1(_03939_),
    .A2(_04050_),
    .B(_04062_),
    .ZN(_00445_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09554_ (.A1(_04055_),
    .A2(\mem[2][11] ),
    .ZN(_04063_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09555_ (.A1(_03941_),
    .A2(_04050_),
    .B(_04063_),
    .ZN(_00446_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09556_ (.A1(_04055_),
    .A2(\mem[2][12] ),
    .ZN(_04064_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09557_ (.A1(_03943_),
    .A2(_04050_),
    .B(_04064_),
    .ZN(_00447_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09558_ (.A1(_04055_),
    .A2(\mem[2][13] ),
    .ZN(_04065_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09559_ (.A1(_03909_),
    .A2(_04050_),
    .B(_04065_),
    .ZN(_00448_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09560_ (.A1(_04048_),
    .A2(\mem[2][14] ),
    .ZN(_04066_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09561_ (.A1(_03911_),
    .A2(_04050_),
    .B(_04066_),
    .ZN(_00449_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09562_ (.A1(_04048_),
    .A2(\mem[2][15] ),
    .ZN(_04067_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09563_ (.A1(_03913_),
    .A2(_04050_),
    .B(_04067_),
    .ZN(_00450_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09564_ (.A1(net119),
    .A2(_01162_),
    .ZN(_04068_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09565_ (.I(_04068_),
    .Z(_04069_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09566_ (.I(_04068_),
    .Z(_04070_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09567_ (.A1(_04070_),
    .A2(\mem[30][0] ),
    .ZN(_04071_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09568_ (.A1(_03915_),
    .A2(_04069_),
    .B(_04071_),
    .ZN(_00451_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09569_ (.A1(_04070_),
    .A2(\mem[30][1] ),
    .ZN(_04072_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09570_ (.A1(_03920_),
    .A2(_04069_),
    .B(_04072_),
    .ZN(_00452_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09571_ (.A1(_04070_),
    .A2(\mem[30][2] ),
    .ZN(_04073_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09572_ (.A1(_03922_),
    .A2(_04069_),
    .B(_04073_),
    .ZN(_00453_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09573_ (.A1(_04070_),
    .A2(\mem[30][3] ),
    .ZN(_04074_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09574_ (.A1(_03924_),
    .A2(_04069_),
    .B(_04074_),
    .ZN(_00454_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09575_ (.I(_04068_),
    .Z(_04075_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09576_ (.A1(_04075_),
    .A2(\mem[30][4] ),
    .ZN(_04076_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09577_ (.A1(_03926_),
    .A2(_04069_),
    .B(_04076_),
    .ZN(_00455_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09578_ (.A1(_04075_),
    .A2(\mem[30][5] ),
    .ZN(_04077_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09579_ (.A1(_03929_),
    .A2(_04069_),
    .B(_04077_),
    .ZN(_00456_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09580_ (.A1(_04075_),
    .A2(\mem[30][6] ),
    .ZN(_04078_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09581_ (.A1(_03931_),
    .A2(_04069_),
    .B(_04078_),
    .ZN(_00457_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09582_ (.A1(_04075_),
    .A2(\mem[30][7] ),
    .ZN(_04079_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09583_ (.A1(_03933_),
    .A2(_04069_),
    .B(_04079_),
    .ZN(_00458_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09584_ (.A1(_04075_),
    .A2(\mem[30][8] ),
    .ZN(_04080_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09585_ (.A1(_03935_),
    .A2(_04069_),
    .B(_04080_),
    .ZN(_00459_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09586_ (.A1(_04075_),
    .A2(\mem[30][9] ),
    .ZN(_04081_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09587_ (.A1(_03937_),
    .A2(_04069_),
    .B(_04081_),
    .ZN(_00460_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09588_ (.A1(_04075_),
    .A2(\mem[30][10] ),
    .ZN(_04082_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09589_ (.A1(_03939_),
    .A2(_04070_),
    .B(_04082_),
    .ZN(_00461_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09590_ (.A1(_04075_),
    .A2(\mem[30][11] ),
    .ZN(_04083_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09591_ (.A1(_03941_),
    .A2(_04070_),
    .B(_04083_),
    .ZN(_00462_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09592_ (.A1(_04075_),
    .A2(\mem[30][12] ),
    .ZN(_04084_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09593_ (.A1(_03943_),
    .A2(_04070_),
    .B(_04084_),
    .ZN(_00463_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09594_ (.A1(_04075_),
    .A2(\mem[30][13] ),
    .ZN(_04085_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09595_ (.A1(_03909_),
    .A2(_04070_),
    .B(_04085_),
    .ZN(_00464_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09596_ (.A1(_04068_),
    .A2(\mem[30][14] ),
    .ZN(_04086_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09597_ (.A1(_03911_),
    .A2(_04070_),
    .B(_04086_),
    .ZN(_00465_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09598_ (.A1(_04068_),
    .A2(\mem[30][15] ),
    .ZN(_04087_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09599_ (.A1(_03913_),
    .A2(_04070_),
    .B(_04087_),
    .ZN(_00466_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09600_ (.A1(net40),
    .A2(_01103_),
    .ZN(_04088_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09601_ (.I(_04088_),
    .Z(_04089_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09602_ (.I(_04088_),
    .Z(_04090_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09603_ (.A1(_04090_),
    .A2(\mem[31][0] ),
    .ZN(_04091_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09604_ (.A1(_03915_),
    .A2(_04089_),
    .B(_04091_),
    .ZN(_00467_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09605_ (.A1(_04090_),
    .A2(\mem[31][1] ),
    .ZN(_04092_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09606_ (.A1(_03920_),
    .A2(_04089_),
    .B(_04092_),
    .ZN(_00468_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09607_ (.A1(_04090_),
    .A2(\mem[31][2] ),
    .ZN(_04093_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09608_ (.A1(_03922_),
    .A2(_04089_),
    .B(_04093_),
    .ZN(_00469_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09609_ (.A1(_04090_),
    .A2(\mem[31][3] ),
    .ZN(_04094_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09610_ (.A1(_03924_),
    .A2(_04089_),
    .B(_04094_),
    .ZN(_00470_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09611_ (.I(_04088_),
    .Z(_04095_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09612_ (.A1(_04095_),
    .A2(\mem[31][4] ),
    .ZN(_04096_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09613_ (.A1(_03926_),
    .A2(_04089_),
    .B(_04096_),
    .ZN(_00471_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09614_ (.A1(_04095_),
    .A2(\mem[31][5] ),
    .ZN(_04097_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09615_ (.A1(_03929_),
    .A2(_04089_),
    .B(_04097_),
    .ZN(_00472_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09616_ (.A1(_04095_),
    .A2(\mem[31][6] ),
    .ZN(_04098_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09617_ (.A1(_03931_),
    .A2(_04089_),
    .B(_04098_),
    .ZN(_00473_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09618_ (.A1(_04095_),
    .A2(\mem[31][7] ),
    .ZN(_04099_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09619_ (.A1(_03933_),
    .A2(_04089_),
    .B(_04099_),
    .ZN(_00474_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09620_ (.A1(_04095_),
    .A2(\mem[31][8] ),
    .ZN(_04100_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09621_ (.A1(_03935_),
    .A2(_04089_),
    .B(_04100_),
    .ZN(_00475_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09622_ (.A1(_04095_),
    .A2(\mem[31][9] ),
    .ZN(_04101_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09623_ (.A1(_03937_),
    .A2(_04089_),
    .B(_04101_),
    .ZN(_00476_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09624_ (.A1(_04095_),
    .A2(\mem[31][10] ),
    .ZN(_04102_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09625_ (.A1(_03939_),
    .A2(_04090_),
    .B(_04102_),
    .ZN(_00477_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09626_ (.A1(_04095_),
    .A2(\mem[31][11] ),
    .ZN(_04103_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09627_ (.A1(_03941_),
    .A2(_04090_),
    .B(_04103_),
    .ZN(_00478_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09628_ (.A1(_04095_),
    .A2(\mem[31][12] ),
    .ZN(_04104_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09629_ (.A1(_03943_),
    .A2(_04090_),
    .B(_04104_),
    .ZN(_00479_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09630_ (.A1(_04095_),
    .A2(\mem[31][13] ),
    .ZN(_04105_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09631_ (.A1(_03909_),
    .A2(_04090_),
    .B(_04105_),
    .ZN(_00480_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09632_ (.A1(_04088_),
    .A2(\mem[31][14] ),
    .ZN(_04106_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09633_ (.A1(_03911_),
    .A2(_04090_),
    .B(_04106_),
    .ZN(_00481_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09634_ (.A1(_04088_),
    .A2(\mem[31][15] ),
    .ZN(_04107_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09635_ (.A1(_03913_),
    .A2(_04090_),
    .B(_04107_),
    .ZN(_00482_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09636_ (.A1(_03588_),
    .A2(_01127_),
    .ZN(_04108_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09637_ (.I(_04108_),
    .Z(_04109_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09638_ (.I(_04108_),
    .Z(_04110_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09639_ (.A1(_04110_),
    .A2(\mem[32][0] ),
    .ZN(_04111_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09640_ (.A1(_03915_),
    .A2(_04109_),
    .B(_04111_),
    .ZN(_00483_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09641_ (.A1(_04110_),
    .A2(\mem[32][1] ),
    .ZN(_04112_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09642_ (.A1(_03920_),
    .A2(_04109_),
    .B(_04112_),
    .ZN(_00484_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09643_ (.A1(_04110_),
    .A2(\mem[32][2] ),
    .ZN(_04113_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09644_ (.A1(_03922_),
    .A2(_04109_),
    .B(_04113_),
    .ZN(_00485_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09645_ (.A1(_04110_),
    .A2(\mem[32][3] ),
    .ZN(_04114_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09646_ (.A1(_03924_),
    .A2(_04109_),
    .B(_04114_),
    .ZN(_00486_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09647_ (.I(_04108_),
    .Z(_04115_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09648_ (.A1(_04115_),
    .A2(\mem[32][4] ),
    .ZN(_04116_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09649_ (.A1(_03926_),
    .A2(_04109_),
    .B(_04116_),
    .ZN(_00487_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09650_ (.A1(_04115_),
    .A2(\mem[32][5] ),
    .ZN(_04117_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09651_ (.A1(_03929_),
    .A2(_04109_),
    .B(_04117_),
    .ZN(_00488_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09652_ (.A1(_04115_),
    .A2(\mem[32][6] ),
    .ZN(_04118_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09653_ (.A1(_03931_),
    .A2(_04109_),
    .B(_04118_),
    .ZN(_00489_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09654_ (.A1(_04115_),
    .A2(\mem[32][7] ),
    .ZN(_04119_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09655_ (.A1(_03933_),
    .A2(_04109_),
    .B(_04119_),
    .ZN(_00490_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09656_ (.A1(_04115_),
    .A2(\mem[32][8] ),
    .ZN(_04120_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09657_ (.A1(_03935_),
    .A2(_04109_),
    .B(_04120_),
    .ZN(_00491_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09658_ (.A1(_04115_),
    .A2(\mem[32][9] ),
    .ZN(_04121_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09659_ (.A1(_03937_),
    .A2(_04109_),
    .B(_04121_),
    .ZN(_00492_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09660_ (.A1(_04115_),
    .A2(\mem[32][10] ),
    .ZN(_04122_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09661_ (.A1(_03939_),
    .A2(_04110_),
    .B(_04122_),
    .ZN(_00493_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09662_ (.A1(_04115_),
    .A2(\mem[32][11] ),
    .ZN(_04123_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09663_ (.A1(_03941_),
    .A2(_04110_),
    .B(_04123_),
    .ZN(_00494_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09664_ (.A1(_04115_),
    .A2(\mem[32][12] ),
    .ZN(_04124_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09665_ (.A1(_03943_),
    .A2(_04110_),
    .B(_04124_),
    .ZN(_00495_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09666_ (.I(_03438_),
    .Z(_04125_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09667_ (.A1(_04115_),
    .A2(\mem[32][13] ),
    .ZN(_04126_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09668_ (.A1(_04125_),
    .A2(_04110_),
    .B(_04126_),
    .ZN(_00496_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09669_ (.I(_03446_),
    .Z(_04127_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09670_ (.A1(_04108_),
    .A2(\mem[32][14] ),
    .ZN(_04128_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09671_ (.A1(_04127_),
    .A2(_04110_),
    .B(_04128_),
    .ZN(_00497_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09672_ (.I(_03449_),
    .Z(_04129_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09673_ (.A1(_04108_),
    .A2(\mem[32][15] ),
    .ZN(_04130_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09674_ (.A1(_04129_),
    .A2(_04110_),
    .B(_04130_),
    .ZN(_00498_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09675_ (.I(_03452_),
    .Z(_04131_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09676_ (.A1(net93),
    .A2(_01127_),
    .ZN(_04132_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09677_ (.I(_04132_),
    .Z(_04133_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09678_ (.I(_04132_),
    .Z(_04134_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09679_ (.A1(_04134_),
    .A2(\mem[33][0] ),
    .ZN(_04135_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09680_ (.A1(_04131_),
    .A2(_04133_),
    .B(_04135_),
    .ZN(_00499_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09681_ (.I(_03461_),
    .Z(_04136_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09682_ (.A1(_04134_),
    .A2(\mem[33][1] ),
    .ZN(_04137_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09683_ (.A1(_04136_),
    .A2(_04133_),
    .B(_04137_),
    .ZN(_00500_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09684_ (.I(_03464_),
    .Z(_04138_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09685_ (.A1(_04134_),
    .A2(\mem[33][2] ),
    .ZN(_04139_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09686_ (.A1(_04138_),
    .A2(_04133_),
    .B(_04139_),
    .ZN(_00501_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09687_ (.I(_03467_),
    .Z(_04140_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09688_ (.A1(_04134_),
    .A2(\mem[33][3] ),
    .ZN(_04141_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09689_ (.A1(_04140_),
    .A2(_04133_),
    .B(_04141_),
    .ZN(_00502_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09690_ (.I(_03470_),
    .Z(_04142_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09691_ (.I(_04132_),
    .Z(_04143_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09692_ (.A1(_04143_),
    .A2(\mem[33][4] ),
    .ZN(_04144_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09693_ (.A1(_04142_),
    .A2(_04133_),
    .B(_04144_),
    .ZN(_00503_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09694_ (.I(_03474_),
    .Z(_04145_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09695_ (.A1(_04143_),
    .A2(\mem[33][5] ),
    .ZN(_04146_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09696_ (.A1(_04145_),
    .A2(_04133_),
    .B(_04146_),
    .ZN(_00504_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09697_ (.I(_03477_),
    .Z(_04147_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09698_ (.A1(_04143_),
    .A2(\mem[33][6] ),
    .ZN(_04148_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09699_ (.A1(_04147_),
    .A2(_04133_),
    .B(_04148_),
    .ZN(_00505_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09700_ (.I(_03480_),
    .Z(_04149_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09701_ (.A1(_04143_),
    .A2(\mem[33][7] ),
    .ZN(_04150_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09702_ (.A1(_04149_),
    .A2(_04133_),
    .B(_04150_),
    .ZN(_00506_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09703_ (.I(_03483_),
    .Z(_04151_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09704_ (.A1(_04143_),
    .A2(\mem[33][8] ),
    .ZN(_04152_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09705_ (.A1(_04151_),
    .A2(_04133_),
    .B(_04152_),
    .ZN(_00507_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09706_ (.I(_03486_),
    .Z(_04153_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09707_ (.A1(_04143_),
    .A2(\mem[33][9] ),
    .ZN(_04154_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09708_ (.D(_00016_),
    .CLK(clknet_leaf_71_i_clk),
    .Q(\mem[7][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09709_ (.D(_00017_),
    .CLK(clknet_leaf_41_i_clk),
    .Q(\mem[7][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09710_ (.D(_00018_),
    .CLK(clknet_leaf_41_i_clk),
    .Q(\mem[7][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09711_ (.D(_00019_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[59][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09712_ (.D(_00020_),
    .CLK(clknet_leaf_22_i_clk),
    .Q(\mem[59][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09713_ (.D(_00021_),
    .CLK(clknet_leaf_22_i_clk),
    .Q(\mem[59][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09714_ (.D(_00022_),
    .CLK(clknet_leaf_22_i_clk),
    .Q(\mem[59][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09715_ (.D(_00023_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[59][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09716_ (.D(_00024_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[59][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09717_ (.D(_00025_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[59][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09718_ (.D(_00026_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[59][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09719_ (.D(_00027_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[59][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09720_ (.D(_00028_),
    .CLK(clknet_leaf_22_i_clk),
    .Q(\mem[59][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09721_ (.D(_00029_),
    .CLK(clknet_leaf_16_i_clk),
    .Q(\mem[59][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09722_ (.D(_00030_),
    .CLK(clknet_leaf_16_i_clk),
    .Q(\mem[59][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09723_ (.D(_00031_),
    .CLK(clknet_leaf_30_i_clk),
    .Q(\mem[59][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09724_ (.D(_00032_),
    .CLK(clknet_leaf_16_i_clk),
    .Q(\mem[59][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09725_ (.D(_00033_),
    .CLK(clknet_leaf_38_i_clk),
    .Q(\mem[59][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09726_ (.D(_00034_),
    .CLK(clknet_leaf_38_i_clk),
    .Q(\mem[59][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09727_ (.D(_00035_),
    .CLK(clknet_leaf_38_i_clk),
    .Q(\mem[63][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09728_ (.D(_00036_),
    .CLK(clknet_leaf_16_i_clk),
    .Q(\mem[63][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09729_ (.D(_00037_),
    .CLK(clknet_leaf_22_i_clk),
    .Q(\mem[63][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09730_ (.D(_00038_),
    .CLK(clknet_leaf_22_i_clk),
    .Q(\mem[63][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09731_ (.D(_00039_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[63][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09732_ (.D(_00040_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[63][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09733_ (.D(_00041_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[63][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09734_ (.D(_00042_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[63][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09735_ (.D(_00043_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[63][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09736_ (.D(_00044_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[63][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09737_ (.D(_00045_),
    .CLK(clknet_leaf_16_i_clk),
    .Q(\mem[63][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09738_ (.D(_00046_),
    .CLK(clknet_leaf_23_i_clk),
    .Q(\mem[63][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09739_ (.D(_00047_),
    .CLK(clknet_leaf_38_i_clk),
    .Q(\mem[63][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09740_ (.D(_00048_),
    .CLK(clknet_leaf_16_i_clk),
    .Q(\mem[63][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09741_ (.D(_00049_),
    .CLK(clknet_leaf_38_i_clk),
    .Q(\mem[63][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09742_ (.D(_00050_),
    .CLK(clknet_leaf_38_i_clk),
    .Q(\mem[63][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09743_ (.D(_00051_),
    .CLK(clknet_leaf_42_i_clk),
    .Q(\mem[6][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09744_ (.D(_00052_),
    .CLK(clknet_leaf_41_i_clk),
    .Q(\mem[6][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09745_ (.D(_00053_),
    .CLK(clknet_leaf_40_i_clk),
    .Q(\mem[6][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09746_ (.D(_00054_),
    .CLK(clknet_leaf_40_i_clk),
    .Q(\mem[6][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09747_ (.D(_00055_),
    .CLK(clknet_leaf_40_i_clk),
    .Q(\mem[6][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09748_ (.D(_00056_),
    .CLK(clknet_leaf_40_i_clk),
    .Q(\mem[6][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09749_ (.D(_00057_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[6][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09750_ (.D(_00058_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[6][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09751_ (.D(_00059_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[6][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09752_ (.D(_00060_),
    .CLK(clknet_leaf_40_i_clk),
    .Q(\mem[6][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09753_ (.D(_00061_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[6][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09754_ (.D(_00062_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[6][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09755_ (.D(_00063_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[6][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09756_ (.D(_00064_),
    .CLK(clknet_leaf_42_i_clk),
    .Q(\mem[6][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09757_ (.D(_00065_),
    .CLK(clknet_leaf_41_i_clk),
    .Q(\mem[6][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09758_ (.D(_00066_),
    .CLK(clknet_leaf_42_i_clk),
    .Q(\mem[6][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09759_ (.D(_00067_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[19][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09760_ (.D(_00068_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[19][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09761_ (.D(_00069_),
    .CLK(clknet_leaf_4_i_clk),
    .Q(\mem[19][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09762_ (.D(_00070_),
    .CLK(clknet_leaf_3_i_clk),
    .Q(\mem[19][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09763_ (.D(_00071_),
    .CLK(clknet_leaf_3_i_clk),
    .Q(\mem[19][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09764_ (.D(_00072_),
    .CLK(clknet_leaf_3_i_clk),
    .Q(\mem[19][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09765_ (.D(_00073_),
    .CLK(clknet_leaf_3_i_clk),
    .Q(\mem[19][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09766_ (.D(_00074_),
    .CLK(clknet_leaf_3_i_clk),
    .Q(\mem[19][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09767_ (.D(_00075_),
    .CLK(clknet_leaf_3_i_clk),
    .Q(\mem[19][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09768_ (.D(_00076_),
    .CLK(clknet_leaf_2_i_clk),
    .Q(\mem[19][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09769_ (.D(_00077_),
    .CLK(clknet_leaf_2_i_clk),
    .Q(\mem[19][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09770_ (.D(_00078_),
    .CLK(clknet_leaf_2_i_clk),
    .Q(\mem[19][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09771_ (.D(_00079_),
    .CLK(clknet_leaf_2_i_clk),
    .Q(\mem[19][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09772_ (.D(_00080_),
    .CLK(clknet_leaf_2_i_clk),
    .Q(\mem[19][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09773_ (.D(_00081_),
    .CLK(clknet_leaf_1_i_clk),
    .Q(\mem[19][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09774_ (.D(_00082_),
    .CLK(clknet_leaf_1_i_clk),
    .Q(\mem[19][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09775_ (.D(_00083_),
    .CLK(clknet_leaf_101_i_clk),
    .Q(\mem[29][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09776_ (.D(_00084_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[29][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09777_ (.D(_00085_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[29][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09778_ (.D(_00086_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[29][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09779_ (.D(_00087_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[29][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09780_ (.D(_00088_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[29][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09781_ (.D(_00089_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[29][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09782_ (.D(_00090_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[29][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09783_ (.D(_00091_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[29][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09784_ (.D(_00092_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[29][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09785_ (.D(_00093_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[29][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09786_ (.D(_00094_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[29][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09787_ (.D(_00095_),
    .CLK(clknet_leaf_101_i_clk),
    .Q(\mem[29][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09788_ (.D(_00096_),
    .CLK(clknet_leaf_101_i_clk),
    .Q(\mem[29][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09789_ (.D(_00097_),
    .CLK(clknet_leaf_101_i_clk),
    .Q(\mem[29][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09790_ (.D(_00098_),
    .CLK(clknet_leaf_101_i_clk),
    .Q(\mem[29][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09791_ (.D(_00099_),
    .CLK(clknet_leaf_11_i_clk),
    .Q(\mem[8][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09792_ (.D(_00100_),
    .CLK(clknet_leaf_11_i_clk),
    .Q(\mem[8][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09793_ (.D(_00101_),
    .CLK(clknet_leaf_10_i_clk),
    .Q(\mem[8][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09794_ (.D(_00102_),
    .CLK(clknet_leaf_10_i_clk),
    .Q(\mem[8][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09795_ (.D(_00103_),
    .CLK(clknet_leaf_10_i_clk),
    .Q(\mem[8][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09796_ (.D(_00104_),
    .CLK(clknet_leaf_10_i_clk),
    .Q(\mem[8][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09797_ (.D(_00105_),
    .CLK(clknet_leaf_11_i_clk),
    .Q(\mem[8][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09798_ (.D(_00106_),
    .CLK(clknet_leaf_7_i_clk),
    .Q(\mem[8][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09799_ (.D(_00107_),
    .CLK(clknet_leaf_7_i_clk),
    .Q(\mem[8][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09800_ (.D(_00108_),
    .CLK(clknet_leaf_7_i_clk),
    .Q(\mem[8][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09801_ (.D(_00109_),
    .CLK(clknet_leaf_7_i_clk),
    .Q(\mem[8][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09802_ (.D(_00110_),
    .CLK(clknet_leaf_6_i_clk),
    .Q(\mem[8][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09803_ (.D(_00111_),
    .CLK(clknet_leaf_6_i_clk),
    .Q(\mem[8][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09804_ (.D(_00112_),
    .CLK(clknet_leaf_17_i_clk),
    .Q(\mem[8][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09805_ (.D(_00113_),
    .CLK(clknet_leaf_17_i_clk),
    .Q(\mem[8][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09806_ (.D(_00114_),
    .CLK(clknet_leaf_17_i_clk),
    .Q(\mem[8][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09807_ (.D(_00115_),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[0][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09808_ (.D(_00116_),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[0][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09809_ (.D(_00117_),
    .CLK(clknet_leaf_103_i_clk),
    .Q(\mem[0][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09810_ (.D(_00118_),
    .CLK(clknet_leaf_12_i_clk),
    .Q(\mem[0][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09811_ (.D(_00119_),
    .CLK(clknet_leaf_13_i_clk),
    .Q(\mem[0][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09812_ (.D(_00120_),
    .CLK(clknet_leaf_12_i_clk),
    .Q(\mem[0][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09813_ (.D(_00121_),
    .CLK(clknet_leaf_12_i_clk),
    .Q(\mem[0][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09814_ (.D(_00122_),
    .CLK(clknet_leaf_13_i_clk),
    .Q(\mem[0][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09815_ (.D(_00123_),
    .CLK(clknet_leaf_13_i_clk),
    .Q(\mem[0][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09816_ (.D(_00124_),
    .CLK(clknet_leaf_13_i_clk),
    .Q(\mem[0][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09817_ (.D(_00125_),
    .CLK(clknet_leaf_13_i_clk),
    .Q(\mem[0][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09818_ (.D(_00126_),
    .CLK(clknet_leaf_40_i_clk),
    .Q(\mem[0][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09819_ (.D(_00127_),
    .CLK(clknet_leaf_41_i_clk),
    .Q(\mem[0][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09820_ (.D(_00128_),
    .CLK(clknet_leaf_41_i_clk),
    .Q(\mem[0][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09821_ (.D(_00129_),
    .CLK(clknet_leaf_41_i_clk),
    .Q(\mem[0][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09822_ (.D(_00130_),
    .CLK(clknet_leaf_41_i_clk),
    .Q(\mem[0][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09823_ (.D(_00131_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[10][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09824_ (.D(_00132_),
    .CLK(clknet_leaf_38_i_clk),
    .Q(\mem[10][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09825_ (.D(_00133_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[10][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09826_ (.D(_00134_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[10][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09827_ (.D(_00135_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[10][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09828_ (.D(_00136_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[10][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09829_ (.D(_00137_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[10][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09830_ (.D(_00138_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[10][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09831_ (.D(_00139_),
    .CLK(clknet_leaf_16_i_clk),
    .Q(\mem[10][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09832_ (.D(_00140_),
    .CLK(clknet_leaf_16_i_clk),
    .Q(\mem[10][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09833_ (.D(_00141_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[10][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09834_ (.D(_00142_),
    .CLK(clknet_leaf_16_i_clk),
    .Q(\mem[10][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09835_ (.D(_00143_),
    .CLK(clknet_leaf_14_i_clk),
    .Q(\mem[10][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09836_ (.D(_00144_),
    .CLK(clknet_leaf_17_i_clk),
    .Q(\mem[10][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09837_ (.D(_00145_),
    .CLK(clknet_leaf_17_i_clk),
    .Q(\mem[10][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09838_ (.D(_00146_),
    .CLK(clknet_leaf_17_i_clk),
    .Q(\mem[10][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09839_ (.D(_00147_),
    .CLK(clknet_leaf_16_i_clk),
    .Q(\mem[11][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09840_ (.D(_00148_),
    .CLK(clknet_leaf_22_i_clk),
    .Q(\mem[11][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09841_ (.D(_00149_),
    .CLK(clknet_leaf_21_i_clk),
    .Q(\mem[11][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09842_ (.D(_00150_),
    .CLK(clknet_leaf_22_i_clk),
    .Q(\mem[11][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09843_ (.D(_00151_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[11][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09844_ (.D(_00152_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[11][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09845_ (.D(_00153_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[11][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09846_ (.D(_00154_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[11][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09847_ (.D(_00155_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[11][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09848_ (.D(_00156_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[11][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09849_ (.D(_00157_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[11][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09850_ (.D(_00158_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[11][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09851_ (.D(_00159_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[11][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09852_ (.D(_00160_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[11][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09853_ (.D(_00161_),
    .CLK(clknet_leaf_17_i_clk),
    .Q(\mem[11][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09854_ (.D(_00162_),
    .CLK(clknet_leaf_17_i_clk),
    .Q(\mem[11][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09855_ (.D(_00163_),
    .CLK(clknet_leaf_17_i_clk),
    .Q(\mem[12][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09856_ (.D(_00164_),
    .CLK(clknet_leaf_17_i_clk),
    .Q(\mem[12][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09857_ (.D(_00165_),
    .CLK(clknet_leaf_18_i_clk),
    .Q(\mem[12][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09858_ (.D(_00166_),
    .CLK(clknet_leaf_18_i_clk),
    .Q(\mem[12][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09859_ (.D(_00167_),
    .CLK(clknet_leaf_19_i_clk),
    .Q(\mem[12][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09860_ (.D(_00168_),
    .CLK(clknet_leaf_19_i_clk),
    .Q(\mem[12][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09861_ (.D(_00169_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[12][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09862_ (.D(_00170_),
    .CLK(clknet_leaf_19_i_clk),
    .Q(\mem[12][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09863_ (.D(_00171_),
    .CLK(clknet_leaf_19_i_clk),
    .Q(\mem[12][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09864_ (.D(_00172_),
    .CLK(clknet_leaf_19_i_clk),
    .Q(\mem[12][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09865_ (.D(_00173_),
    .CLK(clknet_leaf_20_i_clk),
    .Q(\mem[12][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09866_ (.D(_00174_),
    .CLK(clknet_leaf_18_i_clk),
    .Q(\mem[12][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09867_ (.D(_00175_),
    .CLK(clknet_leaf_18_i_clk),
    .Q(\mem[12][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09868_ (.D(_00176_),
    .CLK(clknet_leaf_18_i_clk),
    .Q(\mem[12][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09869_ (.D(_00177_),
    .CLK(clknet_leaf_18_i_clk),
    .Q(\mem[12][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09870_ (.D(_00178_),
    .CLK(clknet_leaf_18_i_clk),
    .Q(\mem[12][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09871_ (.D(_00179_),
    .CLK(clknet_leaf_6_i_clk),
    .Q(\mem[13][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09872_ (.D(_00180_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[13][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09873_ (.D(_00181_),
    .CLK(clknet_leaf_6_i_clk),
    .Q(\mem[13][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09874_ (.D(_00182_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[13][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09875_ (.D(_00183_),
    .CLK(clknet_leaf_4_i_clk),
    .Q(\mem[13][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09876_ (.D(_00184_),
    .CLK(clknet_leaf_4_i_clk),
    .Q(\mem[13][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09877_ (.D(_00185_),
    .CLK(clknet_leaf_4_i_clk),
    .Q(\mem[13][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09878_ (.D(_00186_),
    .CLK(clknet_leaf_5_i_clk),
    .Q(\mem[13][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09879_ (.D(_00187_),
    .CLK(clknet_leaf_4_i_clk),
    .Q(\mem[13][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09880_ (.D(_00188_),
    .CLK(clknet_leaf_5_i_clk),
    .Q(\mem[13][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09881_ (.D(_00189_),
    .CLK(clknet_leaf_5_i_clk),
    .Q(\mem[13][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09882_ (.D(_00190_),
    .CLK(clknet_leaf_5_i_clk),
    .Q(\mem[13][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09883_ (.D(_00191_),
    .CLK(clknet_leaf_5_i_clk),
    .Q(\mem[13][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09884_ (.D(_00192_),
    .CLK(clknet_leaf_5_i_clk),
    .Q(\mem[13][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09885_ (.D(_00193_),
    .CLK(clknet_leaf_6_i_clk),
    .Q(\mem[13][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09886_ (.D(_00194_),
    .CLK(clknet_leaf_6_i_clk),
    .Q(\mem[13][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09887_ (.D(_00195_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[14][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09888_ (.D(_00196_),
    .CLK(clknet_leaf_7_i_clk),
    .Q(\mem[14][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09889_ (.D(_00197_),
    .CLK(clknet_leaf_6_i_clk),
    .Q(\mem[14][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09890_ (.D(_00198_),
    .CLK(clknet_leaf_6_i_clk),
    .Q(\mem[14][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09891_ (.D(_00199_),
    .CLK(clknet_leaf_5_i_clk),
    .Q(\mem[14][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09892_ (.D(_00200_),
    .CLK(clknet_leaf_4_i_clk),
    .Q(\mem[14][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09893_ (.D(_00201_),
    .CLK(clknet_leaf_4_i_clk),
    .Q(\mem[14][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09894_ (.D(_00202_),
    .CLK(clknet_leaf_5_i_clk),
    .Q(\mem[14][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09895_ (.D(_00203_),
    .CLK(clknet_leaf_5_i_clk),
    .Q(\mem[14][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09896_ (.D(_00204_),
    .CLK(clknet_leaf_19_i_clk),
    .Q(\mem[14][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09897_ (.D(_00205_),
    .CLK(clknet_leaf_19_i_clk),
    .Q(\mem[14][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09898_ (.D(_00206_),
    .CLK(clknet_leaf_5_i_clk),
    .Q(\mem[14][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09899_ (.D(_00207_),
    .CLK(clknet_leaf_6_i_clk),
    .Q(\mem[14][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09900_ (.D(_00208_),
    .CLK(clknet_leaf_18_i_clk),
    .Q(\mem[14][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09901_ (.D(_00209_),
    .CLK(clknet_leaf_6_i_clk),
    .Q(\mem[14][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09902_ (.D(_00210_),
    .CLK(clknet_leaf_18_i_clk),
    .Q(\mem[14][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09903_ (.D(_00211_),
    .CLK(clknet_leaf_10_i_clk),
    .Q(\mem[15][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09904_ (.D(_00212_),
    .CLK(clknet_leaf_9_i_clk),
    .Q(\mem[15][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09905_ (.D(_00213_),
    .CLK(clknet_leaf_9_i_clk),
    .Q(\mem[15][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09906_ (.D(_00214_),
    .CLK(clknet_leaf_10_i_clk),
    .Q(\mem[15][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09907_ (.D(_00215_),
    .CLK(clknet_leaf_9_i_clk),
    .Q(\mem[15][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09908_ (.D(_00216_),
    .CLK(clknet_leaf_9_i_clk),
    .Q(\mem[15][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09909_ (.D(_00217_),
    .CLK(clknet_leaf_9_i_clk),
    .Q(\mem[15][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09910_ (.D(_00218_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[15][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09911_ (.D(_00219_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[15][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09912_ (.D(_00220_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[15][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09913_ (.D(_00221_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[15][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09914_ (.D(_00222_),
    .CLK(clknet_leaf_7_i_clk),
    .Q(\mem[15][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09915_ (.D(_00223_),
    .CLK(clknet_leaf_7_i_clk),
    .Q(\mem[15][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09916_ (.D(_00224_),
    .CLK(clknet_leaf_7_i_clk),
    .Q(\mem[15][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09917_ (.D(_00225_),
    .CLK(clknet_leaf_11_i_clk),
    .Q(\mem[15][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09918_ (.D(_00226_),
    .CLK(clknet_leaf_7_i_clk),
    .Q(\mem[15][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09919_ (.D(_00227_),
    .CLK(clknet_leaf_105_i_clk),
    .Q(\mem[16][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09920_ (.D(_00228_),
    .CLK(clknet_leaf_106_i_clk),
    .Q(\mem[16][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09921_ (.D(_00229_),
    .CLK(clknet_leaf_106_i_clk),
    .Q(\mem[16][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09922_ (.D(_00230_),
    .CLK(clknet_leaf_106_i_clk),
    .Q(\mem[16][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09923_ (.D(_00231_),
    .CLK(clknet_leaf_112_i_clk),
    .Q(\mem[16][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09924_ (.D(_00232_),
    .CLK(clknet_leaf_111_i_clk),
    .Q(\mem[16][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09925_ (.D(_00233_),
    .CLK(clknet_leaf_111_i_clk),
    .Q(\mem[16][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09926_ (.D(_00234_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[16][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09927_ (.D(_00235_),
    .CLK(clknet_leaf_111_i_clk),
    .Q(\mem[16][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09928_ (.D(_00236_),
    .CLK(clknet_leaf_111_i_clk),
    .Q(\mem[16][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09929_ (.D(_00237_),
    .CLK(clknet_leaf_111_i_clk),
    .Q(\mem[16][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09930_ (.D(_00238_),
    .CLK(clknet_leaf_111_i_clk),
    .Q(\mem[16][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09931_ (.D(_00239_),
    .CLK(clknet_leaf_111_i_clk),
    .Q(\mem[16][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09932_ (.D(_00240_),
    .CLK(clknet_leaf_112_i_clk),
    .Q(\mem[16][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09933_ (.D(_00241_),
    .CLK(clknet_leaf_112_i_clk),
    .Q(\mem[16][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09934_ (.D(_00242_),
    .CLK(clknet_leaf_106_i_clk),
    .Q(\mem[16][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09935_ (.D(_00243_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[17][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09936_ (.D(_00244_),
    .CLK(clknet_leaf_8_i_clk),
    .Q(\mem[17][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09937_ (.D(_00245_),
    .CLK(clknet_leaf_9_i_clk),
    .Q(\mem[17][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09938_ (.D(_00246_),
    .CLK(clknet_leaf_1_i_clk),
    .Q(\mem[17][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09939_ (.D(_00247_),
    .CLK(clknet_leaf_113_i_clk),
    .Q(\mem[17][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09940_ (.D(_00248_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[17][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09941_ (.D(_00249_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[17][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09942_ (.D(_00250_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[17][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09943_ (.D(_00251_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[17][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09944_ (.D(_00252_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[17][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09945_ (.D(_00253_),
    .CLK(clknet_leaf_114_i_clk),
    .Q(\mem[17][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09946_ (.D(_00254_),
    .CLK(clknet_leaf_114_i_clk),
    .Q(\mem[17][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09947_ (.D(_00255_),
    .CLK(clknet_leaf_113_i_clk),
    .Q(\mem[17][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09948_ (.D(_00256_),
    .CLK(clknet_leaf_113_i_clk),
    .Q(\mem[17][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09949_ (.D(_00257_),
    .CLK(clknet_leaf_113_i_clk),
    .Q(\mem[17][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09950_ (.D(_00258_),
    .CLK(clknet_leaf_1_i_clk),
    .Q(\mem[17][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09951_ (.D(_00259_),
    .CLK(clknet_leaf_9_i_clk),
    .Q(\mem[18][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09952_ (.D(_00260_),
    .CLK(clknet_leaf_9_i_clk),
    .Q(\mem[18][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09953_ (.D(_00261_),
    .CLK(clknet_leaf_9_i_clk),
    .Q(\mem[18][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09954_ (.D(_00262_),
    .CLK(clknet_leaf_1_i_clk),
    .Q(\mem[18][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09955_ (.D(_00263_),
    .CLK(clknet_leaf_113_i_clk),
    .Q(\mem[18][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09956_ (.D(_00264_),
    .CLK(clknet_leaf_114_i_clk),
    .Q(\mem[18][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09957_ (.D(_00265_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[18][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09958_ (.D(_00266_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[18][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09959_ (.D(_00267_),
    .CLK(clknet_leaf_114_i_clk),
    .Q(\mem[18][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09960_ (.D(_00268_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[18][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09961_ (.D(_00269_),
    .CLK(clknet_leaf_114_i_clk),
    .Q(\mem[18][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09962_ (.D(_00270_),
    .CLK(clknet_leaf_114_i_clk),
    .Q(\mem[18][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09963_ (.D(_00271_),
    .CLK(clknet_leaf_113_i_clk),
    .Q(\mem[18][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09964_ (.D(_00272_),
    .CLK(clknet_leaf_113_i_clk),
    .Q(\mem[18][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09965_ (.D(_00273_),
    .CLK(clknet_leaf_113_i_clk),
    .Q(\mem[18][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09966_ (.D(_00274_),
    .CLK(clknet_leaf_113_i_clk),
    .Q(\mem[18][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09967_ (.D(_00275_),
    .CLK(clknet_leaf_11_i_clk),
    .Q(\mem[1][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09968_ (.D(_00276_),
    .CLK(clknet_leaf_12_i_clk),
    .Q(\mem[1][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09969_ (.D(_00277_),
    .CLK(clknet_leaf_11_i_clk),
    .Q(\mem[1][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09970_ (.D(_00278_),
    .CLK(clknet_leaf_10_i_clk),
    .Q(\mem[1][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09971_ (.D(_00279_),
    .CLK(clknet_leaf_10_i_clk),
    .Q(\mem[1][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09972_ (.D(_00280_),
    .CLK(clknet_leaf_10_i_clk),
    .Q(\mem[1][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09973_ (.D(_00281_),
    .CLK(clknet_leaf_105_i_clk),
    .Q(\mem[1][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09974_ (.D(_00282_),
    .CLK(clknet_leaf_105_i_clk),
    .Q(\mem[1][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09975_ (.D(_00283_),
    .CLK(clknet_leaf_105_i_clk),
    .Q(\mem[1][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09976_ (.D(_00284_),
    .CLK(clknet_leaf_12_i_clk),
    .Q(\mem[1][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09977_ (.D(_00285_),
    .CLK(clknet_leaf_12_i_clk),
    .Q(\mem[1][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09978_ (.D(_00286_),
    .CLK(clknet_leaf_11_i_clk),
    .Q(\mem[1][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09979_ (.D(_00287_),
    .CLK(clknet_leaf_12_i_clk),
    .Q(\mem[1][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09980_ (.D(_00288_),
    .CLK(clknet_leaf_11_i_clk),
    .Q(\mem[1][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09981_ (.D(_00289_),
    .CLK(clknet_leaf_12_i_clk),
    .Q(\mem[1][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09982_ (.D(_00290_),
    .CLK(clknet_leaf_13_i_clk),
    .Q(\mem[1][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09983_ (.D(_00291_),
    .CLK(clknet_leaf_1_i_clk),
    .Q(\mem[20][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09984_ (.D(_00292_),
    .CLK(clknet_leaf_1_i_clk),
    .Q(\mem[20][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09985_ (.D(_00293_),
    .CLK(clknet_leaf_2_i_clk),
    .Q(\mem[20][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09986_ (.D(_00294_),
    .CLK(clknet_leaf_2_i_clk),
    .Q(\mem[20][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09987_ (.D(_00295_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[20][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09988_ (.D(_00296_),
    .CLK(clknet_leaf_2_i_clk),
    .Q(\mem[20][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09989_ (.D(_00297_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[20][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09990_ (.D(_00298_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[20][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09991_ (.D(_00299_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[20][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09992_ (.D(_00300_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[20][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09993_ (.D(_00301_),
    .CLK(clknet_leaf_0_i_clk),
    .Q(\mem[20][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09994_ (.D(_00302_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[20][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09995_ (.D(_00303_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[20][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09996_ (.D(_00304_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[20][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09997_ (.D(_00305_),
    .CLK(clknet_leaf_0_i_clk),
    .Q(\mem[20][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09998_ (.D(_00306_),
    .CLK(clknet_leaf_1_i_clk),
    .Q(\mem[20][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09999_ (.D(_00307_),
    .CLK(clknet_leaf_1_i_clk),
    .Q(\mem[21][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10000_ (.D(_00308_),
    .CLK(clknet_leaf_2_i_clk),
    .Q(\mem[21][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10001_ (.D(_00309_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[21][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10002_ (.D(_00310_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[21][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10003_ (.D(_00311_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[21][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10004_ (.D(_00312_),
    .CLK(clknet_leaf_117_i_clk),
    .Q(\mem[21][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10005_ (.D(_00313_),
    .CLK(clknet_leaf_116_i_clk),
    .Q(\mem[21][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10006_ (.D(_00314_),
    .CLK(clknet_leaf_116_i_clk),
    .Q(\mem[21][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10007_ (.D(_00315_),
    .CLK(clknet_leaf_116_i_clk),
    .Q(\mem[21][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10008_ (.D(_00316_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[21][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10009_ (.D(_00317_),
    .CLK(clknet_leaf_116_i_clk),
    .Q(\mem[21][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10010_ (.D(_00318_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[21][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10011_ (.D(_00319_),
    .CLK(clknet_leaf_116_i_clk),
    .Q(\mem[21][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10012_ (.D(_00320_),
    .CLK(clknet_leaf_0_i_clk),
    .Q(\mem[21][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10013_ (.D(_00321_),
    .CLK(clknet_leaf_0_i_clk),
    .Q(\mem[21][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10014_ (.D(_00322_),
    .CLK(clknet_leaf_0_i_clk),
    .Q(\mem[21][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10015_ (.D(_00323_),
    .CLK(clknet_leaf_1_i_clk),
    .Q(\mem[22][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10016_ (.D(_00324_),
    .CLK(clknet_leaf_3_i_clk),
    .Q(\mem[22][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10017_ (.D(_00325_),
    .CLK(clknet_leaf_3_i_clk),
    .Q(\mem[22][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10018_ (.D(_00326_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[22][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10019_ (.D(_00327_),
    .CLK(clknet_leaf_118_i_clk),
    .Q(\mem[22][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10020_ (.D(_00328_),
    .CLK(clknet_leaf_117_i_clk),
    .Q(\mem[22][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10021_ (.D(_00329_),
    .CLK(clknet_leaf_117_i_clk),
    .Q(\mem[22][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10022_ (.D(_00330_),
    .CLK(clknet_leaf_116_i_clk),
    .Q(\mem[22][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10023_ (.D(_00331_),
    .CLK(clknet_leaf_116_i_clk),
    .Q(\mem[22][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10024_ (.D(_00332_),
    .CLK(clknet_leaf_115_i_clk),
    .Q(\mem[22][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10025_ (.D(_00333_),
    .CLK(clknet_leaf_116_i_clk),
    .Q(\mem[22][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10026_ (.D(_00334_),
    .CLK(clknet_leaf_116_i_clk),
    .Q(\mem[22][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10027_ (.D(_00335_),
    .CLK(clknet_leaf_114_i_clk),
    .Q(\mem[22][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10028_ (.D(_00336_),
    .CLK(clknet_leaf_114_i_clk),
    .Q(\mem[22][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10029_ (.D(_00337_),
    .CLK(clknet_leaf_113_i_clk),
    .Q(\mem[22][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10030_ (.D(_00338_),
    .CLK(clknet_leaf_0_i_clk),
    .Q(\mem[22][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10031_ (.D(_00339_),
    .CLK(clknet_leaf_106_i_clk),
    .Q(\mem[23][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10032_ (.D(_00340_),
    .CLK(clknet_leaf_105_i_clk),
    .Q(\mem[23][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10033_ (.D(_00341_),
    .CLK(clknet_leaf_106_i_clk),
    .Q(\mem[23][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10034_ (.D(_00342_),
    .CLK(clknet_leaf_106_i_clk),
    .Q(\mem[23][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10035_ (.D(_00343_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[23][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10036_ (.D(_00344_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[23][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10037_ (.D(_00345_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[23][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10038_ (.D(_00346_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[23][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10039_ (.D(_00347_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[23][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10040_ (.D(_00348_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[23][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10041_ (.D(_00349_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[23][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10042_ (.D(_00350_),
    .CLK(clknet_leaf_111_i_clk),
    .Q(\mem[23][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10043_ (.D(_00351_),
    .CLK(clknet_leaf_112_i_clk),
    .Q(\mem[23][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10044_ (.D(_00352_),
    .CLK(clknet_leaf_112_i_clk),
    .Q(\mem[23][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10045_ (.D(_00353_),
    .CLK(clknet_leaf_106_i_clk),
    .Q(\mem[23][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10046_ (.D(_00354_),
    .CLK(clknet_leaf_106_i_clk),
    .Q(\mem[23][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10047_ (.D(_00355_),
    .CLK(clknet_leaf_91_i_clk),
    .Q(\mem[24][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10048_ (.D(_00356_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[24][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10049_ (.D(_00357_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[24][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10050_ (.D(_00358_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[24][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10051_ (.D(_00359_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[24][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10052_ (.D(_00360_),
    .CLK(clknet_leaf_93_i_clk),
    .Q(\mem[24][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10053_ (.D(_00361_),
    .CLK(clknet_leaf_93_i_clk),
    .Q(\mem[24][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10054_ (.D(_00362_),
    .CLK(clknet_leaf_93_i_clk),
    .Q(\mem[24][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10055_ (.D(_00363_),
    .CLK(clknet_leaf_93_i_clk),
    .Q(\mem[24][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10056_ (.D(_00364_),
    .CLK(clknet_leaf_93_i_clk),
    .Q(\mem[24][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10057_ (.D(_00365_),
    .CLK(clknet_leaf_93_i_clk),
    .Q(\mem[24][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10058_ (.D(_00366_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[24][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10059_ (.D(_00367_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[24][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10060_ (.D(_00368_),
    .CLK(clknet_leaf_94_i_clk),
    .Q(\mem[24][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10061_ (.D(_00369_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[24][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10062_ (.D(_00370_),
    .CLK(clknet_leaf_98_i_clk),
    .Q(\mem[24][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10063_ (.D(_00371_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[25][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10064_ (.D(_00372_),
    .CLK(clknet_leaf_108_i_clk),
    .Q(\mem[25][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10065_ (.D(_00373_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[25][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10066_ (.D(_00374_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[25][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10067_ (.D(_00375_),
    .CLK(clknet_leaf_109_i_clk),
    .Q(\mem[25][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10068_ (.D(_00376_),
    .CLK(clknet_leaf_109_i_clk),
    .Q(\mem[25][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10069_ (.D(_00377_),
    .CLK(clknet_leaf_109_i_clk),
    .Q(\mem[25][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10070_ (.D(_00378_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[25][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10071_ (.D(_00379_),
    .CLK(clknet_leaf_109_i_clk),
    .Q(\mem[25][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10072_ (.D(_00380_),
    .CLK(clknet_leaf_109_i_clk),
    .Q(\mem[25][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10073_ (.D(_00381_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[25][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10074_ (.D(_00382_),
    .CLK(clknet_leaf_109_i_clk),
    .Q(\mem[25][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10075_ (.D(_00383_),
    .CLK(clknet_leaf_110_i_clk),
    .Q(\mem[25][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10076_ (.D(_00384_),
    .CLK(clknet_leaf_108_i_clk),
    .Q(\mem[25][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10077_ (.D(_00385_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[25][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10078_ (.D(_00386_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[25][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10079_ (.D(_00387_),
    .CLK(clknet_leaf_96_i_clk),
    .Q(\mem[26][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10080_ (.D(_00388_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[26][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10081_ (.D(_00389_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[26][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10082_ (.D(_00390_),
    .CLK(clknet_leaf_108_i_clk),
    .Q(\mem[26][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10083_ (.D(_00391_),
    .CLK(clknet_leaf_95_i_clk),
    .Q(\mem[26][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10084_ (.D(_00392_),
    .CLK(clknet_leaf_95_i_clk),
    .Q(\mem[26][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10085_ (.D(_00393_),
    .CLK(clknet_leaf_109_i_clk),
    .Q(\mem[26][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10086_ (.D(_00394_),
    .CLK(clknet_leaf_109_i_clk),
    .Q(\mem[26][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10087_ (.D(_00395_),
    .CLK(clknet_leaf_109_i_clk),
    .Q(\mem[26][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10088_ (.D(_00396_),
    .CLK(clknet_leaf_109_i_clk),
    .Q(\mem[26][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10089_ (.D(_00397_),
    .CLK(clknet_leaf_108_i_clk),
    .Q(\mem[26][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10090_ (.D(_00398_),
    .CLK(clknet_leaf_95_i_clk),
    .Q(\mem[26][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10091_ (.D(_00399_),
    .CLK(clknet_leaf_95_i_clk),
    .Q(\mem[26][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10092_ (.D(_00400_),
    .CLK(clknet_leaf_108_i_clk),
    .Q(\mem[26][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10093_ (.D(_00401_),
    .CLK(clknet_leaf_96_i_clk),
    .Q(\mem[26][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10094_ (.D(_00402_),
    .CLK(clknet_leaf_96_i_clk),
    .Q(\mem[26][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10095_ (.D(_00403_),
    .CLK(clknet_leaf_98_i_clk),
    .Q(\mem[27][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10096_ (.D(_00404_),
    .CLK(clknet_leaf_98_i_clk),
    .Q(\mem[27][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10097_ (.D(_00405_),
    .CLK(clknet_leaf_91_i_clk),
    .Q(\mem[27][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10098_ (.D(_00406_),
    .CLK(clknet_leaf_99_i_clk),
    .Q(\mem[27][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10099_ (.D(_00407_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[27][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10100_ (.D(_00408_),
    .CLK(clknet_leaf_99_i_clk),
    .Q(\mem[27][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10101_ (.D(_00409_),
    .CLK(clknet_leaf_99_i_clk),
    .Q(\mem[27][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10102_ (.D(_00410_),
    .CLK(clknet_leaf_99_i_clk),
    .Q(\mem[27][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10103_ (.D(_00411_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[27][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10104_ (.D(_00412_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[27][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10105_ (.D(_00413_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[27][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10106_ (.D(_00414_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[27][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10107_ (.D(_00415_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[27][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10108_ (.D(_00416_),
    .CLK(clknet_leaf_99_i_clk),
    .Q(\mem[27][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10109_ (.D(_00417_),
    .CLK(clknet_leaf_98_i_clk),
    .Q(\mem[27][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10110_ (.D(_00418_),
    .CLK(clknet_leaf_99_i_clk),
    .Q(\mem[27][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10111_ (.D(_00419_),
    .CLK(clknet_leaf_101_i_clk),
    .Q(\mem[28][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10112_ (.D(_00420_),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[28][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10113_ (.D(_00421_),
    .CLK(clknet_leaf_101_i_clk),
    .Q(\mem[28][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10114_ (.D(_00422_),
    .CLK(clknet_leaf_101_i_clk),
    .Q(\mem[28][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10115_ (.D(_00423_),
    .CLK(clknet_leaf_100_i_clk),
    .Q(\mem[28][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10116_ (.D(_00424_),
    .CLK(clknet_leaf_100_i_clk),
    .Q(\mem[28][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10117_ (.D(_00425_),
    .CLK(clknet_leaf_100_i_clk),
    .Q(\mem[28][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10118_ (.D(_00426_),
    .CLK(clknet_leaf_100_i_clk),
    .Q(\mem[28][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10119_ (.D(_00427_),
    .CLK(clknet_leaf_100_i_clk),
    .Q(\mem[28][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10120_ (.D(_00428_),
    .CLK(clknet_leaf_100_i_clk),
    .Q(\mem[28][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10121_ (.D(_00429_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[28][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10122_ (.D(_00430_),
    .CLK(clknet_leaf_99_i_clk),
    .Q(\mem[28][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10123_ (.D(_00431_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[28][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10124_ (.D(_00432_),
    .CLK(clknet_leaf_72_i_clk),
    .Q(\mem[28][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10125_ (.D(_00433_),
    .CLK(clknet_leaf_101_i_clk),
    .Q(\mem[28][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10126_ (.D(_00434_),
    .CLK(clknet_leaf_100_i_clk),
    .Q(\mem[28][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10127_ (.D(_00435_),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[2][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10128_ (.D(_00436_),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[2][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10129_ (.D(_00437_),
    .CLK(clknet_leaf_103_i_clk),
    .Q(\mem[2][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10130_ (.D(_00438_),
    .CLK(clknet_leaf_103_i_clk),
    .Q(\mem[2][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10131_ (.D(_00439_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[2][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10132_ (.D(_00440_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[2][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10133_ (.D(_00441_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[2][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10134_ (.D(_00442_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[2][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10135_ (.D(_00443_),
    .CLK(clknet_leaf_104_i_clk),
    .Q(\mem[2][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10136_ (.D(_00444_),
    .CLK(clknet_leaf_103_i_clk),
    .Q(\mem[2][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10137_ (.D(_00445_),
    .CLK(clknet_leaf_103_i_clk),
    .Q(\mem[2][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10138_ (.D(_00446_),
    .CLK(clknet_leaf_103_i_clk),
    .Q(\mem[2][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10139_ (.D(_00447_),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[2][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10140_ (.D(_00448_),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[2][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10141_ (.D(_00449_),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[2][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10142_ (.D(_00450_),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[2][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10143_ (.D(_00451_),
    .CLK(clknet_leaf_96_i_clk),
    .Q(\mem[30][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10144_ (.D(_00452_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[30][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10145_ (.D(_00453_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[30][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10146_ (.D(_00454_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[30][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10147_ (.D(_00455_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[30][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10148_ (.D(_00456_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[30][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10149_ (.D(_00457_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[30][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10150_ (.D(_00458_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[30][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10151_ (.D(_00459_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[30][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10152_ (.D(_00460_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[30][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10153_ (.D(_00461_),
    .CLK(clknet_leaf_107_i_clk),
    .Q(\mem[30][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10154_ (.D(_00462_),
    .CLK(clknet_leaf_97_i_clk),
    .Q(\mem[30][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10155_ (.D(_00463_),
    .CLK(clknet_leaf_96_i_clk),
    .Q(\mem[30][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10156_ (.D(_00464_),
    .CLK(clknet_leaf_97_i_clk),
    .Q(\mem[30][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10157_ (.D(_00465_),
    .CLK(clknet_leaf_97_i_clk),
    .Q(\mem[30][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10158_ (.D(_00466_),
    .CLK(clknet_leaf_97_i_clk),
    .Q(\mem[30][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10159_ (.D(_00467_),
    .CLK(clknet_leaf_96_i_clk),
    .Q(\mem[31][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10160_ (.D(_00468_),
    .CLK(clknet_leaf_95_i_clk),
    .Q(\mem[31][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10161_ (.D(_00469_),
    .CLK(clknet_leaf_96_i_clk),
    .Q(\mem[31][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10162_ (.D(_00470_),
    .CLK(clknet_leaf_95_i_clk),
    .Q(\mem[31][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10163_ (.D(_00471_),
    .CLK(clknet_leaf_95_i_clk),
    .Q(\mem[31][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10164_ (.D(_00472_),
    .CLK(clknet_leaf_95_i_clk),
    .Q(\mem[31][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10165_ (.D(_00473_),
    .CLK(clknet_leaf_95_i_clk),
    .Q(\mem[31][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10166_ (.D(_00474_),
    .CLK(clknet_leaf_94_i_clk),
    .Q(\mem[31][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10167_ (.D(_00475_),
    .CLK(clknet_leaf_94_i_clk),
    .Q(\mem[31][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10168_ (.D(_00476_),
    .CLK(clknet_leaf_94_i_clk),
    .Q(\mem[31][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10169_ (.D(_00477_),
    .CLK(clknet_leaf_94_i_clk),
    .Q(\mem[31][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10170_ (.D(_00478_),
    .CLK(clknet_leaf_94_i_clk),
    .Q(\mem[31][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10171_ (.D(_00479_),
    .CLK(clknet_leaf_96_i_clk),
    .Q(\mem[31][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10172_ (.D(_00480_),
    .CLK(clknet_leaf_94_i_clk),
    .Q(\mem[31][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10173_ (.D(_00481_),
    .CLK(clknet_leaf_96_i_clk),
    .Q(\mem[31][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10174_ (.D(_00482_),
    .CLK(clknet_leaf_97_i_clk),
    .Q(\mem[31][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10175_ (.D(_00483_),
    .CLK(clknet_leaf_91_i_clk),
    .Q(\mem[32][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10176_ (.D(_00484_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[32][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10177_ (.D(_00485_),
    .CLK(clknet_leaf_91_i_clk),
    .Q(\mem[32][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10178_ (.D(_00486_),
    .CLK(clknet_leaf_91_i_clk),
    .Q(\mem[32][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10179_ (.D(_00487_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[32][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10180_ (.D(_00488_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[32][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10181_ (.D(_00489_),
    .CLK(clknet_leaf_92_i_clk),
    .Q(\mem[32][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10182_ (.D(_00490_),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[32][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10183_ (.D(_00491_),
    .CLK(clknet_leaf_93_i_clk),
    .Q(\mem[32][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10184_ (.D(_00492_),
    .CLK(clknet_leaf_93_i_clk),
    .Q(\mem[32][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10185_ (.D(_00493_),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[32][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10186_ (.D(_00494_),
    .CLK(clknet_leaf_93_i_clk),
    .Q(\mem[32][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10187_ (.D(_00495_),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[32][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10188_ (.D(_00496_),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[32][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10189_ (.D(_00497_),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[32][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10190_ (.D(_00498_),
    .CLK(clknet_leaf_91_i_clk),
    .Q(\mem[32][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10191_ (.D(_00499_),
    .CLK(clknet_leaf_90_i_clk),
    .Q(\mem[33][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10192_ (.D(_00500_),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[33][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10193_ (.D(_00501_),
    .CLK(clknet_leaf_86_i_clk),
    .Q(\mem[33][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10194_ (.D(_00502_),
    .CLK(clknet_leaf_90_i_clk),
    .Q(\mem[33][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10195_ (.D(_00503_),
    .CLK(clknet_leaf_86_i_clk),
    .Q(\mem[33][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10196_ (.D(_00504_),
    .CLK(clknet_leaf_86_i_clk),
    .Q(\mem[33][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10197_ (.D(_00505_),
    .CLK(clknet_leaf_86_i_clk),
    .Q(\mem[33][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10198_ (.D(_00506_),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[33][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10199_ (.D(_00507_),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[33][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10200_ (.D(_00508_),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[33][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10201_ (.D(_00509_),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[33][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10202_ (.D(_00510_),
    .CLK(clknet_leaf_88_i_clk),
    .Q(\mem[33][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10203_ (.D(_00511_),
    .CLK(clknet_leaf_88_i_clk),
    .Q(\mem[33][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10204_ (.D(_00512_),
    .CLK(clknet_leaf_88_i_clk),
    .Q(\mem[33][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10205_ (.D(_00513_),
    .CLK(clknet_leaf_90_i_clk),
    .Q(\mem[33][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10206_ (.D(_00514_),
    .CLK(clknet_leaf_90_i_clk),
    .Q(\mem[33][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10207_ (.D(_00515_),
    .CLK(clknet_leaf_90_i_clk),
    .Q(\mem[34][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10208_ (.D(_00516_),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[34][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10209_ (.D(_00517_),
    .CLK(clknet_leaf_84_i_clk),
    .Q(\mem[34][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10210_ (.D(_00518_),
    .CLK(clknet_leaf_88_i_clk),
    .Q(\mem[34][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10211_ (.D(_00519_),
    .CLK(clknet_leaf_88_i_clk),
    .Q(\mem[34][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10212_ (.D(_00520_),
    .CLK(clknet_leaf_86_i_clk),
    .Q(\mem[34][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10213_ (.D(_00521_),
    .CLK(clknet_leaf_85_i_clk),
    .Q(\mem[34][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10214_ (.D(_00522_),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[34][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10215_ (.D(_00523_),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[34][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10216_ (.D(_00524_),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[34][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10217_ (.D(_00525_),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[34][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10218_ (.D(_00526_),
    .CLK(clknet_leaf_88_i_clk),
    .Q(\mem[34][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10219_ (.D(_00527_),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[34][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10220_ (.D(_00528_),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[34][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10221_ (.D(_00529_),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[34][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10222_ (.D(_00530_),
    .CLK(clknet_leaf_90_i_clk),
    .Q(\mem[34][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10223_ (.D(_00531_),
    .CLK(clknet_leaf_90_i_clk),
    .Q(\mem[35][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10224_ (.D(_00532_),
    .CLK(clknet_leaf_91_i_clk),
    .Q(\mem[35][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10225_ (.D(_00533_),
    .CLK(clknet_leaf_84_i_clk),
    .Q(\mem[35][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10226_ (.D(_00534_),
    .CLK(clknet_leaf_83_i_clk),
    .Q(\mem[35][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10227_ (.D(_00535_),
    .CLK(clknet_leaf_84_i_clk),
    .Q(\mem[35][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10228_ (.D(_00536_),
    .CLK(clknet_leaf_85_i_clk),
    .Q(\mem[35][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10229_ (.D(_00537_),
    .CLK(clknet_leaf_85_i_clk),
    .Q(\mem[35][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10230_ (.D(_00538_),
    .CLK(clknet_leaf_85_i_clk),
    .Q(\mem[35][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10231_ (.D(_00539_),
    .CLK(clknet_leaf_85_i_clk),
    .Q(\mem[35][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10232_ (.D(_00540_),
    .CLK(clknet_leaf_84_i_clk),
    .Q(\mem[35][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10233_ (.D(_00541_),
    .CLK(clknet_leaf_84_i_clk),
    .Q(\mem[35][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10234_ (.D(_00542_),
    .CLK(clknet_leaf_83_i_clk),
    .Q(\mem[35][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10235_ (.D(_00543_),
    .CLK(clknet_leaf_83_i_clk),
    .Q(\mem[35][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10236_ (.D(_00544_),
    .CLK(clknet_leaf_83_i_clk),
    .Q(\mem[35][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10237_ (.D(_00545_),
    .CLK(clknet_leaf_83_i_clk),
    .Q(\mem[35][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10238_ (.D(_00546_),
    .CLK(clknet_leaf_83_i_clk),
    .Q(\mem[35][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10239_ (.D(_00547_),
    .CLK(clknet_leaf_75_i_clk),
    .Q(\mem[36][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10240_ (.D(_00548_),
    .CLK(clknet_leaf_75_i_clk),
    .Q(\mem[36][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10241_ (.D(_00549_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[36][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10242_ (.D(_00550_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[36][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10243_ (.D(_00551_),
    .CLK(clknet_leaf_81_i_clk),
    .Q(\mem[36][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10244_ (.D(_00552_),
    .CLK(clknet_leaf_81_i_clk),
    .Q(\mem[36][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10245_ (.D(_00553_),
    .CLK(clknet_leaf_85_i_clk),
    .Q(\mem[36][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10246_ (.D(_00554_),
    .CLK(clknet_leaf_85_i_clk),
    .Q(\mem[36][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10247_ (.D(_00555_),
    .CLK(clknet_leaf_81_i_clk),
    .Q(\mem[36][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10248_ (.D(_00556_),
    .CLK(clknet_leaf_81_i_clk),
    .Q(\mem[36][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10249_ (.D(_00557_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[36][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10250_ (.D(_00558_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[36][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10251_ (.D(_00559_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[36][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10252_ (.D(_00560_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[36][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10253_ (.D(_00561_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[36][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10254_ (.D(_00562_),
    .CLK(clknet_leaf_75_i_clk),
    .Q(\mem[36][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10255_ (.D(_00563_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[37][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10256_ (.D(_00564_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[37][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10257_ (.D(_00565_),
    .CLK(clknet_leaf_78_i_clk),
    .Q(\mem[37][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10258_ (.D(_00566_),
    .CLK(clknet_leaf_78_i_clk),
    .Q(\mem[37][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10259_ (.D(_00567_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[37][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10260_ (.D(_00568_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[37][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10261_ (.D(_00569_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[37][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10262_ (.D(_00570_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[37][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10263_ (.D(_00571_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[37][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10264_ (.D(_00572_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[37][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10265_ (.D(_00573_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[37][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10266_ (.D(_00574_),
    .CLK(clknet_leaf_76_i_clk),
    .Q(\mem[37][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10267_ (.D(_00575_),
    .CLK(clknet_leaf_76_i_clk),
    .Q(\mem[37][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10268_ (.D(_00576_),
    .CLK(clknet_leaf_76_i_clk),
    .Q(\mem[37][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10269_ (.D(_00577_),
    .CLK(clknet_leaf_76_i_clk),
    .Q(\mem[37][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10270_ (.D(_00578_),
    .CLK(clknet_leaf_76_i_clk),
    .Q(\mem[37][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10271_ (.D(_00579_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[38][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10272_ (.D(_00580_),
    .CLK(clknet_leaf_74_i_clk),
    .Q(\mem[38][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10273_ (.D(_00581_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[38][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10274_ (.D(_00582_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[38][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10275_ (.D(_00583_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[38][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10276_ (.D(_00584_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[38][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10277_ (.D(_00585_),
    .CLK(clknet_leaf_81_i_clk),
    .Q(\mem[38][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10278_ (.D(_00586_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[38][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10279_ (.D(_00587_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(\mem[38][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10280_ (.D(_00588_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[38][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10281_ (.D(_00589_),
    .CLK(clknet_leaf_82_i_clk),
    .Q(\mem[38][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10282_ (.D(_00590_),
    .CLK(clknet_leaf_76_i_clk),
    .Q(\mem[38][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10283_ (.D(_00591_),
    .CLK(clknet_leaf_76_i_clk),
    .Q(\mem[38][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10284_ (.D(_00592_),
    .CLK(clknet_leaf_75_i_clk),
    .Q(\mem[38][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10285_ (.D(_00593_),
    .CLK(clknet_leaf_75_i_clk),
    .Q(\mem[38][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10286_ (.D(_00594_),
    .CLK(clknet_leaf_75_i_clk),
    .Q(\mem[38][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10287_ (.D(_00595_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[3][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10288_ (.D(_00596_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[3][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10289_ (.D(_00597_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[3][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10290_ (.D(_00598_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[3][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10291_ (.D(_00599_),
    .CLK(clknet_leaf_66_i_clk),
    .Q(\mem[3][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10292_ (.D(_00600_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[3][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10293_ (.D(_00601_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[3][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10294_ (.D(_00602_),
    .CLK(clknet_leaf_66_i_clk),
    .Q(\mem[3][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10295_ (.D(_00603_),
    .CLK(clknet_leaf_69_i_clk),
    .Q(\mem[3][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10296_ (.D(_00604_),
    .CLK(clknet_leaf_69_i_clk),
    .Q(\mem[3][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10297_ (.D(_00605_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[3][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10298_ (.D(_00606_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[3][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10299_ (.D(_00607_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[3][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10300_ (.D(_00608_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[3][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10301_ (.D(_00609_),
    .CLK(clknet_leaf_72_i_clk),
    .Q(\mem[3][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10302_ (.D(_00610_),
    .CLK(clknet_leaf_73_i_clk),
    .Q(\mem[3][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10303_ (.D(_00611_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[40][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10304_ (.D(_00612_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[40][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10305_ (.D(_00613_),
    .CLK(clknet_leaf_78_i_clk),
    .Q(\mem[40][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10306_ (.D(_00614_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[40][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10307_ (.D(_00615_),
    .CLK(clknet_leaf_64_i_clk),
    .Q(\mem[40][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10308_ (.D(_00616_),
    .CLK(clknet_leaf_79_i_clk),
    .Q(\mem[40][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10309_ (.D(_00617_),
    .CLK(clknet_leaf_64_i_clk),
    .Q(\mem[40][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10310_ (.D(_00618_),
    .CLK(clknet_leaf_63_i_clk),
    .Q(\mem[40][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10311_ (.D(_00619_),
    .CLK(clknet_leaf_63_i_clk),
    .Q(\mem[40][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10312_ (.D(_00620_),
    .CLK(clknet_leaf_63_i_clk),
    .Q(\mem[40][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10313_ (.D(_00621_),
    .CLK(clknet_leaf_64_i_clk),
    .Q(\mem[40][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10314_ (.D(_00622_),
    .CLK(clknet_leaf_65_i_clk),
    .Q(\mem[40][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10315_ (.D(_00623_),
    .CLK(clknet_leaf_66_i_clk),
    .Q(\mem[40][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10316_ (.D(_00624_),
    .CLK(clknet_leaf_65_i_clk),
    .Q(\mem[40][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10317_ (.D(_00625_),
    .CLK(clknet_leaf_66_i_clk),
    .Q(\mem[40][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10318_ (.D(_00626_),
    .CLK(clknet_leaf_66_i_clk),
    .Q(\mem[40][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10319_ (.D(_00627_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[41][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10320_ (.D(_00628_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[41][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10321_ (.D(_00629_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[41][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10322_ (.D(_00630_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[41][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10323_ (.D(_00631_),
    .CLK(clknet_leaf_79_i_clk),
    .Q(\mem[41][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10324_ (.D(_00632_),
    .CLK(clknet_leaf_79_i_clk),
    .Q(\mem[41][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10325_ (.D(_00633_),
    .CLK(clknet_leaf_79_i_clk),
    .Q(\mem[41][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10326_ (.D(_00634_),
    .CLK(clknet_leaf_64_i_clk),
    .Q(\mem[41][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10327_ (.D(_00635_),
    .CLK(clknet_leaf_63_i_clk),
    .Q(\mem[41][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10328_ (.D(_00636_),
    .CLK(clknet_leaf_64_i_clk),
    .Q(\mem[41][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10329_ (.D(_00637_),
    .CLK(clknet_leaf_65_i_clk),
    .Q(\mem[41][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10330_ (.D(_00638_),
    .CLK(clknet_leaf_65_i_clk),
    .Q(\mem[41][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10331_ (.D(_00639_),
    .CLK(clknet_leaf_65_i_clk),
    .Q(\mem[41][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10332_ (.D(_00640_),
    .CLK(clknet_leaf_65_i_clk),
    .Q(\mem[41][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10333_ (.D(_00641_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[41][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10334_ (.D(_00642_),
    .CLK(clknet_leaf_66_i_clk),
    .Q(\mem[41][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10335_ (.D(_00643_),
    .CLK(clknet_leaf_76_i_clk),
    .Q(\mem[42][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10336_ (.D(_00644_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[42][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10337_ (.D(_00645_),
    .CLK(clknet_leaf_78_i_clk),
    .Q(\mem[42][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10338_ (.D(_00646_),
    .CLK(clknet_leaf_77_i_clk),
    .Q(\mem[42][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10339_ (.D(_00647_),
    .CLK(clknet_leaf_78_i_clk),
    .Q(\mem[42][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10340_ (.D(_00648_),
    .CLK(clknet_leaf_79_i_clk),
    .Q(\mem[42][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10341_ (.D(_00649_),
    .CLK(clknet_leaf_79_i_clk),
    .Q(\mem[42][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10342_ (.D(_00650_),
    .CLK(clknet_leaf_64_i_clk),
    .Q(\mem[42][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10343_ (.D(_00651_),
    .CLK(clknet_leaf_63_i_clk),
    .Q(\mem[42][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10344_ (.D(_00652_),
    .CLK(clknet_leaf_63_i_clk),
    .Q(\mem[42][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10345_ (.D(_00653_),
    .CLK(clknet_leaf_64_i_clk),
    .Q(\mem[42][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10346_ (.D(_00654_),
    .CLK(clknet_leaf_63_i_clk),
    .Q(\mem[42][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10347_ (.D(_00655_),
    .CLK(clknet_leaf_65_i_clk),
    .Q(\mem[42][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10348_ (.D(_00656_),
    .CLK(clknet_leaf_66_i_clk),
    .Q(\mem[42][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10349_ (.D(_00657_),
    .CLK(clknet_leaf_66_i_clk),
    .Q(\mem[42][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10350_ (.D(_00658_),
    .CLK(clknet_leaf_66_i_clk),
    .Q(\mem[42][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10351_ (.D(_00659_),
    .CLK(clknet_leaf_59_i_clk),
    .Q(\mem[43][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10352_ (.D(_00660_),
    .CLK(clknet_leaf_59_i_clk),
    .Q(\mem[43][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10353_ (.D(_00661_),
    .CLK(clknet_leaf_58_i_clk),
    .Q(\mem[43][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10354_ (.D(_00662_),
    .CLK(clknet_leaf_59_i_clk),
    .Q(\mem[43][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10355_ (.D(_00663_),
    .CLK(clknet_leaf_57_i_clk),
    .Q(\mem[43][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10356_ (.D(_00664_),
    .CLK(clknet_leaf_57_i_clk),
    .Q(\mem[43][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10357_ (.D(_00665_),
    .CLK(clknet_leaf_57_i_clk),
    .Q(\mem[43][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10358_ (.D(_00666_),
    .CLK(clknet_leaf_57_i_clk),
    .Q(\mem[43][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10359_ (.D(_00667_),
    .CLK(clknet_leaf_57_i_clk),
    .Q(\mem[43][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10360_ (.D(_00668_),
    .CLK(clknet_leaf_57_i_clk),
    .Q(\mem[43][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10361_ (.D(_00669_),
    .CLK(clknet_leaf_58_i_clk),
    .Q(\mem[43][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10362_ (.D(_00670_),
    .CLK(clknet_leaf_59_i_clk),
    .Q(\mem[43][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10363_ (.D(_00671_),
    .CLK(clknet_leaf_59_i_clk),
    .Q(\mem[43][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10364_ (.D(_00672_),
    .CLK(clknet_leaf_59_i_clk),
    .Q(\mem[43][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10365_ (.D(_00673_),
    .CLK(clknet_leaf_52_i_clk),
    .Q(\mem[43][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10366_ (.D(_00674_),
    .CLK(clknet_leaf_52_i_clk),
    .Q(\mem[43][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10367_ (.D(_00675_),
    .CLK(clknet_leaf_60_i_clk),
    .Q(\mem[44][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10368_ (.D(_00676_),
    .CLK(clknet_leaf_60_i_clk),
    .Q(\mem[44][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10369_ (.D(_00677_),
    .CLK(clknet_leaf_61_i_clk),
    .Q(\mem[44][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10370_ (.D(_00678_),
    .CLK(clknet_leaf_61_i_clk),
    .Q(\mem[44][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10371_ (.D(_00679_),
    .CLK(clknet_leaf_58_i_clk),
    .Q(\mem[44][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10372_ (.D(_00680_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(\mem[44][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10373_ (.D(_00681_),
    .CLK(clknet_leaf_58_i_clk),
    .Q(\mem[44][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10374_ (.D(_00682_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(\mem[44][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10375_ (.D(_00683_),
    .CLK(clknet_leaf_61_i_clk),
    .Q(\mem[44][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10376_ (.D(_00684_),
    .CLK(clknet_leaf_61_i_clk),
    .Q(\mem[44][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10377_ (.D(_00685_),
    .CLK(clknet_leaf_61_i_clk),
    .Q(\mem[44][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10378_ (.D(_00686_),
    .CLK(clknet_leaf_60_i_clk),
    .Q(\mem[44][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10379_ (.D(_00687_),
    .CLK(clknet_leaf_60_i_clk),
    .Q(\mem[44][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10380_ (.D(_00688_),
    .CLK(clknet_leaf_60_i_clk),
    .Q(\mem[44][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10381_ (.D(_00689_),
    .CLK(clknet_leaf_60_i_clk),
    .Q(\mem[44][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10382_ (.D(_00690_),
    .CLK(clknet_leaf_60_i_clk),
    .Q(\mem[44][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10383_ (.D(_00691_),
    .CLK(clknet_leaf_53_i_clk),
    .Q(\mem[45][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10384_ (.D(_00692_),
    .CLK(clknet_leaf_53_i_clk),
    .Q(\mem[45][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10385_ (.D(_00693_),
    .CLK(clknet_leaf_55_i_clk),
    .Q(\mem[45][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10386_ (.D(_00694_),
    .CLK(clknet_leaf_59_i_clk),
    .Q(\mem[45][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10387_ (.D(_00695_),
    .CLK(clknet_leaf_55_i_clk),
    .Q(\mem[45][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10388_ (.D(_00696_),
    .CLK(clknet_leaf_56_i_clk),
    .Q(\mem[45][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10389_ (.D(_00697_),
    .CLK(clknet_leaf_56_i_clk),
    .Q(\mem[45][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10390_ (.D(_00698_),
    .CLK(clknet_leaf_56_i_clk),
    .Q(\mem[45][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10391_ (.D(_00699_),
    .CLK(clknet_leaf_55_i_clk),
    .Q(\mem[45][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10392_ (.D(_00700_),
    .CLK(clknet_leaf_55_i_clk),
    .Q(\mem[45][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10393_ (.D(_00701_),
    .CLK(clknet_leaf_55_i_clk),
    .Q(\mem[45][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10394_ (.D(_00702_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[45][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10395_ (.D(_00703_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[45][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10396_ (.D(_00704_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[45][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10397_ (.D(_00705_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[45][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10398_ (.D(_00706_),
    .CLK(clknet_leaf_53_i_clk),
    .Q(\mem[45][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10399_ (.D(_00707_),
    .CLK(clknet_leaf_53_i_clk),
    .Q(\mem[46][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10400_ (.D(_00708_),
    .CLK(clknet_leaf_53_i_clk),
    .Q(\mem[46][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10401_ (.D(_00709_),
    .CLK(clknet_leaf_55_i_clk),
    .Q(\mem[46][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10402_ (.D(_00710_),
    .CLK(clknet_leaf_57_i_clk),
    .Q(\mem[46][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10403_ (.D(_00711_),
    .CLK(clknet_leaf_56_i_clk),
    .Q(\mem[46][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10404_ (.D(_00712_),
    .CLK(clknet_leaf_56_i_clk),
    .Q(\mem[46][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10405_ (.D(_00713_),
    .CLK(clknet_leaf_56_i_clk),
    .Q(\mem[46][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10406_ (.D(_00714_),
    .CLK(clknet_leaf_55_i_clk),
    .Q(\mem[46][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10407_ (.D(_00715_),
    .CLK(clknet_leaf_55_i_clk),
    .Q(\mem[46][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10408_ (.D(_00716_),
    .CLK(clknet_leaf_55_i_clk),
    .Q(\mem[46][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10409_ (.D(_00717_),
    .CLK(clknet_leaf_55_i_clk),
    .Q(\mem[46][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10410_ (.D(_00718_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[46][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10411_ (.D(_00719_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[46][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10412_ (.D(_00720_),
    .CLK(clknet_leaf_53_i_clk),
    .Q(\mem[46][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10413_ (.D(_00721_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[46][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10414_ (.D(_00722_),
    .CLK(clknet_leaf_53_i_clk),
    .Q(\mem[46][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10415_ (.D(_00723_),
    .CLK(clknet_leaf_67_i_clk),
    .Q(\mem[47][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10416_ (.D(_00724_),
    .CLK(clknet_leaf_67_i_clk),
    .Q(\mem[47][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10417_ (.D(_00725_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(\mem[47][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10418_ (.D(_00726_),
    .CLK(clknet_leaf_61_i_clk),
    .Q(\mem[47][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10419_ (.D(_00727_),
    .CLK(clknet_leaf_61_i_clk),
    .Q(\mem[47][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10420_ (.D(_00728_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(\mem[47][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10421_ (.D(_00729_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(\mem[47][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10422_ (.D(_00730_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(\mem[47][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10423_ (.D(_00731_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(\mem[47][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10424_ (.D(_00732_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(\mem[47][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10425_ (.D(_00733_),
    .CLK(clknet_leaf_61_i_clk),
    .Q(\mem[47][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10426_ (.D(_00734_),
    .CLK(clknet_leaf_60_i_clk),
    .Q(\mem[47][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10427_ (.D(_00735_),
    .CLK(clknet_leaf_67_i_clk),
    .Q(\mem[47][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10428_ (.D(_00736_),
    .CLK(clknet_leaf_60_i_clk),
    .Q(\mem[47][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10429_ (.D(_00737_),
    .CLK(clknet_leaf_67_i_clk),
    .Q(\mem[47][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10430_ (.D(_00738_),
    .CLK(clknet_leaf_67_i_clk),
    .Q(\mem[47][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10431_ (.D(_00739_),
    .CLK(clknet_leaf_69_i_clk),
    .Q(\mem[48][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10432_ (.D(_00740_),
    .CLK(clknet_leaf_69_i_clk),
    .Q(\mem[48][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10433_ (.D(_00741_),
    .CLK(clknet_leaf_51_i_clk),
    .Q(\mem[48][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10434_ (.D(_00742_),
    .CLK(clknet_leaf_51_i_clk),
    .Q(\mem[48][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10435_ (.D(_00743_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[48][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10436_ (.D(_00744_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[48][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10437_ (.D(_00745_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[48][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10438_ (.D(_00746_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[48][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10439_ (.D(_00747_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[48][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10440_ (.D(_00748_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[48][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10441_ (.D(_00749_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[48][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10442_ (.D(_00750_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[48][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10443_ (.D(_00751_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[48][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10444_ (.D(_00752_),
    .CLK(clknet_leaf_46_i_clk),
    .Q(\mem[48][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10445_ (.D(_00753_),
    .CLK(clknet_leaf_51_i_clk),
    .Q(\mem[48][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10446_ (.D(_00754_),
    .CLK(clknet_leaf_45_i_clk),
    .Q(\mem[48][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10447_ (.D(_00755_),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[4][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10448_ (.D(_00756_),
    .CLK(clknet_leaf_66_i_clk),
    .Q(\mem[4][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10449_ (.D(_00757_),
    .CLK(clknet_leaf_67_i_clk),
    .Q(\mem[4][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10450_ (.D(_00758_),
    .CLK(clknet_leaf_69_i_clk),
    .Q(\mem[4][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10451_ (.D(_00759_),
    .CLK(clknet_leaf_67_i_clk),
    .Q(\mem[4][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10452_ (.D(_00760_),
    .CLK(clknet_leaf_67_i_clk),
    .Q(\mem[4][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10453_ (.D(_00761_),
    .CLK(clknet_leaf_68_i_clk),
    .Q(\mem[4][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10454_ (.D(_00762_),
    .CLK(clknet_leaf_68_i_clk),
    .Q(\mem[4][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10455_ (.D(_00763_),
    .CLK(clknet_leaf_68_i_clk),
    .Q(\mem[4][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10456_ (.D(_00764_),
    .CLK(clknet_leaf_68_i_clk),
    .Q(\mem[4][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10457_ (.D(_00765_),
    .CLK(clknet_leaf_69_i_clk),
    .Q(\mem[4][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10458_ (.D(_00766_),
    .CLK(clknet_leaf_68_i_clk),
    .Q(\mem[4][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10459_ (.D(_00767_),
    .CLK(clknet_leaf_69_i_clk),
    .Q(\mem[4][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10460_ (.D(_00768_),
    .CLK(clknet_leaf_69_i_clk),
    .Q(\mem[4][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10461_ (.D(_00769_),
    .CLK(clknet_leaf_69_i_clk),
    .Q(\mem[4][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10462_ (.D(_00770_),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[4][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10463_ (.D(_00771_),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[50][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10464_ (.D(_00772_),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[50][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10465_ (.D(_00773_),
    .CLK(clknet_leaf_68_i_clk),
    .Q(\mem[50][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10466_ (.D(_00774_),
    .CLK(clknet_leaf_44_i_clk),
    .Q(\mem[50][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10467_ (.D(_00775_),
    .CLK(clknet_leaf_44_i_clk),
    .Q(\mem[50][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10468_ (.D(_00776_),
    .CLK(clknet_leaf_68_i_clk),
    .Q(\mem[50][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10469_ (.D(_00777_),
    .CLK(clknet_leaf_45_i_clk),
    .Q(\mem[50][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10470_ (.D(_00778_),
    .CLK(clknet_leaf_45_i_clk),
    .Q(\mem[50][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10471_ (.D(_00779_),
    .CLK(clknet_leaf_45_i_clk),
    .Q(\mem[50][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10472_ (.D(_00780_),
    .CLK(clknet_leaf_45_i_clk),
    .Q(\mem[50][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10473_ (.D(_00781_),
    .CLK(clknet_leaf_45_i_clk),
    .Q(\mem[50][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10474_ (.D(_00782_),
    .CLK(clknet_leaf_45_i_clk),
    .Q(\mem[50][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10475_ (.D(_00783_),
    .CLK(clknet_leaf_43_i_clk),
    .Q(\mem[50][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10476_ (.D(_00784_),
    .CLK(clknet_leaf_46_i_clk),
    .Q(\mem[50][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10477_ (.D(_00785_),
    .CLK(clknet_leaf_45_i_clk),
    .Q(\mem[50][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10478_ (.D(_00786_),
    .CLK(clknet_leaf_45_i_clk),
    .Q(\mem[50][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10479_ (.D(_00787_),
    .CLK(clknet_leaf_45_i_clk),
    .Q(\mem[51][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10480_ (.D(_00788_),
    .CLK(clknet_leaf_52_i_clk),
    .Q(\mem[51][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10481_ (.D(_00789_),
    .CLK(clknet_leaf_52_i_clk),
    .Q(\mem[51][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10482_ (.D(_00790_),
    .CLK(clknet_leaf_52_i_clk),
    .Q(\mem[51][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10483_ (.D(_00791_),
    .CLK(clknet_leaf_52_i_clk),
    .Q(\mem[51][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10484_ (.D(_00792_),
    .CLK(clknet_leaf_53_i_clk),
    .Q(\mem[51][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10485_ (.D(_00793_),
    .CLK(clknet_leaf_53_i_clk),
    .Q(\mem[51][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10486_ (.D(_00794_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[51][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10487_ (.D(_00795_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[51][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10488_ (.D(_00796_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[51][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10489_ (.D(_00797_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[51][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10490_ (.D(_00798_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[51][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10491_ (.D(_00799_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[51][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10492_ (.D(_00800_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[51][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10493_ (.D(_00801_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[51][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10494_ (.D(_00802_),
    .CLK(clknet_leaf_51_i_clk),
    .Q(\mem[51][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10495_ (.D(_00803_),
    .CLK(clknet_leaf_51_i_clk),
    .Q(\mem[52][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10496_ (.D(_00804_),
    .CLK(clknet_leaf_51_i_clk),
    .Q(\mem[52][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10497_ (.D(_00805_),
    .CLK(clknet_leaf_51_i_clk),
    .Q(\mem[52][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10498_ (.D(_00806_),
    .CLK(clknet_leaf_51_i_clk),
    .Q(\mem[52][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10499_ (.D(_00807_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[52][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10500_ (.D(_00808_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[52][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10501_ (.D(_00809_),
    .CLK(clknet_leaf_51_i_clk),
    .Q(\mem[52][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10502_ (.D(_00810_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[52][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10503_ (.D(_00811_),
    .CLK(clknet_leaf_54_i_clk),
    .Q(\mem[52][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10504_ (.D(_00812_),
    .CLK(clknet_leaf_50_i_clk),
    .Q(\mem[52][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10505_ (.D(_00813_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[52][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10506_ (.D(_00814_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[52][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10507_ (.D(_00815_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[52][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10508_ (.D(_00816_),
    .CLK(clknet_leaf_49_i_clk),
    .Q(\mem[52][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10509_ (.D(_00817_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[52][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10510_ (.D(_00818_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[52][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10511_ (.D(_00819_),
    .CLK(clknet_leaf_36_i_clk),
    .Q(\mem[53][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10512_ (.D(_00820_),
    .CLK(clknet_leaf_36_i_clk),
    .Q(\mem[53][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10513_ (.D(_00821_),
    .CLK(clknet_leaf_36_i_clk),
    .Q(\mem[53][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10514_ (.D(_00822_),
    .CLK(clknet_leaf_35_i_clk),
    .Q(\mem[53][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10515_ (.D(_00823_),
    .CLK(clknet_leaf_33_i_clk),
    .Q(\mem[53][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10516_ (.D(_00824_),
    .CLK(clknet_leaf_35_i_clk),
    .Q(\mem[53][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10517_ (.D(_00825_),
    .CLK(clknet_leaf_34_i_clk),
    .Q(\mem[53][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10518_ (.D(_00826_),
    .CLK(clknet_leaf_33_i_clk),
    .Q(\mem[53][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10519_ (.D(_00827_),
    .CLK(clknet_leaf_33_i_clk),
    .Q(\mem[53][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10520_ (.D(_00828_),
    .CLK(clknet_leaf_33_i_clk),
    .Q(\mem[53][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10521_ (.D(_00829_),
    .CLK(clknet_leaf_33_i_clk),
    .Q(\mem[53][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10522_ (.D(_00830_),
    .CLK(clknet_leaf_33_i_clk),
    .Q(\mem[53][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10523_ (.D(_00831_),
    .CLK(clknet_leaf_34_i_clk),
    .Q(\mem[53][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10524_ (.D(_00832_),
    .CLK(clknet_leaf_34_i_clk),
    .Q(\mem[53][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10525_ (.D(_00833_),
    .CLK(clknet_leaf_34_i_clk),
    .Q(\mem[53][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10526_ (.D(_00834_),
    .CLK(clknet_leaf_35_i_clk),
    .Q(\mem[53][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10527_ (.D(_00835_),
    .CLK(clknet_leaf_47_i_clk),
    .Q(\mem[54][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10528_ (.D(_00836_),
    .CLK(clknet_leaf_35_i_clk),
    .Q(\mem[54][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10529_ (.D(_00837_),
    .CLK(clknet_leaf_35_i_clk),
    .Q(\mem[54][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10530_ (.D(_00838_),
    .CLK(clknet_leaf_35_i_clk),
    .Q(\mem[54][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10531_ (.D(_00839_),
    .CLK(clknet_leaf_35_i_clk),
    .Q(\mem[54][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10532_ (.D(_00840_),
    .CLK(clknet_leaf_34_i_clk),
    .Q(\mem[54][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10533_ (.D(_00841_),
    .CLK(clknet_leaf_34_i_clk),
    .Q(\mem[54][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10534_ (.D(_00842_),
    .CLK(clknet_leaf_34_i_clk),
    .Q(\mem[54][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10535_ (.D(_00843_),
    .CLK(clknet_leaf_34_i_clk),
    .Q(\mem[54][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10536_ (.D(_00844_),
    .CLK(clknet_leaf_34_i_clk),
    .Q(\mem[54][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10537_ (.D(_00845_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[54][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10538_ (.D(_00846_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[54][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10539_ (.D(_00847_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[54][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10540_ (.D(_00848_),
    .CLK(clknet_leaf_34_i_clk),
    .Q(\mem[54][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10541_ (.D(_00849_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[54][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10542_ (.D(_00850_),
    .CLK(clknet_leaf_47_i_clk),
    .Q(\mem[54][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10543_ (.D(_00851_),
    .CLK(clknet_leaf_43_i_clk),
    .Q(\mem[55][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10544_ (.D(_00852_),
    .CLK(clknet_leaf_42_i_clk),
    .Q(\mem[55][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10545_ (.D(_00853_),
    .CLK(clknet_leaf_47_i_clk),
    .Q(\mem[55][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10546_ (.D(_00854_),
    .CLK(clknet_leaf_47_i_clk),
    .Q(\mem[55][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10547_ (.D(_00855_),
    .CLK(clknet_leaf_47_i_clk),
    .Q(\mem[55][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10548_ (.D(_00856_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[55][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10549_ (.D(_00857_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[55][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10550_ (.D(_00858_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[55][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10551_ (.D(_00859_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[55][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10552_ (.D(_00860_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[55][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10553_ (.D(_00861_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[55][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10554_ (.D(_00862_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[55][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10555_ (.D(_00863_),
    .CLK(clknet_leaf_47_i_clk),
    .Q(\mem[55][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10556_ (.D(_00864_),
    .CLK(clknet_leaf_48_i_clk),
    .Q(\mem[55][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10557_ (.D(_00865_),
    .CLK(clknet_leaf_47_i_clk),
    .Q(\mem[55][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10558_ (.D(_00866_),
    .CLK(clknet_leaf_46_i_clk),
    .Q(\mem[55][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10559_ (.D(_00867_),
    .CLK(clknet_leaf_38_i_clk),
    .Q(\mem[56][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10560_ (.D(_00868_),
    .CLK(clknet_leaf_22_i_clk),
    .Q(\mem[56][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10561_ (.D(_00869_),
    .CLK(clknet_leaf_23_i_clk),
    .Q(\mem[56][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10562_ (.D(_00870_),
    .CLK(clknet_leaf_22_i_clk),
    .Q(\mem[56][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10563_ (.D(_00871_),
    .CLK(clknet_leaf_25_i_clk),
    .Q(\mem[56][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10564_ (.D(_00872_),
    .CLK(clknet_leaf_25_i_clk),
    .Q(\mem[56][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10565_ (.D(_00873_),
    .CLK(clknet_leaf_25_i_clk),
    .Q(\mem[56][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10566_ (.D(_00874_),
    .CLK(clknet_leaf_24_i_clk),
    .Q(\mem[56][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10567_ (.D(_00875_),
    .CLK(clknet_leaf_25_i_clk),
    .Q(\mem[56][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10568_ (.D(_00876_),
    .CLK(clknet_leaf_24_i_clk),
    .Q(\mem[56][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10569_ (.D(_00877_),
    .CLK(clknet_leaf_30_i_clk),
    .Q(\mem[56][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10570_ (.D(_00878_),
    .CLK(clknet_leaf_30_i_clk),
    .Q(\mem[56][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10571_ (.D(_00879_),
    .CLK(clknet_leaf_30_i_clk),
    .Q(\mem[56][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10572_ (.D(_00880_),
    .CLK(clknet_leaf_38_i_clk),
    .Q(\mem[56][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10573_ (.D(_00881_),
    .CLK(clknet_leaf_37_i_clk),
    .Q(\mem[56][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10574_ (.D(_00882_),
    .CLK(clknet_leaf_37_i_clk),
    .Q(\mem[56][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10575_ (.D(_00883_),
    .CLK(clknet_leaf_37_i_clk),
    .Q(\mem[57][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10576_ (.D(_00884_),
    .CLK(clknet_leaf_23_i_clk),
    .Q(\mem[57][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10577_ (.D(_00885_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[57][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10578_ (.D(_00886_),
    .CLK(clknet_leaf_30_i_clk),
    .Q(\mem[57][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10579_ (.D(_00887_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[57][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10580_ (.D(_00888_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[57][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10581_ (.D(_00889_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[57][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10582_ (.D(_00890_),
    .CLK(clknet_leaf_28_i_clk),
    .Q(\mem[57][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10583_ (.D(_00891_),
    .CLK(clknet_leaf_28_i_clk),
    .Q(\mem[57][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10584_ (.D(_00892_),
    .CLK(clknet_leaf_28_i_clk),
    .Q(\mem[57][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10585_ (.D(_00893_),
    .CLK(clknet_leaf_28_i_clk),
    .Q(\mem[57][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10586_ (.D(_00894_),
    .CLK(clknet_leaf_31_i_clk),
    .Q(\mem[57][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10587_ (.D(_00895_),
    .CLK(clknet_leaf_31_i_clk),
    .Q(\mem[57][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10588_ (.D(_00896_),
    .CLK(clknet_leaf_31_i_clk),
    .Q(\mem[57][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10589_ (.D(_00897_),
    .CLK(clknet_leaf_31_i_clk),
    .Q(\mem[57][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10590_ (.D(_00898_),
    .CLK(clknet_leaf_37_i_clk),
    .Q(\mem[57][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10591_ (.D(_00899_),
    .CLK(clknet_leaf_37_i_clk),
    .Q(\mem[58][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10592_ (.D(_00900_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[58][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10593_ (.D(_00901_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[58][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10594_ (.D(_00902_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[58][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10595_ (.D(_00903_),
    .CLK(clknet_leaf_25_i_clk),
    .Q(\mem[58][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10596_ (.D(_00904_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[58][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10597_ (.D(_00905_),
    .CLK(clknet_leaf_27_i_clk),
    .Q(\mem[58][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10598_ (.D(_00906_),
    .CLK(clknet_leaf_27_i_clk),
    .Q(\mem[58][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10599_ (.D(_00907_),
    .CLK(clknet_leaf_27_i_clk),
    .Q(\mem[58][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10600_ (.D(_00908_),
    .CLK(clknet_leaf_24_i_clk),
    .Q(\mem[58][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10601_ (.D(_00909_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[58][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10602_ (.D(_00910_),
    .CLK(clknet_leaf_31_i_clk),
    .Q(\mem[58][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10603_ (.D(_00911_),
    .CLK(clknet_leaf_31_i_clk),
    .Q(\mem[58][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10604_ (.D(_00912_),
    .CLK(clknet_leaf_31_i_clk),
    .Q(\mem[58][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10605_ (.D(_00913_),
    .CLK(clknet_leaf_31_i_clk),
    .Q(\mem[58][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10606_ (.D(_00914_),
    .CLK(clknet_leaf_37_i_clk),
    .Q(\mem[58][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10607_ (.D(_00915_),
    .CLK(clknet_leaf_42_i_clk),
    .Q(\mem[5][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10608_ (.D(_00916_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[5][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10609_ (.D(_00917_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[5][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10610_ (.D(_00918_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[5][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10611_ (.D(_00919_),
    .CLK(clknet_leaf_36_i_clk),
    .Q(\mem[5][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10612_ (.D(_00920_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[5][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10613_ (.D(_00921_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[5][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10614_ (.D(_00922_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[5][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10615_ (.D(_00923_),
    .CLK(clknet_leaf_36_i_clk),
    .Q(\mem[5][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10616_ (.D(_00924_),
    .CLK(clknet_leaf_36_i_clk),
    .Q(\mem[5][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10617_ (.D(_00925_),
    .CLK(clknet_leaf_36_i_clk),
    .Q(\mem[5][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10618_ (.D(_00926_),
    .CLK(clknet_leaf_39_i_clk),
    .Q(\mem[5][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10619_ (.D(_00927_),
    .CLK(clknet_leaf_43_i_clk),
    .Q(\mem[5][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10620_ (.D(_00928_),
    .CLK(clknet_leaf_47_i_clk),
    .Q(\mem[5][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10621_ (.D(_00929_),
    .CLK(clknet_leaf_47_i_clk),
    .Q(\mem[5][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10622_ (.D(_00930_),
    .CLK(clknet_leaf_43_i_clk),
    .Q(\mem[5][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10623_ (.D(_00931_),
    .CLK(clknet_leaf_36_i_clk),
    .Q(\mem[60][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10624_ (.D(_00932_),
    .CLK(clknet_leaf_23_i_clk),
    .Q(\mem[60][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10625_ (.D(_00933_),
    .CLK(clknet_leaf_23_i_clk),
    .Q(\mem[60][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10626_ (.D(_00934_),
    .CLK(clknet_leaf_24_i_clk),
    .Q(\mem[60][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10627_ (.D(_00935_),
    .CLK(clknet_leaf_25_i_clk),
    .Q(\mem[60][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10628_ (.D(_00936_),
    .CLK(clknet_leaf_25_i_clk),
    .Q(\mem[60][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10629_ (.D(_00937_),
    .CLK(clknet_leaf_25_i_clk),
    .Q(\mem[60][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10630_ (.D(_00938_),
    .CLK(clknet_leaf_24_i_clk),
    .Q(\mem[60][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10631_ (.D(_00939_),
    .CLK(clknet_leaf_25_i_clk),
    .Q(\mem[60][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10632_ (.D(_00940_),
    .CLK(clknet_leaf_24_i_clk),
    .Q(\mem[60][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10633_ (.D(_00941_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[60][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10634_ (.D(_00942_),
    .CLK(clknet_leaf_30_i_clk),
    .Q(\mem[60][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10635_ (.D(_00943_),
    .CLK(clknet_leaf_30_i_clk),
    .Q(\mem[60][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10636_ (.D(_00944_),
    .CLK(clknet_leaf_30_i_clk),
    .Q(\mem[60][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10637_ (.D(_00945_),
    .CLK(clknet_leaf_36_i_clk),
    .Q(\mem[60][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10638_ (.D(_00946_),
    .CLK(clknet_leaf_36_i_clk),
    .Q(\mem[60][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10639_ (.D(_00947_),
    .CLK(clknet_leaf_33_i_clk),
    .Q(\mem[61][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10640_ (.D(_00948_),
    .CLK(clknet_leaf_27_i_clk),
    .Q(\mem[61][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10641_ (.D(_00949_),
    .CLK(clknet_leaf_28_i_clk),
    .Q(\mem[61][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10642_ (.D(_00950_),
    .CLK(clknet_leaf_27_i_clk),
    .Q(\mem[61][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10643_ (.D(_00951_),
    .CLK(clknet_leaf_25_i_clk),
    .Q(\mem[61][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10644_ (.D(_00952_),
    .CLK(clknet_leaf_26_i_clk),
    .Q(\mem[61][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10645_ (.D(_00953_),
    .CLK(clknet_leaf_26_i_clk),
    .Q(\mem[61][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10646_ (.D(_00954_),
    .CLK(clknet_leaf_27_i_clk),
    .Q(\mem[61][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10647_ (.D(_00955_),
    .CLK(clknet_leaf_26_i_clk),
    .Q(\mem[61][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10648_ (.D(_00956_),
    .CLK(clknet_leaf_28_i_clk),
    .Q(\mem[61][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10649_ (.D(_00957_),
    .CLK(clknet_leaf_28_i_clk),
    .Q(\mem[61][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10650_ (.D(_00958_),
    .CLK(clknet_leaf_32_i_clk),
    .Q(\mem[61][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10651_ (.D(_00959_),
    .CLK(clknet_leaf_32_i_clk),
    .Q(\mem[61][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10652_ (.D(_00960_),
    .CLK(clknet_leaf_32_i_clk),
    .Q(\mem[61][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10653_ (.D(_00961_),
    .CLK(clknet_leaf_32_i_clk),
    .Q(\mem[61][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10654_ (.D(_00962_),
    .CLK(clknet_leaf_32_i_clk),
    .Q(\mem[61][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10655_ (.D(_00963_),
    .CLK(clknet_leaf_33_i_clk),
    .Q(\mem[62][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10656_ (.D(_00964_),
    .CLK(clknet_leaf_27_i_clk),
    .Q(\mem[62][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10657_ (.D(_00965_),
    .CLK(clknet_leaf_27_i_clk),
    .Q(\mem[62][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10658_ (.D(_00966_),
    .CLK(clknet_leaf_29_i_clk),
    .Q(\mem[62][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10659_ (.D(_00967_),
    .CLK(clknet_leaf_26_i_clk),
    .Q(\mem[62][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10660_ (.D(_00968_),
    .CLK(clknet_leaf_26_i_clk),
    .Q(\mem[62][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10661_ (.D(_00969_),
    .CLK(clknet_leaf_26_i_clk),
    .Q(\mem[62][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10662_ (.D(_00970_),
    .CLK(clknet_leaf_27_i_clk),
    .Q(\mem[62][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10663_ (.D(_00971_),
    .CLK(clknet_leaf_26_i_clk),
    .Q(\mem[62][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10664_ (.D(_00972_),
    .CLK(clknet_leaf_27_i_clk),
    .Q(\mem[62][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10665_ (.D(_00973_),
    .CLK(clknet_leaf_28_i_clk),
    .Q(\mem[62][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10666_ (.D(_00974_),
    .CLK(clknet_leaf_32_i_clk),
    .Q(\mem[62][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10667_ (.D(_00975_),
    .CLK(clknet_leaf_32_i_clk),
    .Q(\mem[62][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10668_ (.D(_00976_),
    .CLK(clknet_leaf_32_i_clk),
    .Q(\mem[62][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10669_ (.D(_00977_),
    .CLK(clknet_leaf_32_i_clk),
    .Q(\mem[62][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10670_ (.D(_00978_),
    .CLK(clknet_leaf_33_i_clk),
    .Q(\mem[62][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10671_ (.D(_00000_),
    .CLK(clknet_leaf_85_i_clk),
    .Q(net24),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10672_ (.D(_00007_),
    .CLK(clknet_leaf_85_i_clk),
    .Q(net31),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10673_ (.D(_00008_),
    .CLK(clknet_leaf_81_i_clk),
    .Q(net32),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10674_ (.D(_00009_),
    .CLK(clknet_leaf_80_i_clk),
    .Q(net33),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10675_ (.D(_00010_),
    .CLK(clknet_leaf_79_i_clk),
    .Q(net34),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10676_ (.D(_00011_),
    .CLK(clknet_leaf_79_i_clk),
    .Q(net35),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10677_ (.D(_00012_),
    .CLK(clknet_leaf_64_i_clk),
    .Q(net36),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10678_ (.D(_00013_),
    .CLK(clknet_leaf_63_i_clk),
    .Q(net37),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10679_ (.D(_00014_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(net38),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10680_ (.D(_00015_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(net39),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10681_ (.D(_00001_),
    .CLK(clknet_leaf_62_i_clk),
    .Q(net25),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10682_ (.D(_00002_),
    .CLK(clknet_leaf_57_i_clk),
    .Q(net26),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10683_ (.D(_00003_),
    .CLK(clknet_leaf_57_i_clk),
    .Q(net27),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10684_ (.D(_00004_),
    .CLK(clknet_leaf_57_i_clk),
    .Q(net28),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10685_ (.D(_00005_),
    .CLK(clknet_leaf_56_i_clk),
    .Q(net29),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10686_ (.D(_00006_),
    .CLK(clknet_leaf_56_i_clk),
    .Q(net30),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10687_ (.D(_00979_),
    .CLK(clknet_leaf_13_i_clk),
    .Q(\mem[9][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10688_ (.D(_00980_),
    .CLK(clknet_leaf_40_i_clk),
    .Q(\mem[9][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10689_ (.D(_00981_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[9][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10690_ (.D(_00982_),
    .CLK(clknet_leaf_40_i_clk),
    .Q(\mem[9][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10691_ (.D(_00983_),
    .CLK(clknet_leaf_11_i_clk),
    .Q(\mem[9][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10692_ (.D(_00984_),
    .CLK(clknet_leaf_14_i_clk),
    .Q(\mem[9][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10693_ (.D(_00985_),
    .CLK(clknet_leaf_14_i_clk),
    .Q(\mem[9][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10694_ (.D(_00986_),
    .CLK(clknet_leaf_14_i_clk),
    .Q(\mem[9][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10695_ (.D(_00987_),
    .CLK(clknet_leaf_14_i_clk),
    .Q(\mem[9][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10696_ (.D(_00988_),
    .CLK(clknet_leaf_14_i_clk),
    .Q(\mem[9][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10697_ (.D(_00989_),
    .CLK(clknet_leaf_14_i_clk),
    .Q(\mem[9][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10698_ (.D(_00990_),
    .CLK(clknet_leaf_13_i_clk),
    .Q(\mem[9][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10699_ (.D(_00991_),
    .CLK(clknet_leaf_13_i_clk),
    .Q(\mem[9][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10700_ (.D(_00992_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[9][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10701_ (.D(_00993_),
    .CLK(clknet_leaf_15_i_clk),
    .Q(\mem[9][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10702_ (.D(_00994_),
    .CLK(clknet_leaf_14_i_clk),
    .Q(\mem[9][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10703_ (.D(_00995_),
    .CLK(clknet_leaf_42_i_clk),
    .Q(\mem[49][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10704_ (.D(net73),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[49][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10705_ (.D(_00997_),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[49][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10706_ (.D(_00998_),
    .CLK(clknet_leaf_42_i_clk),
    .Q(\mem[49][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10707_ (.D(_00999_),
    .CLK(clknet_leaf_68_i_clk),
    .Q(\mem[49][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10708_ (.D(_01000_),
    .CLK(clknet_leaf_44_i_clk),
    .Q(\mem[49][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10709_ (.D(_01001_),
    .CLK(clknet_leaf_44_i_clk),
    .Q(\mem[49][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10710_ (.D(_01002_),
    .CLK(clknet_leaf_44_i_clk),
    .Q(\mem[49][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10711_ (.D(_01003_),
    .CLK(clknet_leaf_44_i_clk),
    .Q(\mem[49][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10712_ (.D(_01004_),
    .CLK(clknet_leaf_44_i_clk),
    .Q(\mem[49][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10713_ (.D(_01005_),
    .CLK(clknet_leaf_43_i_clk),
    .Q(\mem[49][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10714_ (.D(_01006_),
    .CLK(clknet_leaf_43_i_clk),
    .Q(\mem[49][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10715_ (.D(_01007_),
    .CLK(clknet_leaf_43_i_clk),
    .Q(\mem[49][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10716_ (.D(_01008_),
    .CLK(clknet_leaf_43_i_clk),
    .Q(\mem[49][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10717_ (.D(_01009_),
    .CLK(clknet_leaf_42_i_clk),
    .Q(\mem[49][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10718_ (.D(_01010_),
    .CLK(clknet_leaf_42_i_clk),
    .Q(\mem[49][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10719_ (.D(net149),
    .CLK(clknet_leaf_91_i_clk),
    .Q(\mem[39][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10720_ (.D(net44),
    .CLK(clknet_leaf_91_i_clk),
    .Q(\mem[39][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10721_ (.D(net128),
    .CLK(clknet_leaf_84_i_clk),
    .Q(\mem[39][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10722_ (.D(net53),
    .CLK(clknet_leaf_83_i_clk),
    .Q(\mem[39][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10723_ (.D(net47),
    .CLK(clknet_leaf_86_i_clk),
    .Q(\mem[39][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10724_ (.D(net78),
    .CLK(clknet_leaf_86_i_clk),
    .Q(\mem[39][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10725_ (.D(net108),
    .CLK(clknet_leaf_85_i_clk),
    .Q(\mem[39][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10726_ (.D(net116),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[39][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10727_ (.D(_01019_),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[39][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10728_ (.D(_01020_),
    .CLK(clknet_leaf_87_i_clk),
    .Q(\mem[39][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10729_ (.D(_01021_),
    .CLK(clknet_leaf_88_i_clk),
    .Q(\mem[39][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10730_ (.D(_01022_),
    .CLK(clknet_leaf_88_i_clk),
    .Q(\mem[39][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10731_ (.D(net152),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[39][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10732_ (.D(net145),
    .CLK(clknet_leaf_89_i_clk),
    .Q(\mem[39][13] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10733_ (.D(_01025_),
    .CLK(clknet_leaf_90_i_clk),
    .Q(\mem[39][14] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10734_ (.D(net56),
    .CLK(clknet_leaf_91_i_clk),
    .Q(\mem[39][15] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10735_ (.D(_01027_),
    .CLK(clknet_leaf_71_i_clk),
    .Q(\mem[7][0] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10736_ (.D(_01028_),
    .CLK(clknet_leaf_72_i_clk),
    .Q(\mem[7][1] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10737_ (.D(_01029_),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[7][2] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10738_ (.D(_01030_),
    .CLK(clknet_leaf_72_i_clk),
    .Q(\mem[7][3] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10739_ (.D(net63),
    .CLK(clknet_leaf_71_i_clk),
    .Q(\mem[7][4] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10740_ (.D(net50),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[7][5] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10741_ (.D(net66),
    .CLK(clknet_leaf_102_i_clk),
    .Q(\mem[7][6] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10742_ (.D(_01034_),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[7][7] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10743_ (.D(_01035_),
    .CLK(clknet_leaf_71_i_clk),
    .Q(\mem[7][8] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10744_ (.D(_01036_),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[7][9] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10745_ (.D(_01037_),
    .CLK(clknet_leaf_71_i_clk),
    .Q(\mem[7][10] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10746_ (.D(_01038_),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[7][11] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10747_ (.D(_01039_),
    .CLK(clknet_leaf_70_i_clk),
    .Q(\mem[7][12] ),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_i_clk (.I(i_clk),
    .Z(clknet_0_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_i_clk (.I(clknet_0_i_clk),
    .Z(clknet_3_0_0_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_i_clk (.I(clknet_0_i_clk),
    .Z(clknet_3_1_0_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_i_clk (.I(clknet_0_i_clk),
    .Z(clknet_3_2_0_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_i_clk (.I(clknet_0_i_clk),
    .Z(clknet_3_3_0_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_i_clk (.I(clknet_0_i_clk),
    .Z(clknet_3_4_0_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_i_clk (.I(clknet_0_i_clk),
    .Z(clknet_3_5_0_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_i_clk (.I(clknet_0_i_clk),
    .Z(clknet_3_6_0_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_i_clk (.I(clknet_0_i_clk),
    .Z(clknet_3_7_0_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_0__f_i_clk (.I(clknet_3_0_0_i_clk),
    .Z(clknet_4_0__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_10__f_i_clk (.I(clknet_3_5_0_i_clk),
    .Z(clknet_4_10__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_11__f_i_clk (.I(clknet_3_5_0_i_clk),
    .Z(clknet_4_11__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_12__f_i_clk (.I(clknet_3_6_0_i_clk),
    .Z(clknet_4_12__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_13__f_i_clk (.I(clknet_3_6_0_i_clk),
    .Z(clknet_4_13__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_14__f_i_clk (.I(clknet_3_7_0_i_clk),
    .Z(clknet_4_14__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_15__f_i_clk (.I(clknet_3_7_0_i_clk),
    .Z(clknet_4_15__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_1__f_i_clk (.I(clknet_3_0_0_i_clk),
    .Z(clknet_4_1__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_2__f_i_clk (.I(clknet_3_1_0_i_clk),
    .Z(clknet_4_2__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_3__f_i_clk (.I(clknet_3_1_0_i_clk),
    .Z(clknet_4_3__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_4__f_i_clk (.I(clknet_3_2_0_i_clk),
    .Z(clknet_4_4__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_5__f_i_clk (.I(clknet_3_2_0_i_clk),
    .Z(clknet_4_5__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_6__f_i_clk (.I(clknet_3_3_0_i_clk),
    .Z(clknet_4_6__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_7__f_i_clk (.I(clknet_3_3_0_i_clk),
    .Z(clknet_4_7__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_8__f_i_clk (.I(clknet_3_4_0_i_clk),
    .Z(clknet_4_8__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_9__f_i_clk (.I(clknet_3_4_0_i_clk),
    .Z(clknet_4_9__leaf_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_i_clk (.I(clknet_4_0__leaf_i_clk),
    .Z(clknet_leaf_0_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_i_clk (.I(clknet_4_9__leaf_i_clk),
    .Z(clknet_leaf_100_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_i_clk (.I(clknet_4_9__leaf_i_clk),
    .Z(clknet_leaf_101_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_i_clk (.I(clknet_4_9__leaf_i_clk),
    .Z(clknet_leaf_102_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_i_clk (.I(clknet_4_3__leaf_i_clk),
    .Z(clknet_leaf_103_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_i_clk (.I(clknet_4_3__leaf_i_clk),
    .Z(clknet_leaf_104_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_i_clk (.I(clknet_4_3__leaf_i_clk),
    .Z(clknet_leaf_105_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_i_clk (.I(clknet_4_2__leaf_i_clk),
    .Z(clknet_leaf_106_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_i_clk (.I(clknet_4_2__leaf_i_clk),
    .Z(clknet_leaf_107_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_i_clk (.I(clknet_4_2__leaf_i_clk),
    .Z(clknet_leaf_108_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_i_clk (.I(clknet_4_2__leaf_i_clk),
    .Z(clknet_leaf_109_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_i_clk (.I(clknet_4_3__leaf_i_clk),
    .Z(clknet_leaf_10_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_i_clk (.I(clknet_4_2__leaf_i_clk),
    .Z(clknet_leaf_110_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_i_clk (.I(clknet_4_2__leaf_i_clk),
    .Z(clknet_leaf_111_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_i_clk (.I(clknet_4_2__leaf_i_clk),
    .Z(clknet_leaf_112_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_i_clk (.I(clknet_4_0__leaf_i_clk),
    .Z(clknet_leaf_113_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_i_clk (.I(clknet_4_0__leaf_i_clk),
    .Z(clknet_leaf_114_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_i_clk (.I(clknet_4_0__leaf_i_clk),
    .Z(clknet_leaf_115_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_i_clk (.I(clknet_4_0__leaf_i_clk),
    .Z(clknet_leaf_116_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_i_clk (.I(clknet_4_0__leaf_i_clk),
    .Z(clknet_leaf_117_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_i_clk (.I(clknet_4_0__leaf_i_clk),
    .Z(clknet_leaf_118_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_i_clk (.I(clknet_4_3__leaf_i_clk),
    .Z(clknet_leaf_11_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_i_clk (.I(clknet_4_3__leaf_i_clk),
    .Z(clknet_leaf_12_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_i_clk (.I(clknet_4_6__leaf_i_clk),
    .Z(clknet_leaf_13_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_i_clk (.I(clknet_4_6__leaf_i_clk),
    .Z(clknet_leaf_14_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_i_clk (.I(clknet_4_6__leaf_i_clk),
    .Z(clknet_leaf_15_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_i_clk (.I(clknet_4_4__leaf_i_clk),
    .Z(clknet_leaf_16_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_i_clk (.I(clknet_4_4__leaf_i_clk),
    .Z(clknet_leaf_17_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_i_clk (.I(clknet_4_4__leaf_i_clk),
    .Z(clknet_leaf_18_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_i_clk (.I(clknet_4_4__leaf_i_clk),
    .Z(clknet_leaf_19_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_i_clk (.I(clknet_4_1__leaf_i_clk),
    .Z(clknet_leaf_1_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_i_clk (.I(clknet_4_4__leaf_i_clk),
    .Z(clknet_leaf_20_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_i_clk (.I(clknet_4_4__leaf_i_clk),
    .Z(clknet_leaf_21_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_i_clk (.I(clknet_4_4__leaf_i_clk),
    .Z(clknet_leaf_22_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_i_clk (.I(clknet_4_5__leaf_i_clk),
    .Z(clknet_leaf_23_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_i_clk (.I(clknet_4_5__leaf_i_clk),
    .Z(clknet_leaf_24_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_i_clk (.I(clknet_4_5__leaf_i_clk),
    .Z(clknet_leaf_25_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_i_clk (.I(clknet_4_5__leaf_i_clk),
    .Z(clknet_leaf_26_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_i_clk (.I(clknet_4_5__leaf_i_clk),
    .Z(clknet_leaf_27_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_i_clk (.I(clknet_4_5__leaf_i_clk),
    .Z(clknet_leaf_28_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_i_clk (.I(clknet_4_5__leaf_i_clk),
    .Z(clknet_leaf_29_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_i_clk (.I(clknet_4_1__leaf_i_clk),
    .Z(clknet_leaf_2_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_i_clk (.I(clknet_4_7__leaf_i_clk),
    .Z(clknet_leaf_30_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_i_clk (.I(clknet_4_7__leaf_i_clk),
    .Z(clknet_leaf_31_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_i_clk (.I(clknet_4_7__leaf_i_clk),
    .Z(clknet_leaf_32_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_i_clk (.I(clknet_4_7__leaf_i_clk),
    .Z(clknet_leaf_33_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_i_clk (.I(clknet_4_7__leaf_i_clk),
    .Z(clknet_leaf_34_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_i_clk (.I(clknet_4_7__leaf_i_clk),
    .Z(clknet_leaf_35_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_i_clk (.I(clknet_4_7__leaf_i_clk),
    .Z(clknet_leaf_36_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_i_clk (.I(clknet_4_7__leaf_i_clk),
    .Z(clknet_leaf_37_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_i_clk (.I(clknet_4_6__leaf_i_clk),
    .Z(clknet_leaf_38_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_i_clk (.I(clknet_4_6__leaf_i_clk),
    .Z(clknet_leaf_39_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_i_clk (.I(clknet_4_1__leaf_i_clk),
    .Z(clknet_leaf_3_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_i_clk (.I(clknet_4_6__leaf_i_clk),
    .Z(clknet_leaf_40_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_i_clk (.I(clknet_4_12__leaf_i_clk),
    .Z(clknet_leaf_41_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_i_clk (.I(clknet_4_12__leaf_i_clk),
    .Z(clknet_leaf_42_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_i_clk (.I(clknet_4_12__leaf_i_clk),
    .Z(clknet_leaf_43_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_i_clk (.I(clknet_4_12__leaf_i_clk),
    .Z(clknet_leaf_44_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_i_clk (.I(clknet_4_13__leaf_i_clk),
    .Z(clknet_leaf_45_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_i_clk (.I(clknet_4_13__leaf_i_clk),
    .Z(clknet_leaf_46_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_i_clk (.I(clknet_4_13__leaf_i_clk),
    .Z(clknet_leaf_47_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_i_clk (.I(clknet_4_13__leaf_i_clk),
    .Z(clknet_leaf_48_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_i_clk (.I(clknet_4_13__leaf_i_clk),
    .Z(clknet_leaf_49_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_i_clk (.I(clknet_4_1__leaf_i_clk),
    .Z(clknet_leaf_4_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_i_clk (.I(clknet_4_13__leaf_i_clk),
    .Z(clknet_leaf_50_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_i_clk (.I(clknet_4_13__leaf_i_clk),
    .Z(clknet_leaf_51_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_i_clk (.I(clknet_4_15__leaf_i_clk),
    .Z(clknet_leaf_52_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_i_clk (.I(clknet_4_15__leaf_i_clk),
    .Z(clknet_leaf_53_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_i_clk (.I(clknet_4_15__leaf_i_clk),
    .Z(clknet_leaf_54_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_i_clk (.I(clknet_4_15__leaf_i_clk),
    .Z(clknet_leaf_55_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_i_clk (.I(clknet_4_15__leaf_i_clk),
    .Z(clknet_leaf_56_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_i_clk (.I(clknet_4_15__leaf_i_clk),
    .Z(clknet_leaf_57_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_i_clk (.I(clknet_4_15__leaf_i_clk),
    .Z(clknet_leaf_58_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_i_clk (.I(clknet_4_15__leaf_i_clk),
    .Z(clknet_leaf_59_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_i_clk (.I(clknet_4_1__leaf_i_clk),
    .Z(clknet_leaf_5_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_i_clk (.I(clknet_4_14__leaf_i_clk),
    .Z(clknet_leaf_60_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_i_clk (.I(clknet_4_14__leaf_i_clk),
    .Z(clknet_leaf_61_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_i_clk (.I(clknet_4_14__leaf_i_clk),
    .Z(clknet_leaf_62_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_i_clk (.I(clknet_4_14__leaf_i_clk),
    .Z(clknet_leaf_63_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_i_clk (.I(clknet_4_14__leaf_i_clk),
    .Z(clknet_leaf_64_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_i_clk (.I(clknet_4_14__leaf_i_clk),
    .Z(clknet_leaf_65_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_i_clk (.I(clknet_4_14__leaf_i_clk),
    .Z(clknet_leaf_66_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_i_clk (.I(clknet_4_14__leaf_i_clk),
    .Z(clknet_leaf_67_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_i_clk (.I(clknet_4_12__leaf_i_clk),
    .Z(clknet_leaf_68_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_i_clk (.I(clknet_4_12__leaf_i_clk),
    .Z(clknet_leaf_69_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_i_clk (.I(clknet_4_1__leaf_i_clk),
    .Z(clknet_leaf_6_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_i_clk (.I(clknet_4_12__leaf_i_clk),
    .Z(clknet_leaf_70_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_i_clk (.I(clknet_4_9__leaf_i_clk),
    .Z(clknet_leaf_71_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_i_clk (.I(clknet_4_9__leaf_i_clk),
    .Z(clknet_leaf_72_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_i_clk (.I(clknet_4_9__leaf_i_clk),
    .Z(clknet_leaf_73_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_i_clk (.I(clknet_4_9__leaf_i_clk),
    .Z(clknet_leaf_74_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_i_clk (.I(clknet_4_11__leaf_i_clk),
    .Z(clknet_leaf_75_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_i_clk (.I(clknet_4_11__leaf_i_clk),
    .Z(clknet_leaf_76_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_i_clk (.I(clknet_4_11__leaf_i_clk),
    .Z(clknet_leaf_77_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_i_clk (.I(clknet_4_11__leaf_i_clk),
    .Z(clknet_leaf_78_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_i_clk (.I(clknet_4_11__leaf_i_clk),
    .Z(clknet_leaf_79_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_i_clk (.I(clknet_4_1__leaf_i_clk),
    .Z(clknet_leaf_7_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_i_clk (.I(clknet_4_11__leaf_i_clk),
    .Z(clknet_leaf_80_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_i_clk (.I(clknet_4_11__leaf_i_clk),
    .Z(clknet_leaf_81_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_i_clk (.I(clknet_4_11__leaf_i_clk),
    .Z(clknet_leaf_82_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_i_clk (.I(clknet_4_10__leaf_i_clk),
    .Z(clknet_leaf_83_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_i_clk (.I(clknet_4_10__leaf_i_clk),
    .Z(clknet_leaf_84_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_i_clk (.I(clknet_4_10__leaf_i_clk),
    .Z(clknet_leaf_85_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_i_clk (.I(clknet_4_10__leaf_i_clk),
    .Z(clknet_leaf_86_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_i_clk (.I(clknet_4_10__leaf_i_clk),
    .Z(clknet_leaf_87_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_i_clk (.I(clknet_4_10__leaf_i_clk),
    .Z(clknet_leaf_88_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_i_clk (.I(clknet_4_10__leaf_i_clk),
    .Z(clknet_leaf_89_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_i_clk (.I(clknet_4_1__leaf_i_clk),
    .Z(clknet_leaf_8_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_i_clk (.I(clknet_4_10__leaf_i_clk),
    .Z(clknet_leaf_90_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_i_clk (.I(clknet_4_8__leaf_i_clk),
    .Z(clknet_leaf_91_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_i_clk (.I(clknet_4_8__leaf_i_clk),
    .Z(clknet_leaf_92_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_i_clk (.I(clknet_4_8__leaf_i_clk),
    .Z(clknet_leaf_93_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_i_clk (.I(clknet_4_8__leaf_i_clk),
    .Z(clknet_leaf_94_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_i_clk (.I(clknet_4_8__leaf_i_clk),
    .Z(clknet_leaf_95_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_i_clk (.I(clknet_4_8__leaf_i_clk),
    .Z(clknet_leaf_96_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_i_clk (.I(clknet_4_8__leaf_i_clk),
    .Z(clknet_leaf_97_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_i_clk (.I(clknet_4_8__leaf_i_clk),
    .Z(clknet_leaf_98_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_i_clk (.I(clknet_4_9__leaf_i_clk),
    .Z(clknet_leaf_99_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_i_clk (.I(clknet_4_3__leaf_i_clk),
    .Z(clknet_leaf_9_i_clk),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold1 (.I(net162),
    .Z(net42),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold10 (.I(net140),
    .Z(net51),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold100 (.I(net51),
    .Z(net141),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold101 (.I(_01078_),
    .Z(net142),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold102 (.I(i_data[13]),
    .Z(net143),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold103 (.I(net99),
    .Z(net144),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold104 (.I(_01024_),
    .Z(net145),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold105 (.I(i_addr[3]),
    .Z(net146),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold106 (.I(i_data[0]),
    .Z(net147),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold107 (.I(net81),
    .Z(net148),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold108 (.I(_01011_),
    .Z(net149),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold109 (.I(i_data[12]),
    .Z(net150),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold11 (.I(net16),
    .Z(net52),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold110 (.I(net101),
    .Z(net151),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold111 (.I(_01023_),
    .Z(net152),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold112 (.I(i_addr[4]),
    .Z(net153),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold113 (.I(i_data[11]),
    .Z(net154),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold114 (.I(net103),
    .Z(net155),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold115 (.I(i_data[15]),
    .Z(net156),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold116 (.I(net54),
    .Z(net157),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold117 (.I(i_data[8]),
    .Z(net158),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold118 (.I(net105),
    .Z(net159),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold119 (.I(i_data[10]),
    .Z(net160),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold12 (.I(_01014_),
    .Z(net53),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold120 (.I(net111),
    .Z(net161),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold121 (.I(i_data[1]),
    .Z(net162),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold122 (.I(net42),
    .Z(net163),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold123 (.I(i_we),
    .Z(net164),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold124 (.I(i_data[14]),
    .Z(net165),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold125 (.I(net83),
    .Z(net166),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold126 (.I(i_addr[1]),
    .Z(net167),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold127 (.I(i_data[9]),
    .Z(net168),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold128 (.I(net113),
    .Z(net169),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold129 (.I(_01154_),
    .Z(net170),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold13 (.I(net156),
    .Z(net54),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold14 (.I(net13),
    .Z(net55),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold15 (.I(_01026_),
    .Z(net56),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold16 (.I(net125),
    .Z(net57),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 hold17 (.I(net2),
    .Z(net58),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 hold18 (.I(_01074_),
    .Z(net59),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 hold19 (.I(_03441_),
    .Z(net60),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold2 (.I(net14),
    .Z(net43),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 hold20 (.I(_03442_),
    .Z(net61),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 hold21 (.I(_03443_),
    .Z(net62),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(_01031_),
    .Z(net63),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(net75),
    .Z(net64),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold24 (.I(net19),
    .Z(net65),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(_01033_),
    .Z(net66),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(net153),
    .Z(net67),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 hold27 (.I(net5),
    .Z(net68),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold28 (.I(_01217_),
    .Z(net69),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 hold29 (.I(_01329_),
    .Z(net70),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold3 (.I(_01012_),
    .Z(net44),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 hold30 (.I(_04800_),
    .Z(net71),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 hold31 (.I(_04801_),
    .Z(net72),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(_00996_),
    .Z(net73),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold33 (.I(net146),
    .Z(net74),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold34 (.I(i_data[6]),
    .Z(net75),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 hold35 (.I(_01126_),
    .Z(net76),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold36 (.I(_04820_),
    .Z(net77),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(_01016_),
    .Z(net78),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(net117),
    .Z(net79),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold39 (.I(net15),
    .Z(net80),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold4 (.I(net135),
    .Z(net45),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(net147),
    .Z(net81),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold41 (.I(net7),
    .Z(net82),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(net165),
    .Z(net83),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold43 (.I(net12),
    .Z(net84),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(net133),
    .Z(net85),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold45 (.I(net6),
    .Z(net86),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 hold46 (.I(_01233_),
    .Z(net87),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 hold47 (.I(_03454_),
    .Z(net88),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold48 (.I(_04760_),
    .Z(net89),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(net123),
    .Z(net90),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold5 (.I(net17),
    .Z(net46),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 hold50 (.I(net23),
    .Z(net91),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold51 (.I(_03789_),
    .Z(net92),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 hold52 (.I(_03790_),
    .Z(net93),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(net109),
    .Z(net94),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold54 (.I(net20),
    .Z(net95),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold55 (.I(i_addr[0]),
    .Z(net96),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 hold56 (.I(net1),
    .Z(net97),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 hold57 (.I(_01160_),
    .Z(net98),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(net143),
    .Z(net99),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold59 (.I(net11),
    .Z(net100),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold6 (.I(_01015_),
    .Z(net47),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(net150),
    .Z(net101),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold61 (.I(net10),
    .Z(net102),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(net154),
    .Z(net103),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold63 (.I(net9),
    .Z(net104),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(net158),
    .Z(net105),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold65 (.I(net21),
    .Z(net106),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold66 (.I(net64),
    .Z(net107),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold67 (.I(_01017_),
    .Z(net108),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold68 (.I(i_data[7]),
    .Z(net109),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold69 (.I(_01198_),
    .Z(net110),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold7 (.I(net129),
    .Z(net48),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(net160),
    .Z(net111),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold71 (.I(net8),
    .Z(net112),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(net168),
    .Z(net113),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold73 (.I(net22),
    .Z(net114),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold74 (.I(net94),
    .Z(net115),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold75 (.I(_01018_),
    .Z(net116),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold76 (.I(i_data[2]),
    .Z(net117),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(_01102_),
    .Z(net118),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 hold78 (.I(_03564_),
    .Z(net119),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold79 (.I(net138),
    .Z(net120),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold8 (.I(net18),
    .Z(net49),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold80 (.I(net79),
    .Z(net121),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold81 (.I(_01056_),
    .Z(net122),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(net164),
    .Z(net123),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold83 (.I(_03521_),
    .Z(net124),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(net167),
    .Z(net125),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(_01048_),
    .Z(net126),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold86 (.I(_03587_),
    .Z(net127),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold87 (.I(_01013_),
    .Z(net128),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold88 (.I(i_data[5]),
    .Z(net129),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold89 (.I(net48),
    .Z(net130),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold9 (.I(_01032_),
    .Z(net50),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold90 (.I(net97),
    .Z(net131),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 hold91 (.I(net170),
    .Z(net132),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold92 (.I(i_addr[5]),
    .Z(net133),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold93 (.I(_01178_),
    .Z(net134),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold94 (.I(i_data[4]),
    .Z(net135),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 hold95 (.I(net68),
    .Z(net136),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold96 (.I(_01080_),
    .Z(net137),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold97 (.I(i_addr[2]),
    .Z(net138),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold98 (.I(net45),
    .Z(net139),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold99 (.I(i_data[3]),
    .Z(net140),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1 (.I(net96),
    .Z(net1),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(net151),
    .Z(net10),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(net144),
    .Z(net11),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(net166),
    .Z(net12),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(net157),
    .Z(net13),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(net163),
    .Z(net14),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(net121),
    .Z(net15),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(net141),
    .Z(net16),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(net139),
    .Z(net17),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(net130),
    .Z(net18),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(net107),
    .Z(net19),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input2 (.I(net57),
    .Z(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(net115),
    .Z(net20),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(net159),
    .Z(net21),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(net169),
    .Z(net22),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input23 (.I(net90),
    .Z(net23),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input3 (.I(net120),
    .Z(net3),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input4 (.I(net74),
    .Z(net4),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input5 (.I(net67),
    .Z(net5),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(net85),
    .Z(net6),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(net148),
    .Z(net7),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(net161),
    .Z(net8),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(net155),
    .Z(net9),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 load_slew41 (.I(net132),
    .Z(net41),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap40 (.I(net60),
    .Z(net40),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output24 (.I(net24),
    .Z(o_data[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output25 (.I(net25),
    .Z(o_data[10]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output26 (.I(net26),
    .Z(o_data[11]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output27 (.I(net27),
    .Z(o_data[12]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output28 (.I(net28),
    .Z(o_data[13]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output29 (.I(net29),
    .Z(o_data[14]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output30 (.I(net30),
    .Z(o_data[15]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output31 (.I(net31),
    .Z(o_data[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output32 (.I(net32),
    .Z(o_data[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output33 (.I(net33),
    .Z(o_data[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output34 (.I(net34),
    .Z(o_data[4]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output35 (.I(net35),
    .Z(o_data[5]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output36 (.I(net36),
    .Z(o_data[6]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output37 (.I(net37),
    .Z(o_data[7]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output38 (.I(net38),
    .Z(o_data[8]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 output39 (.I(net39),
    .Z(o_data[9]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
endmodule
