* NGSPICE file created from interconnect_outer.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

.subckt interconnect_outer c0_clk c1_clk dcache_clk ic0_clk ic1_clk inner_clock inner_disable
+ inner_embed_mode inner_ext_irq inner_reset inner_wb_4_burst inner_wb_8_burst inner_wb_ack
+ inner_wb_adr[0] inner_wb_adr[10] inner_wb_adr[11] inner_wb_adr[12] inner_wb_adr[13]
+ inner_wb_adr[14] inner_wb_adr[15] inner_wb_adr[16] inner_wb_adr[17] inner_wb_adr[18]
+ inner_wb_adr[19] inner_wb_adr[1] inner_wb_adr[20] inner_wb_adr[21] inner_wb_adr[22]
+ inner_wb_adr[23] inner_wb_adr[2] inner_wb_adr[3] inner_wb_adr[4] inner_wb_adr[5]
+ inner_wb_adr[6] inner_wb_adr[7] inner_wb_adr[8] inner_wb_adr[9] inner_wb_cyc inner_wb_err
+ inner_wb_i_dat[0] inner_wb_i_dat[10] inner_wb_i_dat[11] inner_wb_i_dat[12] inner_wb_i_dat[13]
+ inner_wb_i_dat[14] inner_wb_i_dat[15] inner_wb_i_dat[1] inner_wb_i_dat[2] inner_wb_i_dat[3]
+ inner_wb_i_dat[4] inner_wb_i_dat[5] inner_wb_i_dat[6] inner_wb_i_dat[7] inner_wb_i_dat[8]
+ inner_wb_i_dat[9] inner_wb_o_dat[0] inner_wb_o_dat[10] inner_wb_o_dat[11] inner_wb_o_dat[12]
+ inner_wb_o_dat[13] inner_wb_o_dat[14] inner_wb_o_dat[15] inner_wb_o_dat[1] inner_wb_o_dat[2]
+ inner_wb_o_dat[3] inner_wb_o_dat[4] inner_wb_o_dat[5] inner_wb_o_dat[6] inner_wb_o_dat[7]
+ inner_wb_o_dat[8] inner_wb_o_dat[9] inner_wb_sel[0] inner_wb_sel[1] inner_wb_stb
+ inner_wb_we iram_addr[0] iram_addr[1] iram_addr[2] iram_addr[3] iram_addr[4] iram_addr[5]
+ iram_clk iram_i_data[0] iram_i_data[10] iram_i_data[11] iram_i_data[12] iram_i_data[13]
+ iram_i_data[14] iram_i_data[15] iram_i_data[1] iram_i_data[2] iram_i_data[3] iram_i_data[4]
+ iram_i_data[5] iram_i_data[6] iram_i_data[7] iram_i_data[8] iram_i_data[9] iram_o_data[0]
+ iram_o_data[10] iram_o_data[11] iram_o_data[12] iram_o_data[13] iram_o_data[14]
+ iram_o_data[15] iram_o_data[1] iram_o_data[2] iram_o_data[3] iram_o_data[4] iram_o_data[5]
+ iram_o_data[6] iram_o_data[7] iram_o_data[8] iram_o_data[9] iram_we la_data_in[0]
+ la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[11] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[22] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] m_io_in[0] m_io_in[10] m_io_in[11] m_io_in[12] m_io_in[13]
+ m_io_in[14] m_io_in[15] m_io_in[16] m_io_in[17] m_io_in[18] m_io_in[19] m_io_in[1]
+ m_io_in[20] m_io_in[21] m_io_in[22] m_io_in[23] m_io_in[24] m_io_in[25] m_io_in[26]
+ m_io_in[27] m_io_in[28] m_io_in[29] m_io_in[2] m_io_in[30] m_io_in[31] m_io_in[32]
+ m_io_in[33] m_io_in[34] m_io_in[35] m_io_in[36] m_io_in[37] m_io_in[3] m_io_in[4]
+ m_io_in[5] m_io_in[6] m_io_in[7] m_io_in[8] m_io_in[9] m_io_oeb[0] m_io_oeb[10]
+ m_io_oeb[11] m_io_oeb[12] m_io_oeb[13] m_io_oeb[14] m_io_oeb[15] m_io_oeb[16] m_io_oeb[17]
+ m_io_oeb[18] m_io_oeb[19] m_io_oeb[1] m_io_oeb[20] m_io_oeb[21] m_io_oeb[22] m_io_oeb[23]
+ m_io_oeb[24] m_io_oeb[25] m_io_oeb[26] m_io_oeb[28] m_io_oeb[29] m_io_oeb[2] m_io_oeb[30]
+ m_io_oeb[31] m_io_oeb[32] m_io_oeb[33] m_io_oeb[34] m_io_oeb[35] m_io_oeb[36] m_io_oeb[37]
+ m_io_oeb[3] m_io_oeb[4] m_io_oeb[5] m_io_oeb[6] m_io_oeb[7] m_io_oeb[8] m_io_oeb[9]
+ m_io_out[0] m_io_out[10] m_io_out[11] m_io_out[12] m_io_out[13] m_io_out[14] m_io_out[15]
+ m_io_out[16] m_io_out[17] m_io_out[18] m_io_out[19] m_io_out[1] m_io_out[20] m_io_out[21]
+ m_io_out[22] m_io_out[23] m_io_out[24] m_io_out[25] m_io_out[26] m_io_out[27] m_io_out[28]
+ m_io_out[29] m_io_out[2] m_io_out[36] m_io_out[37] m_io_out[3] m_io_out[4] m_io_out[5]
+ m_io_out[6] m_io_out[7] m_io_out[8] m_io_out[9] mgt_wb_ack_o mgt_wb_adr_i[0] mgt_wb_adr_i[10]
+ mgt_wb_adr_i[11] mgt_wb_adr_i[12] mgt_wb_adr_i[13] mgt_wb_adr_i[14] mgt_wb_adr_i[15]
+ mgt_wb_adr_i[16] mgt_wb_adr_i[17] mgt_wb_adr_i[18] mgt_wb_adr_i[19] mgt_wb_adr_i[1]
+ mgt_wb_adr_i[20] mgt_wb_adr_i[21] mgt_wb_adr_i[22] mgt_wb_adr_i[23] mgt_wb_adr_i[24]
+ mgt_wb_adr_i[25] mgt_wb_adr_i[26] mgt_wb_adr_i[27] mgt_wb_adr_i[28] mgt_wb_adr_i[29]
+ mgt_wb_adr_i[2] mgt_wb_adr_i[30] mgt_wb_adr_i[31] mgt_wb_adr_i[3] mgt_wb_adr_i[4]
+ mgt_wb_adr_i[5] mgt_wb_adr_i[6] mgt_wb_adr_i[7] mgt_wb_adr_i[8] mgt_wb_adr_i[9]
+ mgt_wb_clk_i mgt_wb_cyc_i mgt_wb_dat_i[0] mgt_wb_dat_i[10] mgt_wb_dat_i[11] mgt_wb_dat_i[12]
+ mgt_wb_dat_i[13] mgt_wb_dat_i[14] mgt_wb_dat_i[15] mgt_wb_dat_i[16] mgt_wb_dat_i[17]
+ mgt_wb_dat_i[18] mgt_wb_dat_i[19] mgt_wb_dat_i[1] mgt_wb_dat_i[20] mgt_wb_dat_i[21]
+ mgt_wb_dat_i[22] mgt_wb_dat_i[23] mgt_wb_dat_i[24] mgt_wb_dat_i[25] mgt_wb_dat_i[26]
+ mgt_wb_dat_i[27] mgt_wb_dat_i[28] mgt_wb_dat_i[29] mgt_wb_dat_i[2] mgt_wb_dat_i[30]
+ mgt_wb_dat_i[31] mgt_wb_dat_i[3] mgt_wb_dat_i[4] mgt_wb_dat_i[5] mgt_wb_dat_i[6]
+ mgt_wb_dat_i[7] mgt_wb_dat_i[8] mgt_wb_dat_i[9] mgt_wb_dat_o[0] mgt_wb_dat_o[10]
+ mgt_wb_dat_o[11] mgt_wb_dat_o[12] mgt_wb_dat_o[13] mgt_wb_dat_o[14] mgt_wb_dat_o[1]
+ mgt_wb_dat_o[20] mgt_wb_dat_o[21] mgt_wb_dat_o[22] mgt_wb_dat_o[23] mgt_wb_dat_o[24]
+ mgt_wb_dat_o[25] mgt_wb_dat_o[26] mgt_wb_dat_o[27] mgt_wb_dat_o[28] mgt_wb_dat_o[29]
+ mgt_wb_dat_o[2] mgt_wb_dat_o[30] mgt_wb_dat_o[31] mgt_wb_dat_o[6] mgt_wb_dat_o[7]
+ mgt_wb_dat_o[8] mgt_wb_dat_o[9] mgt_wb_rst_i mgt_wb_sel_i[0] mgt_wb_sel_i[1] mgt_wb_sel_i[2]
+ mgt_wb_sel_i[3] mgt_wb_stb_i mgt_wb_we_i user_clock2 vccd1 vssd1 la_data_out[39]
+ la_data_out[38] la_data_out[59] la_data_out[58] la_data_out[57] la_data_out[56]
+ m_io_out[35] la_data_out[55] m_io_out[34] mgt_wb_dat_o[19] mgt_wb_dat_o[18] m_io_out[33]
+ m_io_out[32] mgt_wb_dat_o[17] m_io_out[31] mgt_wb_dat_o[5] mgt_wb_dat_o[16] mgt_wb_dat_o[4]
+ mgt_wb_dat_o[15] m_io_out[30] mgt_wb_dat_o[3] m_io_oeb[27] irq[2] la_data_out[10]
+ la_data_out[21] irq[1] la_data_out[9] la_data_out[20] irq[0] la_data_out[8] la_data_out[29]
+ la_data_out[7] la_data_out[6] la_data_out[28] la_data_out[5] la_data_out[27] la_data_out[4]
+ la_data_out[15] la_data_out[26] la_data_out[3] la_data_out[14] la_data_out[25] la_data_out[13]
+ la_data_out[24] la_data_out[2] la_data_out[12] la_data_out[23]
X_3155_ m_arbiter.wb0_adr\[9\] sspi.req_addr\[9\] _1478_ _1483_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2106_ iram_wb_ack net53 _0733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3086_ _1431_ _1432_ _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2037_ wb_compressor.wb_i_dat\[6\] wb_cross_clk.s_m_sync.s_data_ff\[8\] _0688_ _0689_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3050__S _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2939_ _1331_ _1333_ _1334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1757__A2 _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input73_I m_io_in[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_20_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2706__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3198__A1 net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1748__A2 _0448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2812__B _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1920__A2 net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3122__B2 sspi.res_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1684__A1 _0391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3773_ net249 net160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2724_ wb_cross_clk.m_s_sync.d_data\[34\] _1080_ _0555_ _1162_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_42_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2655_ _0553_ _1102_ _0238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1606_ _1527_ m_arbiter.wb0_o_dat\[6\] _1530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_2_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2586_ wb_compressor.wb_i_dat\[10\] net78 net213 _1050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1852__I net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3207_ net186 _1509_ _1511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1675__A1 net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3138_ m_arbiter.wb0_adr\[1\] sspi.req_addr\[1\] _1400_ _1474_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3779__I net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_50_user_clock2 clknet_2_0__leaf_user_clock2 clknet_leaf_50_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3069_ clk_div.cnt\[0\] clk_div.cnt\[1\] clk_div.cnt\[2\] _1422_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2927__A1 _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2079__B _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1711__B _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2091__A1 iram_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2034__S _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2440_ wb_cross_clk.m_s_sync.s_data_ff\[26\] _0937_ _0958_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2371_ _0437_ _0889_ _0918_ _0917_ _0138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1672__I _1588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_30_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2909__A1 _0609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2385__A2 _0926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2707_ wb_cross_clk.m_s_sync.d_data\[32\] _1080_ _0555_ _1147_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2638_ net141 _1086_ _1079_ _0929_ _1087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2569_ _1041_ _0213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input36_I inner_wb_o_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1648__A1 _1563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3320__CLK clknet_4_11_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1671__I1 net14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2376__A2 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3470__CLK clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2128__A2 _0525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1887__A1 _0569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_18_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_18_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2300__A2 _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1940_ _0617_ _0618_ _0620_ _0621_ _0623_ _0002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1811__B2 _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1871_ _0553_ _0557_ _0011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1662__I1 net15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3610_ _0375_ clknet_leaf_27_user_clock2 net169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2367__A2 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3541_ _0306_ clknet_leaf_9_user_clock2 sspi.req_addr\[16\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3472_ _0010_ clknet_4_2_0_net196 wb_compressor.state\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2423_ net211 _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__2498__I _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3167__I1 sspi.req_addr\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2354_ _0907_ _0908_ _0895_ _0131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2285_ wb_cross_clk.m_s_sync.d_data\[38\] _0771_ _0861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3343__CLK clknet_4_8_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1802__A1 _0492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2182__B _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1653__I1 net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2358__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output142_I net142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2357__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1688__S _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2092__B _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1644__I1 net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2349__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_10_0_net196 clknet_0_net196 clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2070_ _0707_ _0708_ _0631_ _0047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2267__B _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Left_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2972_ _0619_ _1298_ _1351_ _1360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_8_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1923_ sspi.bit_cnt\[2\] _0607_ sspi.bit_cnt\[3\] _0608_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1854_ _0543_ _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1785_ net173 net227 net223 net200 _0482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2730__B _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3524_ _0289_ clknet_leaf_12_user_clock2 sspi.req_data\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3455_ _0235_ clknet_4_3_0_net196 net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2406_ _1539_ _0934_ _0940_ _0151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_4_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_1_user_clock2_I clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3386_ _0166_ clknet_leaf_39_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[24\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2337_ wb_cross_clk.m_wb_i_dat\[0\] _0896_ _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2268_ wb_cross_clk.m_s_sync.d_data\[33\] _0835_ _0849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2199_ _0799_ net415 _0794_ _0083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2751__A2 _0590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold30 _0791_ net417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold41 wb_cross_clk.m_s_sync.s_data_ff\[10\] net428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3190__C _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold74 _0868_ net461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold52 _0855_ net439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold63 wb_cross_clk.m_s_sync.s_data_ff\[13\] net450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold85 wb_cross_clk.m_s_sync.s_data_ff\[29\] net472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold96 net517 net483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2815__B _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2114__S1 clk_div.curr_div\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1778__B1 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3138__S _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2742__A2 _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1881__S _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3240_ net530 clknet_leaf_13_user_clock2 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2776__I _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1680__I net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3171_ m_arbiter.wb0_adr\[17\] sspi.req_addr\[17\] _1399_ _1491_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2122_ _0736_ _0745_ _0746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2053_ wb_compressor.wb_i_dat\[14\] wb_cross_clk.s_m_sync.s_data_ff\[16\] _0688_
+ _0697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ _0641_ _1346_ _1347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2886_ _1287_ _1290_ _1291_ _0280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1906_ _0525_ _0526_ _0591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3048__S _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2981__A2 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1837_ _0525_ _0526_ _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_13_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3507_ _0272_ clknet_leaf_18_user_clock2 sspi.res_data\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xmax_cap230 _0637_ net230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3531__CLK clknet_leaf_8_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1768_ _0465_ _0466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xmax_cap252 _1328_ net252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1699_ _1563_ _1564_ _0405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3438_ _0218_ clknet_4_15_0_net196 wb_compressor.wb_i_dat\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3369_ _0149_ clknet_leaf_39_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1775__A3 net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1765__I net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2724__A2 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2037__S _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2660__A1 _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2660__B2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1876__S _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2412__A1 net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2740_ _0822_ _1074_ _1158_ _1174_ _1175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_2671_ _0774_ _1116_ _0240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2280__B _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1622_ _1524_ m_arbiter.wb0_o_dat\[2\] _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3223_ net98 _1520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3154_ _1555_ _1400_ _1482_ _0357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2105_ _0699_ iram_latched\[14\] _0732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3085_ _1431_ _1432_ _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2036_ _0676_ _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2938_ _1208_ _0605_ _1265_ _1332_ _1333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_60_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2869_ sspi.req_data\[3\] _1277_ _1278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input66_I m_io_in[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Left_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2890__A1 sspi.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3198__A2 _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3122__A2 _0603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2881__A1 net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3151__S _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1684__A2 _1579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2633__A1 _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3772_ net249 net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3189__A2 _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2723_ _1074_ net496 _1161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2654_ net178 _1072_ _1101_ _1102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2585_ _1049_ _0221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1605_ net237 net147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2169__C _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3206_ _1552_ _1509_ _1510_ _1253_ _0381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2872__A1 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1675__A2 net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3137_ _1473_ _0349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_4_1_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3068_ clk_div.cnt\[0\] clk_div.cnt\[1\] clk_div.cnt\[2\] _1421_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2185__B _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2019_ wb_cross_clk.s_m_sync.s_data_ff\[0\] _0677_ _0679_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2475__I1 _1572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Left_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_17_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_17_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2095__B _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2918__A2 _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2370_ wb_cross_clk.s_m_sync.s_data_ff\[14\] _0888_ _0918_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2717__C _1071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2606__A1 _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2909__A2 _0610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2706_ _1073_ net509 _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2637_ _1077_ _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3056__S _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2568_ wb_compressor.wb_i_dat\[1\] net68 _1039_ _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2499_ _1527_ net1 _0989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input29_I inner_wb_o_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1648__A2 _1564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2448__I1 _0396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2362__C _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_8_0_net196 clknet_0_net196 clknet_4_8_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_34_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1974__S _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_36_Left_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_30_Right_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2128__A3 _0656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Left_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2818__B _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2537__C _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1639__A2 net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__S _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_54_Left_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1811__A2 _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1870_ _0554_ wb_compressor.state\[2\] _0556_ _0557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1884__S _0558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3013__A1 _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3540_ _0305_ clknet_leaf_9_user_clock2 sspi.req_addr\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3295__CLK clknet_4_3_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3471_ _0251_ clknet_4_12_0_net196 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2422_ _0948_ _0159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_63_Left_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2353_ wb_cross_clk.s_m_sync.s_data_ff\[7\] _0891_ _0908_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2284_ net466 _0852_ _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1999_ _1525_ _0596_ net109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2818__A1 sspi.res_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output135_I net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2294__A2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3188__C _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_3_Left_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2285__A2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1879__S _0558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2971_ _1296_ _1336_ sspi.req_addr\[8\] _1359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2283__B _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1922_ _0601_ _0602_ _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_32_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1853_ _0542_ _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_16_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1784_ net96 _0471_ _0481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3523_ _0288_ clknet_leaf_16_user_clock2 sspi.req_data\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3454_ _0234_ clknet_4_3_0_net196 net168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2405_ wb_cross_clk.m_s_sync.s_data_ff\[9\] _0937_ _0940_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_4_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3385_ _0165_ clknet_leaf_38_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[23\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2336_ _0888_ _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__3310__CLK clknet_4_11_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2267_ _0847_ net465 _0846_ _0104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1789__S _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2198_ net414 _0800_ _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2276__A2 _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3460__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input96_I m_io_in[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1787__A1 _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2200__A2 _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2736__B1 _0571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1711__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold31 wb_cross_clk.m_s_sync.s_data_ff\[8\] net418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2503__A3 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold20 _0862_ net407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold42 _0798_ net429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold53 wb_cross_clk.m_s_sync.s_data_ff\[24\] net440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold64 _0805_ net451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold75 wb_cross_clk.m_s_sync.s_data_ff\[27\] net462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold86 _0841_ net473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold97 net523 net484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3216__A1 net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2019__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3333__CLK clknet_4_6_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3170_ _1490_ _0365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2121_ clk_div.cnt\[0\] clk_div.cnt\[1\] clk_div.cnt\[2\] clk_div.cnt\[3\] _0737_
+ clk_div.curr_div\[1\] _0745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_2052_ _0696_ _0041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_65_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2258__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3058__I1 m_arbiter.wb0_o_dat\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2954_ _0619_ sspi.req_addr\[4\] _1345_ _1346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1769__A1 _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2885_ sspi.req_data\[6\] _1290_ _0763_ _1291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1905_ _1587_ _0583_ _0587_ net219 _0590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XPHY_EDGE_ROW_6_Right_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1836_ _1524_ net46 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_53_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1767_ net128 _0463_ _0465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3506_ _0271_ clknet_leaf_18_user_clock2 sspi.res_data\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xmax_cap253 _1266_ net253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1698_ _1570_ net255 net246 _0400_ _0404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3437_ _0217_ clknet_4_15_0_net196 wb_compressor.wb_i_dat\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3368_ _0148_ clknet_leaf_42_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2497__A2 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2319_ net210 _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3299_ _0079_ clknet_4_10_0_net196 wb_cross_clk.m_s_sync.d_data\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input11_I inner_wb_adr[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2249__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_38_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2709__B1 _1148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1982__S _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2098__B _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2660__A2 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3149__S _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2412__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2053__S _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2670_ net180 _1084_ _1115_ _1116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1621_ _1540_ net36 _1541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1691__I _0398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3222_ net65 _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA_input3_I inner_wb_adr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3153_ sspi.req_addr\[8\] _1400_ _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2104_ _0730_ _0731_ _0721_ _0058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3084_ clk_div.cnt\[4\] clk_div.cnt\[5\] clk_div.cnt\[6\] _1423_ _1432_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_2035_ _0687_ _0033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2100__A1 iram_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2937_ sspi.bit_cnt\[4\] _0611_ net92 _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__2403__A2 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1866__I _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2868_ net239 _1275_ _1277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1819_ net77 _0471_ _0511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2799_ _0988_ _1225_ _1226_ _0258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_41_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1914__A1 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input59_I iram_o_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_16_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_16_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_26_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2890__A2 _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3196__C _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2400__I _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2881__A2 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3771_ net249 net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2397__A1 _0933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2722_ wb_cross_clk.m_s_sync.d_data\[18\] _1033_ _1160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_15_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2653_ _1073_ _1096_ _1100_ _1093_ _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_23_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2584_ wb_compressor.wb_i_dat\[9\] net76 _1039_ _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1604_ _1525_ net41 _1528_ _1529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3205_ net175 _1509_ _1510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2321__A1 _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3136_ m_arbiter.wb0_adr\[0\] sspi.req_addr\[0\] _1400_ _1473_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3067_ _1419_ _1420_ _0332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2018_ _0521_ wb_cross_clk.ack_xor_flag _0678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_57_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2421__S _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold150 net390 net537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2560__A1 net487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2312__A1 _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2863__A2 _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_9_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3000__B sspi.req_addr\[17\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2286__B _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2733__C _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer1_I _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2909__A3 _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3031__A2 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _0774_ _1145_ _0245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput200 net200 m_io_out[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2636_ _1072_ _1083_ _1085_ _0660_ _0236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_64_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2567_ _1040_ _0212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2542__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2498_ _0524_ _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3119_ sspi.res_data\[0\] _0607_ _1270_ sspi.res_data\[2\] _1457_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_2_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2781__A1 _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1887__A3 _0571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2836__A2 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2772__A1 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3157__S _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3470_ _0250_ clknet_4_12_0_net196 net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2421_ wb_cross_clk.m_s_sync.s_data_ff\[17\] net136 _0923_ _0948_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2352_ wb_cross_clk.m_wb_i_dat\[5\] _0896_ _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2283_ _0858_ net477 _0846_ _0109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2728__C _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2827__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1998_ _0663_ _0000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2619_ _0543_ _1068_ _1069_ _0235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3599_ _0364_ clknet_leaf_20_user_clock2 m_arbiter.wb0_adr\[15\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input41_I inner_wb_o_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2818__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output128_I net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2373__C _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2754__A1 sspi.state\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2809__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3262__CLK clknet_4_13_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2970_ _0580_ _1358_ _0297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1921_ _0603_ _0605_ _0606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_44_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1852_ net193 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_24_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1783_ iram_latched\[6\] _0457_ _0479_ _0413_ _0480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2745__A1 sspi.state\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3522_ _0287_ clknet_leaf_16_user_clock2 sspi.req_data\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2596__I1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3453_ _0233_ clknet_leaf_0_user_clock2 sspi.sy_clk\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2404_ _1544_ _0934_ _0939_ _0150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3384_ _0164_ clknet_leaf_35_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[22\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2335_ _0893_ _0894_ _0895_ _0125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_4_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2266_ net464 _0829_ _0848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2197_ _0776_ _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__1869__I _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1787__A2 _0483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input89_I m_io_in[32] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2736__A1 _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2736__B2 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold32 _0793_ net419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold10 _0843_ net397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold21 wb_cross_clk.m_s_sync.s_data_ff\[14\] net408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold54 _0830_ net441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold43 wb_cross_clk.m_s_sync.s_data_ff\[23\] net430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold65 wb_cross_clk.m_s_sync.s_data_ff\[12\] net452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold87 wb_cross_clk.m_s_sync.s_data_ff\[16\] net474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold76 _0837_ net463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold98 net520 net485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3216__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__A2 net228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2831__C _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2727__A1 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3628__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2120_ clk_div.curr_div\[2\] _0743_ clk_div.curr_div\[3\] _0744_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2051_ wb_compressor.wb_i_dat\[13\] wb_cross_clk.s_m_sync.s_data_ff\[15\] _0688_
+ _0696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3207__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2953_ _1330_ _1344_ _1345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1904_ _0462_ _0588_ _0589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2884_ _1261_ _1289_ _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1835_ _0522_ _0523_ _0524_ _0525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__2718__A1 net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1766_ net128 _0463_ _0464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xmax_cap221 net222 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3505_ _0270_ clknet_leaf_17_user_clock2 sspi.res_data\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2194__A2 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap232 net233 net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xmax_cap254 _1179_ net254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1697_ net248 _0392_ _0393_ _0403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_3436_ _0216_ clknet_4_15_0_net196 wb_compressor.wb_i_dat\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_15_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_15_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3367_ _0147_ clknet_leaf_42_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2318_ _0394_ _0395_ _0880_ _0883_ _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_32_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3298_ _0078_ clknet_4_10_0_net196 wb_cross_clk.m_s_sync.d_data\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2249_ wb_cross_clk.m_s_sync.d_data\[27\] _0835_ _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2424__S _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output195_I net195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2709__B2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2709__A1 _0566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1932__A2 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3134__A1 net195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput99 net99 c0_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1999__A2 _0596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3003__B _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2948__A1 sspi.bit_cnt\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3300__CLK clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1620_ _1526_ _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_22_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1923__A2 _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3165__S _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2289__B _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3221_ net64 _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3152_ _1481_ _0356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1687__A1 _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2103_ iram_wb_ack net52 _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3083_ clk_div.cnt\[7\] _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2736__C _1171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2034_ wb_compressor.wb_i_dat\[5\] wb_cross_clk.s_m_sync.s_data_ff\[7\] _0677_ _0687_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2939__A1 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2936_ _1330_ _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2867_ _0629_ net239 _1275_ _1276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_45_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1818_ iram_latched\[1\] _0457_ _0509_ _0413_ _0510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_5_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2798_ _0516_ _0520_ _1223_ _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_5_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1749_ wb_cross_clk.m_wb_i_dat\[9\] _0449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2199__B _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1914__A2 _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3419_ _0199_ clknet_leaf_0_user_clock2 wb_cross_clk.m_burst_cnt\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2419__S _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3323__CLK clknet_4_8_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3473__CLK clknet_4_2_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1741__B _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2330__A2 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2094__A1 iram_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1841__A1 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1692__I1 net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3770_ net249 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2397__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2721_ _1554_ net137 _1159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2652_ _0555_ _1097_ _1099_ _1074_ _1100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2583_ _1048_ _0220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1603_ _1527_ m_arbiter.wb0_o_dat\[7\] _1528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_2_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3204_ _1508_ _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3135_ _0761_ _1472_ _0348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3066_ clk_div.cnt\[0\] clk_div.cnt\[1\] _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2017_ _0676_ _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__1683__I1 net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1832__A1 _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2919_ _1287_ _1316_ _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input71_I m_io_in[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold151 net503 net538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2560__A2 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2657__B _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2312__A2 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1823__A1 _0510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1736__B _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2551__A2 _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2303__A2 _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1665__I1 net4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2909__A4 _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2704_ net185 _1084_ net513 _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput201 net201 m_io_out[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2635_ net176 _1084_ _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2566_ wb_compressor.wb_i_dat\[0\] net67 _1039_ _1040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2497_ wb_cross_clk.m_burst_cnt\[0\] _0878_ _0885_ _0987_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3118_ sspi.res_data\[3\] _1200_ _1265_ sspi.res_data\[1\] _1456_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_2_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinterconnect_outer_380 m_io_oeb[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tieh
X_3049_ _1411_ _0323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1887__A4 _0572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2834__C _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1647__I1 net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2420_ _0947_ _0158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2351_ _0905_ _0906_ _0895_ _0130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3173__S _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2282_ net476 _0852_ _0859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1997_ _0543_ _0533_ _0540_ _0662_ _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_43_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3534__CLK clknet_leaf_8_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3598_ _0363_ clknet_leaf_20_user_clock2 m_arbiter.wb0_adr\[14\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2618_ wb_compressor.state\[5\] wb_compressor.state\[2\] _0551_ _1024_ _1069_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_11_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2549_ _1024_ _1025_ _1026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_11_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input34_I inner_wb_o_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3006__B _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2690__A1 net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1920_ sspi.bit_cnt\[2\] net259 _0605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_4
XTAP_TAPCELL_ROW_32_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1851_ wb_compressor.state\[4\] _0534_ _0540_ _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_65_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1782_ wb_compressor.wb_i_dat\[6\] wb_cross_clk.m_wb_i_dat\[6\] _0458_ _0479_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3521_ _0286_ clknet_leaf_19_user_clock2 sspi.req_data\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3452_ _0232_ clknet_leaf_0_user_clock2 sspi.sy_clk\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_14_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_14_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2403_ wb_cross_clk.m_s_sync.s_data_ff\[8\] _0937_ _0939_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3383_ _0163_ clknet_leaf_31_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[21\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2334_ _0579_ _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_4_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2265_ wb_cross_clk.m_s_sync.d_data\[32\] _0835_ _0847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2196_ wb_cross_clk.m_s_sync.d_data\[11\] _0783_ _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2681__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2984__A2 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output140_I net140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold11 wb_cross_clk.m_s_sync.s_data_ff\[26\] net398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold22 _0808_ net409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold55 wb_cross_clk.m_s_sync.s_data_ff\[4\] net442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold44 _0827_ net431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold33 wb_cross_clk.m_s_sync.s_data_ff\[28\] net420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold99 inner_wb_8_burst net486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold66 _0803_ net453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2665__B _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold88 _0812_ net475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold77 wb_cross_clk.m_s_sync.s_data_ff\[32\] net464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2672__A1 _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2727__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ _0695_ _0040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_65_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2663__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2952_ sspi.bit_cnt\[3\] _0610_ _0607_ _1344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_45_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1903_ _0403_ net500 _0407_ _0409_ _0588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2883_ _1288_ _1283_ _1289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1834_ net108 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_52_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2718__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1765_ net127 _0463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xmax_cap222 net223 net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3504_ _0269_ clknet_leaf_18_user_clock2 sspi.res_data\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xmax_cap244 _0747_ net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3128__C1 _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3435_ _0215_ clknet_4_14_0_net196 wb_compressor.wb_i_dat\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xmax_cap255 _0395_ net255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1696_ _1590_ _1594_ _0394_ _0401_ _0402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_40_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3366_ _0146_ clknet_leaf_45_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3297_ _0077_ clknet_4_8_0_net196 wb_cross_clk.m_s_sync.d_data\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2317_ _0881_ wb_cross_clk.prev_ack _0882_ _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2248_ _0770_ _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_25_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2179_ _0786_ net445 _0544_ _0077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2654__A1 net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2406__A1 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2957__A2 _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output188_I net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2709__A2 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3252__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2893__A1 _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1696__A2 _1594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire237_I _1529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2645__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2948__A2 _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3070__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3220_ net237 _1509_ _1517_ _0988_ _0388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3125__A2 net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3151_ m_arbiter.wb0_adr\[7\] sspi.req_addr\[7\] _1478_ _1481_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2102_ _0699_ iram_latched\[13\] _0730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2884__A1 _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3181__S _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3082_ _1419_ _1430_ _0337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2033_ _0686_ _0032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2636__A1 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold131_I _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2935_ _1323_ _1328_ _1330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2866_ _1200_ _0605_ _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1817_ wb_compressor.wb_i_dat\[1\] wb_cross_clk.m_wb_i_dat\[1\] _0458_ _0509_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2797_ sspi.res_data\[0\] _1224_ _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_2_2__f_user_clock2_I clknet_0_user_clock2 vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_1748_ _0447_ _0448_ net112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1679_ _1592_ net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3418_ _0198_ clknet_leaf_1_user_clock2 wb_cross_clk.m_burst_cnt\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3349_ _0129_ clknet_leaf_30_user_clock2 wb_cross_clk.m_wb_i_dat\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2866__A1 _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1841__A2 _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2720_ wb_compressor.state\[5\] wb_compressor.state\[6\] wb_compressor.state\[2\]
+ _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__3298__CLK clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2651_ _1098_ _1099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1602_ _1526_ _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2582_ wb_compressor.wb_i_dat\[8\] net75 _1039_ _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3203_ net241 _0464_ net233 _0658_ _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
X_3134_ net195 _1455_ _1471_ _1454_ _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3065_ clk_div.cnt\[0\] _1419_ _0331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2016_ wb_compressor.wb_ack wb_compressor.wb_err _0676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_54_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Left_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1832__A2 m_arbiter.i_wb0_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2918_ _0605_ _0636_ _1288_ _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2849_ sspi.state\[6\] _0582_ _1221_ _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_5_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1893__I sspi.state\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input64_I la_data_in[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold152 clk_div.clock_sel net539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_14_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold130 clk_div.clock_sel net526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold141 net130 net528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2673__B _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3440__CLK clknet_4_13_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2000__A2 _0590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_13_0_net196 clknet_0_net196 clknet_4_13_0_net196 vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_59_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2703_ _1140_ _1141_ _1143_ _1093_ _1144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2634_ net206 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput202 net202 m_io_out[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2565_ net213 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_2_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2496_ wb_cross_clk.m_burst_cnt\[0\] _0878_ _0986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3313__CLK clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3117_ _0597_ _1179_ _1454_ _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinterconnect_outer_370 mgt_wb_dat_o[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_381 m_io_oeb[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tieh
X_3048_ sspi.req_data\[8\] m_arbiter.wb0_o_dat\[8\] _1402_ _1411_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1805__A2 _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2230__A2 _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1741__A1 _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2297__A2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_0_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3336__CLK clknet_4_1_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_13_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_13_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1732__A1 iram_latched\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2350_ wb_cross_clk.s_m_sync.s_data_ff\[6\] _0891_ _0906_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2281_ wb_cross_clk.m_s_sync.d_data\[37\] _0772_ _0858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2288__A2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Left_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1996_ wb_compressor.state\[5\] wb_compressor.state\[4\] _0662_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_16_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3597_ _0362_ clknet_leaf_20_user_clock2 m_arbiter.wb0_adr\[13\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2617_ _1025_ _1067_ net202 _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2548_ wb_compressor.state\[5\] wb_compressor.state\[2\] _1025_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2479_ wb_cross_clk.m_s_sync.s_data_ff\[45\] _0391_ _0885_ _0978_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input27_I inner_wb_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2279__A2 _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2708__S _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__A2 _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1714__A1 _0405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2690__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2442__A2 _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1850_ _0535_ _0536_ _0538_ _0539_ _0540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_25_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1781_ _0460_ _0478_ net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3520_ _0285_ clknet_leaf_19_user_clock2 sspi.req_data\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3451_ _0231_ clknet_leaf_0_user_clock2 sspi.sy_clk\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_wire1_I net495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2402_ _1548_ _0934_ _0938_ _0149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3382_ _0162_ clknet_leaf_31_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[20\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2101__B _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2333_ wb_cross_clk.s_m_sync.s_data_ff\[1\] _0891_ _0894_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2264_ _0844_ net457 _0846_ _0103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2195_ _0797_ net429 _0794_ _0082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2130__A1 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2327__I _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2681__A2 net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3501__CLK clknet_leaf_16_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2433__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ _0650_ net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2062__I iram_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1944__A1 _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold23 wb_cross_clk.m_s_sync.s_data_ff\[25\] net410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold12 _0834_ net399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold45 wb_cross_clk.m_s_sync.s_data_ff\[6\] net432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold56 _0785_ net443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold34 _0839_ net421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2438__S _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold78 _0848_ net465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold89 wb_cross_clk.m_s_sync.s_data_ff\[37\] net476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold67 wb_cross_clk.m_s_sync.s_data_ff\[17\] net454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_7_Left_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_1_0_net196 clknet_0_net196 clknet_4_1_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_65_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3179__S _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2951_ _0988_ _1342_ _1343_ _0293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1902_ _1587_ _0402_ _0410_ _0586_ _0587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_57_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2882_ _0601_ sspi.bit_cnt\[0\] _1288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_5_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1833_ _1526_ net27 _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_53_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1926__A1 _0609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1764_ _0461_ _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xmax_cap223 net224 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xmax_cap212 net213 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3503_ _0268_ clknet_leaf_17_user_clock2 sspi.res_data\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3128__B1 _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3434_ _0214_ clknet_4_15_0_net196 wb_compressor.wb_i_dat\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xmax_cap256 net257 net256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1695_ _1570_ net255 net247 _0400_ _0401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_0_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3365_ _0145_ clknet_leaf_45_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3296_ _0076_ clknet_4_8_0_net196 wb_cross_clk.m_s_sync.d_data\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2316_ wb_cross_clk.m_burst_cnt\[3\] wb_cross_clk.m_burst_cnt\[2\] wb_cross_clk.m_burst_cnt\[1\]
+ wb_cross_clk.m_burst_cnt\[0\] _0882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2247_ _0833_ net399 _0817_ _0098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1670__B net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2103__A1 iram_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2057__I iram_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2178_ net444 _0777_ _0787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2654__A2 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2406__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input94_I m_io_in[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3119__B1 _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_max_cap227_I net228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3547__CLK clknet_leaf_8_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Right_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3150_ _1480_ _0355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2101_ _0728_ _0729_ _0721_ _0057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3081_ clk_div.cnt\[6\] _1429_ _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1687__A3 _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2032_ wb_compressor.wb_i_dat\[4\] wb_cross_clk.s_m_sync.s_data_ff\[6\] _0677_ _0686_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_37_Right_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2934_ _1327_ net252 sspi.req_addr\[1\] _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2865_ _1272_ _1274_ _1207_ _0276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1816_ _0504_ _0508_ net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_46_Right_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2796_ _1223_ _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_13_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1747_ iram_latched\[10\] _0426_ _0448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1678_ m_arbiter.wb0_adr\[4\] net21 _1522_ _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3417_ _0197_ clknet_leaf_2_user_clock2 wb_cross_clk.m_burst_cnt\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3348_ _0128_ clknet_leaf_29_user_clock2 wb_cross_clk.m_wb_i_dat\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2324__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Right_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3279_ _0060_ clknet_leaf_30_user_clock2 iram_latched\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Right_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_47_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2650_ wb_cross_clk.m_s_sync.d_data\[8\] _1077_ _1078_ wb_cross_clk.m_s_sync.d_data\[4\]
+ _1098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1601_ _1523_ _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_2581_ _1047_ _0219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2160__I _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3202_ net237 _1499_ _1507_ _0623_ _0380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input1_I inner_wb_4_burst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2857__A2 net253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3133_ sspi.state\[1\] _1470_ _0621_ _1471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3064_ net244 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2015_ _0668_ _0670_ _0674_ _0675_ _0025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_57_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2917_ _1314_ _1315_ _1207_ _0287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2848_ net92 _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_5_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3392__CLK clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2779_ _0610_ net259 _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold142 embed_s_ff\[0\] net529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold131 _1560_ net518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold120 _1567_ net507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input57_I iram_o_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2446__S _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2784__A1 _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_12_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Left_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2775__A1 _0603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2702_ _0569_ _1078_ _1142_ _1086_ _1143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_54_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2104__B _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2633_ _0556_ _1076_ _1079_ _1082_ _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xoutput203 net203 m_io_out[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2564_ _0542_ _0533_ _0662_ _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1750__A2 _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2495_ _0634_ _0985_ _0195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3116_ _0621_ _1453_ _0618_ _1454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2774__B _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_360 mgt_wb_dat_o[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_371 mgt_wb_dat_o[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3047_ _1410_ _0322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinterconnect_outer_382 m_io_oeb[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_38_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2518__A1 _0933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1741__A2 wb_compressor.wb_i_dat\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2757__A1 sspi.state\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2509__A1 _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2859__B _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1732__A2 _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2280_ _0856_ net447 _0846_ _0108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3624__263 net263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_35_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3202__C _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1995_ _0660_ _0661_ _0575_ _0001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_7_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2616_ _0575_ _1024_ _1067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3596_ _0361_ clknet_leaf_7_user_clock2 m_arbiter.wb0_adr\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3430__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2547_ wb_compressor.state\[6\] wb_compressor.state\[3\] _1023_ _1024_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__2920__A1 _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2478_ _0977_ _0186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_54_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2739__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2911__A1 _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1803__S _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3219__A2 _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1602__I _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3303__CLK clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1780_ _0462_ _0477_ _0478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_47_user_clock2_I clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3450_ _0230_ clknet_leaf_0_user_clock2 sspi.sy_clk\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2401_ wb_cross_clk.m_s_sync.s_data_ff\[7\] _0937_ _0938_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3381_ _0161_ clknet_leaf_31_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[19\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2902__A1 _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2332_ wb_cross_clk.msy_xor_err _0889_ _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2263_ _0543_ _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2194_ net428 _0777_ _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1940__C _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2130__A2 _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2969__A1 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2969__B2 sspi.req_addr\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Left_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ m_arbiter.wb0_o_dat\[13\] net32 _1540_ _0650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3579_ _0344_ clknet_leaf_49_user_clock2 clk_div.cnt\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold13 wb_cross_clk.m_s_sync.s_xfer_xor_flag net400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold46 _0789_ net433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold24 _0832_ net411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold35 wb_cross_clk.m_s_sync.s_data_ff\[22\] net422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold57 wb_cross_clk.m_s_sync.s_data_ff\[5\] net444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold79 wb_cross_clk.m_s_sync.s_data_ff\[38\] net466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold68 _0814_ net455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output126_I net126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3123__B _0610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3326__CLK clknet_4_6_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2962__B _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Left_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3476__CLK clknet_4_2_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_60_Left_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2202__B _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1699__A1 _1563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2648__B1 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_35_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1871__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2950_ _1336_ _1332_ net251 _1343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_45_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2881_ net92 _0611_ _1287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1901_ wb_compressor.wb_err _1553_ _0585_ _0586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1832_ _1524_ m_arbiter.i_wb0_cyc _0522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1763_ _1590_ _1594_ _0394_ _0401_ _0461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3502_ _0267_ clknet_leaf_16_user_clock2 sspi.res_data\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xmax_cap213 net214 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1926__A2 _0610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1694_ net130 net129 _0400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3433_ _0213_ clknet_4_15_0_net196 wb_compressor.wb_i_dat\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xmax_cap257 _1209_ net257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xmax_cap246 net247 net246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3364_ _0144_ clknet_leaf_1_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3295_ _0075_ clknet_4_3_0_net196 wb_cross_clk.m_s_sync.d_data\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2315_ wb_cross_clk.prev_stb _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2246_ net398 _0829_ _0834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3151__I1 sspi.req_addr\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2177_ wb_cross_clk.m_s_sync.d_data\[5\] _0783_ _0786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input87_I m_io_in[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_23_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2708__I1 net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2333__A2 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2100_ iram_wb_ack net51 _0729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3080_ clk_div.cnt\[4\] clk_div.cnt\[5\] _1423_ _1429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2031_ _0685_ _0031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2097__A1 iram_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3210__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2933_ _0600_ _0611_ _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2107__B _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2864_ sspi.req_data\[2\] _1273_ _1274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1815_ _0462_ _0507_ _0508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2795_ _0582_ _0597_ _1222_ _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_32_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold117_I _1564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1746_ _0428_ wb_compressor.wb_i_dat\[10\] _0412_ _0446_ _0447_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2021__A1 wb_compressor.wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1677_ _1591_ net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2777__B _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3416_ _0196_ clknet_leaf_1_user_clock2 wb_cross_clk.m_burst_cnt\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3347_ _0127_ clknet_leaf_29_user_clock2 wb_cross_clk.m_wb_i_dat\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3278_ _0059_ clknet_leaf_29_user_clock2 iram_latched\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2229_ wb_cross_clk.m_s_sync.d_data\[21\] _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1700__I net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output193_I net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_11_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_11_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3514__CLK clknet_leaf_16_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_11_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1600_ _1524_ _1525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2003__A1 wb_compressor.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2580_ wb_compressor.wb_i_dat\[7\] net74 _1039_ _1047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2554__A2 _1027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_user_clock2_I clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3201_ net174 _1498_ _1507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2306__A2 _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3132_ sspi.resp_err _0617_ _1469_ _1470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3063_ _1418_ _0330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2014_ _0536_ _0668_ wb_compressor.burst_cnt\[2\] _0675_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2916_ _1261_ _1312_ sspi.req_data\[13\] _1315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2847_ _1258_ _1229_ _1259_ _1253_ _0273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_33_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2778_ sspi.bit_cnt\[3\] _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_14_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold110 _1163_ net497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1729_ wb_cross_clk.m_wb_i_dat\[13\] _0433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold143 disable_s_ff\[0\] net530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2545__A2 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold132 _1172_ net519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold121 wb_cross_clk.m_s_sync.s_data_ff\[19\] net517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_1_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1808__A1 _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_52_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1605__I net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2701_ wb_cross_clk.m_s_sync.d_data\[15\] net149 _1033_ _1142_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2632_ _1080_ _1552_ _1081_ _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2563_ _1037_ _0211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ _0922_ net209 _0985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_4_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3115_ net258 _1452_ _1453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3046_ sspi.req_data\[7\] m_arbiter.wb0_o_dat\[7\] _1402_ _1410_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinterconnect_outer_361 mgt_wb_dat_o[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_350 mgt_wb_dat_o[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_372 mgt_wb_dat_o[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_383 m_io_oeb[32] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_18_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3191__A2 _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3126__B _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2757__A2 sspi.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2205__B _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3382__CLK clknet_leaf_31_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ wb_compressor.state\[0\] _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2615_ _1064_ _1066_ _0549_ _0234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3595_ _0360_ clknet_leaf_19_user_clock2 m_arbiter.wb0_adr\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2546_ wb_compressor.state\[4\] wb_compressor.state\[1\] _1023_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
X_2477_ wb_cross_clk.m_s_sync.s_data_ff\[44\] _1571_ _0885_ _0977_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2684__A1 net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3029_ sspi.state\[1\] _1399_ _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_34_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2739__A2 net140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3255__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout250 net168 net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_6_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2675__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2978__A2 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2450__I1 _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2400_ _0885_ _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_24_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3380_ _0160_ clknet_leaf_31_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[18\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2902__A2 _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2331_ _0890_ _0892_ _0721_ _0124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2262_ net456 _0829_ _0845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2666__A1 wb_cross_clk.m_s_sync.d_data\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2193_ wb_cross_clk.m_s_sync.d_data\[10\] _0783_ _0797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_2_1__f_user_clock2 clknet_0_user_clock2 clknet_2_1__leaf_user_clock2 vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold147_I net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3091__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2624__I _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1977_ _0649_ net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_16_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3578_ _0343_ clknet_leaf_49_user_clock2 clk_div.cnt\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2529_ _1008_ _1013_ _0549_ _0201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold14 _0879_ net401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input32_I inner_wb_o_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold25 wb_cross_clk.m_s_sync.s_data_ff\[1\] net412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold36 _0825_ net423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold47 wb_cross_clk.m_s_sync.s_data_ff\[15\] net434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold58 _0787_ net445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold69 wb_cross_clk.m_s_sync.s_data_ff\[31\] net456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output119_I net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3082__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2896__A1 _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1699__A2 _1564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2648__B2 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2648__A1 net142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3073__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2880_ _1260_ _1285_ _1286_ _0279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2820__A1 _0460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3420__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1900_ _1553_ net262 _0585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1831_ wb_compressor.wb_ack _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_32_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2380__S _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1762_ iram_latched\[7\] _0457_ _0459_ _0413_ _0460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_52_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap225 net226 net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3501_ _0266_ clknet_leaf_16_user_clock2 sspi.res_data\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1926__A3 net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1693_ _0399_ net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3208__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3128__A2 _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3432_ _0212_ clknet_4_15_0_net196 wb_compressor.wb_i_dat\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap258 _1181_ net258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xmax_cap247 _0397_ net247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3363_ _0143_ clknet_leaf_1_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3294_ _0074_ clknet_4_1_0_net196 wb_cross_clk.m_s_sync.d_data\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2314_ _1540_ m_arbiter.i_wb0_cyc _0412_ _0526_ _0880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_57_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2245_ wb_cross_clk.m_s_sync.d_data\[26\] _0806_ _0833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2176_ _0784_ net443 _0544_ _0076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_64_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2811__A1 _0492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_10_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_10_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3119__A2 _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Right_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2878__A1 _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2465__S _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3443__CLK clknet_4_5_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_29_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_29_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1608__I net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2030_ wb_compressor.wb_i_dat\[3\] wb_cross_clk.s_m_sync.s_data_ff\[5\] _0677_ _0685_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2932_ _0612_ net253 _1326_ _1327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_57_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2863_ net239 _1271_ _1273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1814_ _0505_ _0506_ _0507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2794_ _1178_ _1190_ _1221_ _1222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1745_ _0445_ _0415_ _0446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1780__A1 _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3316__CLK clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1676_ m_arbiter.wb0_adr\[5\] net22 _1557_ _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3415_ _0195_ clknet_leaf_0_user_clock2 wb_cross_clk.m_new_req_flag vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3346_ _0126_ clknet_leaf_32_user_clock2 wb_cross_clk.m_wb_i_dat\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3277_ _0058_ clknet_leaf_28_user_clock2 iram_latched\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3466__CLK clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2228_ _0820_ _0771_ _0821_ _0774_ _0092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2159_ net482 _0772_ _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_64_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3129__B sspi.bit_cnt\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3060__I1 m_arbiter.wb0_o_dat\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1771__A1 net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap232_I net233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire235_I _1533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1826__A2 _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3200__A1 net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3339__CLK clknet_leaf_5_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1762__A1 iram_latched\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1762__B2 _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3200_ net236 _1499_ _1506_ _0761_ _0379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_38_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3131_ sspi.state\[3\] net492 _0617_ _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3062_ sspi.req_data\[15\] m_arbiter.wb0_o_dat\[15\] _1401_ _1418_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2013_ wb_compressor.burst_cnt\[2\] _0536_ _0668_ _0674_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_18_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2915_ _1295_ _1313_ _1314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2242__A2 _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2846_ sspi.res_data\[15\] _1227_ _1259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2793__A3 _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2777_ _1205_ _1206_ _1207_ _0255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xhold100 _1032_ net487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold144 m_arbiter.wb0_o_dat\[0\] net531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1728_ _0431_ _0432_ net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold133 wb_cross_clk.m_s_sync.s_data_ff\[41\] net527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold111 _1164_ net498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold122 _1582_ net509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1659_ _1574_ _1575_ _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2702__B1 _1142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3329_ _0109_ clknet_4_7_0_net196 wb_cross_clk.m_s_sync.d_data\[37\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1808__A2 _0501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2233__A2 _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3631__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2224__A2 _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2700_ wb_cross_clk.m_s_sync.d_data\[31\] _1080_ _0556_ _1141_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2631_ wb_cross_clk.m_s_sync.d_data\[6\] _1080_ _1077_ _1081_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2562_ wb_compressor.burst_end\[2\] net487 _1027_ _1037_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3216__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2493_ _0984_ _0194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3114_ _1187_ _1451_ _1452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3045_ _1409_ _0321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinterconnect_outer_362 mgt_wb_dat_o[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_351 mgt_wb_dat_o[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_340 m_io_out[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_373 mgt_wb_dat_o[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_384 m_io_oeb[33] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_58_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2829_ net112 _1247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1726__A1 _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input62_I iram_o_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output149_I net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2473__S _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2272__I _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1965__A1 _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1817__S _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2142__A1 _0737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2693__A2 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3527__CLK clknet_leaf_9_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1993_ _0542_ _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_16_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2614_ wb_compressor.state\[5\] wb_compressor.state\[4\] _0666_ _1065_ _1066_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3594_ _0359_ clknet_leaf_20_user_clock2 m_arbiter.wb0_adr\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2545_ _0768_ _0544_ _0208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2476_ _0976_ _0185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2684__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3028_ _1399_ _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_66_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2976__B _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1970__I1 net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2675__A2 net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2902__A3 _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2330_ wb_cross_clk.s_m_sync.s_data_ff\[0\] _0891_ _0892_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2261_ wb_cross_clk.m_s_sync.d_data\[31\] _0835_ _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2666__A2 _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2192_ _0795_ net405 _0794_ _0081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_62_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ m_arbiter.wb0_o_dat\[12\] net31 _1540_ _0649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_19_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3577_ _0342_ clknet_leaf_44_user_clock2 clk_div.cnt\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2528_ _1012_ wb_cross_clk.s_burst_cnt\[1\] _1010_ _1013_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2106__A1 iram_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold26 _0778_ net413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2459_ wb_cross_clk.m_s_sync.s_data_ff\[35\] _1567_ _0964_ _0968_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold15 wb_cross_clk.m_s_sync.s_data_ff\[40\] net402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold37 wb_cross_clk.m_s_sync.s_data_ff\[18\] net424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input25_I inner_wb_adr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2657__A2 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold59 wb_cross_clk.m_s_sync.s_data_ff\[36\] net446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold48 _0810_ net435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2409__A2 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_28_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_62_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2648__A2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2820__A2 _0478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ _0520_ _0516_ net111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_37_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3500_ _0265_ clknet_leaf_16_user_clock2 sspi.res_data\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1761_ wb_compressor.wb_i_dat\[7\] wb_cross_clk.m_wb_i_dat\[7\] _0458_ _0459_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap226 net227 net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap204 _1195_ net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1692_ m_arbiter.wb0_adr\[2\] net19 net388 _0399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xmax_cap259 _0604_ net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3431_ _0211_ clknet_4_0_0_net196 wb_compressor.burst_end\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3362_ _0142_ clknet_leaf_1_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2887__A2 _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2313_ net400 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3293_ _0073_ clknet_4_1_0_net196 wb_cross_clk.m_s_sync.d_data\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2639__A2 _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2244_ _0831_ net411 _0817_ _0097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2175_ net442 _0777_ _0785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3245__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1959_ sspi.state\[4\] _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3629_ rst_cw_sync.reset_sync_ff\[0\] _0020_ clknet_4_0_0_net196 rst_cw_sync.reset_sync_ff\[1\]
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA_output131_I net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1650__S _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2481__S _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1624__I _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3268__CLK clknet_leaf_31_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2931_ _0639_ _1180_ _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2862_ _0629_ _0611_ net239 _1271_ _1272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_38_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1813_ net169 net225 net221 net194 _0506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2793_ sspi.state\[0\] sspi.state\[2\] _0639_ _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1744_ wb_cross_clk.m_wb_i_dat\[10\] _0445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3414_ _0194_ clknet_leaf_21_user_clock2 wb_cross_clk.prev_xor_err vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1675_ net128 net127 _1590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3345_ _0125_ clknet_leaf_21_user_clock2 wb_cross_clk.msy_xor_err vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3276_ _0057_ clknet_leaf_29_user_clock2 iram_latched\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2566__S _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2227_ net484 _0772_ _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2158_ _0770_ _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_17_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2089_ _0719_ _0720_ _0721_ _0053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_24_Right_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input92_I m_io_in[35] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1709__I _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2314__B _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Left_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output179_I net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1771__A2 net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Right_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_48_Left_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_47_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_wire228_I _0474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_57_Left_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1619__I _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Right_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3200__A2 _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2003__A3 _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1762__A2 _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3130_ sspi.bit_cnt\[3\] net242 _1461_ _1464_ _1467_ _1468_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2711__A1 net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2562__I1 net487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Left_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_60_Right_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3061_ _1417_ _0329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2012_ _0673_ _0024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3019__A2 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2914_ _1260_ _1312_ _1313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2845_ net117 _1258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_hold122_I _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2776_ _0579_ _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold101 _1036_ net488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_13_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1727_ iram_latched\[14\] _0426_ _0432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3433__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold134 _1572_ net521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold112 m_arbiter.wb0_we net499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold123 _1150_ net510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold145 split_s_ff\[0\] net532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1658_ m_arbiter.wb0_adr\[18\] net12 _1557_ _1575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2950__A1 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3328_ _0108_ clknet_4_6_0_net196 wb_cross_clk.m_s_sync.d_data\[36\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2702__A1 _0569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2702__B2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3259_ _0040_ clknet_4_5_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2823__I net125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2769__A1 _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3194__A1 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3306__CLK clknet_4_11_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2630_ _1033_ _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_40_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2561_ _0535_ _1027_ net488 _0210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1735__A2 _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2492_ wb_cross_clk.msy_xor_err _0623_ _0984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_49_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3113_ sspi.state\[5\] sspi.state\[7\] _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3044_ sspi.req_data\[6\] m_arbiter.wb0_o_dat\[6\] _1402_ _1409_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinterconnect_outer_352 mgt_wb_dat_o[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_330 la_data_out[62] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_341 m_io_out[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_363 mgt_wb_dat_o[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_374 mgt_wb_dat_o[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_385 m_io_oeb[34] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2999__A1 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2828_ _1245_ _1229_ _1246_ _0917_ _0267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_5_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2759_ _1190_ _1191_ sspi.state\[2\] _1192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2923__A1 _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input55_I iram_o_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2151__A2 _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3329__CLK clknet_4_7_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3479__CLK clknet_leaf_5_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1965__A2 _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2502__B _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2914__A1 _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_4_0_net196 clknet_0_net196 clknet_4_4_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__2142__A2 _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1992_ _0659_ net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3593_ _0358_ clknet_leaf_7_user_clock2 m_arbiter.wb0_adr\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2613_ net250 _0533_ _0540_ _0545_ _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_51_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2905__A1 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2544_ _1022_ _0207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2475_ wb_cross_clk.m_s_sync.s_data_ff\[43\] _1572_ _0885_ _0976_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2133__A2 _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2574__S _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3027_ _1398_ _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_27_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_27_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_62_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2372__A2 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2124__A2 net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire210_I _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2363__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2260_ _0842_ net397 _0817_ _0102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3163__I1 sspi.req_addr\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2191_ net404 _0777_ _0796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1626__A1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1975_ _0648_ net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1929__A2 _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3576_ _0341_ clknet_leaf_44_user_clock2 clk_div.cnt\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2527_ wb_cross_clk.s_burst_cnt\[1\] _1006_ _1012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2458_ _0468_ _0925_ _0967_ _0176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2368__I _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold27 wb_cross_clk.m_s_sync.s_data_ff\[11\] net414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold16 _0865_ net403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold38 _0816_ net425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2389_ wb_cross_clk.m_s_sync.s_data_ff\[3\] _0929_ _0923_ _0930_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold49 wb_cross_clk.m_s_sync.s_data_ff\[34\] net436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1865__A1 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input18_I inner_wb_adr[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3517__CLK clknet_leaf_16_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2987__B sspi.req_addr\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2479__S _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2820__A3 _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1760_ _1553_ _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_52_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1691_ _0398_ net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xmax_cap227 net228 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3430_ net489 clknet_4_0_0_net196 wb_compressor.burst_end\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap238 _1324_ net238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3361_ _0141_ clknet_leaf_23_user_clock2 wb_cross_clk.m_wb_i_dat\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2389__S _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2887__A3 _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2312_ _0634_ _0878_ _0119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_27_Left_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3292_ _0072_ clknet_4_1_0_net196 wb_cross_clk.m_s_sync.d_data\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2188__I _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3136__I1 sspi.req_addr\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2243_ net410 _0829_ _0832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2174_ wb_cross_clk.m_s_sync.d_data\[4\] _0783_ _0784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Left_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2811__A3 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1958_ _0582_ net230 _0638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1889_ _0411_ net491 _0574_ _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_16_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3628_ net264 _0019_ clknet_4_0_0_net196 rst_cw_sync.reset_sync_ff\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_12_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3559_ _0324_ clknet_leaf_21_user_clock2 m_arbiter.wb0_o_dat\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2826__I net126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1829__A1 _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1640__I _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2930_ _1260_ net238 _1325_ _0290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2861_ _0605_ _1270_ _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1812_ net86 _0471_ _0505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2792_ _1217_ _1220_ _1207_ _0257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1743_ _0443_ _0444_ net113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1674_ _1589_ net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_40_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2309__A2 _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3413_ _0193_ clknet_leaf_5_user_clock2 wb_cross_clk.prev_stb vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3344_ _0124_ clknet_leaf_32_user_clock2 wb_cross_clk.msy_xor_ack vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3275_ _0056_ clknet_leaf_29_user_clock2 iram_latched\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2226_ wb_cross_clk.m_s_sync.d_data\[20\] _0820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2157_ _0770_ _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2088_ _0579_ _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2582__S _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2314__C _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input85_I m_io_in[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2720__A2 wb_compressor.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2484__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2505__B _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1635__I _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3235__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2711__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3060_ sspi.req_data\[14\] m_arbiter.wb0_o_dat\[14\] _1401_ _1417_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2011_ wb_compressor.burst_cnt\[1\] _0672_ _0668_ _0673_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3385__CLK clknet_leaf_38_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2913_ _0605_ _0636_ _1282_ _1312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_61_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2844_ _1256_ _1229_ _1257_ _1253_ _0272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_5_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2775_ _0603_ _1204_ _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold113 net107 net508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1726_ _0428_ wb_compressor.wb_i_dat\[14\] _0413_ _0430_ _0431_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xhold102 _0210_ net489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold135 _1168_ net522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold124 wb_cross_clk.m_s_sync.s_data_ff\[21\] net520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1657_ m_arbiter.wb0_adr\[16\] net10 _1557_ _1574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2950__A2 _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2702__A2 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3327_ _0107_ clknet_4_6_0_net196 wb_cross_clk.m_s_sync.d_data\[35\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3258_ _0039_ clknet_4_7_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3189_ net162 _1499_ _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2209_ _0807_ net409 _0794_ _0086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_14_Left_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2769__A2 _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output191_I net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3258__CLK clknet_4_7_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3194__A2 _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2560_ net487 net220 _1027_ _1036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2932__A2 net253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2491_ _0634_ _0880_ _0193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_outer_320 la_data_out[52] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3112_ _1184_ _1450_ _0347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3043_ _1408_ _0320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinterconnect_outer_353 mgt_wb_dat_o[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_331 la_data_out[63] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_342 m_io_out[32] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_386 m_io_oeb[35] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tieh
Xinterconnect_outer_364 mgt_wb_dat_o[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_375 mgt_wb_dat_o[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xclkbuf_leaf_26_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_26_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2827_ sspi.res_data\[9\] _1224_ _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2758_ sspi.state\[3\] sspi.state\[7\] _0617_ _1191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1709_ _1553_ _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__1982__I0 m_arbiter.wb0_o_dat\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2689_ _1086_ _1130_ _1131_ _0556_ _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_10_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input48_I iram_o_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2687__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2678__A1 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2850__A1 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3423__CLK clknet_4_3_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1991_ _0457_ _0658_ _0659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_55_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2453__I1 _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2612_ net250 _1063_ _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3592_ _0357_ clknet_leaf_20_user_clock2 m_arbiter.wb0_adr\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2905__A2 _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2543_ wb_cross_clk.msy_xor_ack _0623_ _1022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_23_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2474_ _0975_ _0184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2669__A1 _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3094__A1 net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3026_ _0524_ net254 _1182_ _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_46_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2444__I1 _1564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3446__CLK clknet_4_7_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2899__A1 _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2190_ wb_cross_clk.m_s_sync.d_data\[9\] _0783_ _0795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1974_ m_arbiter.wb0_o_dat\[11\] net30 _1526_ _0648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2426__I1 net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3319__CLK clknet_4_8_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3575_ _0340_ clknet_leaf_44_user_clock2 clk_div.cnt\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2526_ _1008_ _1011_ _0549_ _0200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2457_ wb_cross_clk.m_s_sync.s_data_ff\[34\] _0923_ _0967_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3469__CLK clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold17 wb_cross_clk.m_s_sync.s_data_ff\[9\] net404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold28 _0801_ net415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2388_ _1525_ net44 _0929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
Xhold39 wb_cross_clk.m_s_sync.s_data_ff\[3\] net426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3067__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3009_ _1332_ net251 _1380_ _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_66_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2290__A2 _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2417__I1 net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1664__S _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2805__A1 _0504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2281__A2 _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_2_Left_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1690_ m_arbiter.wb0_adr\[3\] net20 _1522_ _0398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xmax_cap206 net207 net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xmax_cap239 _1264_ net239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3360_ _0140_ clknet_leaf_23_user_clock2 wb_cross_clk.m_wb_i_dat\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2592__I0 wb_compressor.wb_i_dat\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2311_ net262 net260 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3291_ net539 clknet_leaf_50_user_clock2 clk_div.clock_sel_r vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2242_ wb_cross_clk.m_s_sync.d_data\[25\] _0806_ _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2173_ _0770_ _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_64_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_20_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1957_ _0600_ _0606_ _0636_ _0637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_7_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1783__A1 iram_latched\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1888_ _0563_ _0568_ _0573_ _0574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1783__B2 _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3627_ rst_soc_sync.reset_sync_ff\[2\] _0018_ clknet_leaf_50_user_clock2 net108 vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3558_ _0323_ clknet_leaf_16_user_clock2 m_arbiter.wb0_o_dat\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2509_ _0623_ _0996_ _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3489_ _0254_ clknet_leaf_11_user_clock2 sspi.bit_cnt\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA_input30_I inner_wb_o_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output117_I net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3212__A1 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1829__A2 _0519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2860_ sspi.bit_cnt\[1\] _0602_ _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1811_ iram_latched\[2\] _0457_ _0503_ _0413_ _0504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_41_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2791_ _0639_ _1219_ _1220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1742_ iram_latched\[11\] _0426_ _0444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1673_ m_arbiter.wb0_adr\[0\] net3 _1523_ _1589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3412_ _0192_ clknet_leaf_22_user_clock2 wb_cross_clk.s_m_sync.d_xfer_xor_sync\[2\]
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2190__A1 wb_cross_clk.m_s_sync.d_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3343_ _0123_ clknet_4_8_0_net196 wb_cross_clk.m_s_sync.d_xfer_xor_sync\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3274_ _0055_ clknet_leaf_29_user_clock2 iram_latched\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1831__I wb_compressor.wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2225_ _0818_ _0771_ _0819_ _0774_ _0091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2156_ wb_cross_clk.m_s_sync.d_xfer_xor_sync\[2\] _0769_ _0770_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_49_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2087_ _0703_ net62 _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_5_Right_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2245__A2 _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2989_ _1317_ _1331_ _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_user_clock2_I clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1756__A1 _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input78_I m_io_in[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2837__I _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2236__A2 _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1995__A1 _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2505__C _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1747__A1 iram_latched\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ _0537_ _0536_ _0670_ _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_9_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2227__A2 _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_25_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_25_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2912_ _0634_ _1311_ _0286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1986__A1 _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2843_ sspi.res_data\[14\] _1227_ _1257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2774_ _1195_ _1204_ _1202_ _1205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1725_ _0429_ _0415_ _0430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold103 net526 net490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold114 _0396_ net501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold125 _1558_ net512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold147 net129 net534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold136 wb_cross_clk.m_s_sync.s_data_ff\[30\] net533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1656_ _1570_ _1571_ _1572_ _1573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_21_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3326_ _0106_ clknet_4_6_0_net196 wb_cross_clk.m_s_sync.d_data\[34\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1910__A1 wb_compressor.wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3257_ _0038_ clknet_4_5_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3188_ _1552_ _1499_ _1500_ _0761_ _0373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2208_ net408 _0800_ _0808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2139_ _0751_ _0757_ _0721_ _0067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output184_I net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1901__A1 wb_compressor.wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2457__A2 _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2251__B _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2490_ _0983_ _0192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3111_ m_arbiter.i_wb0_cyc _1183_ _0763_ _1450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinterconnect_outer_310 la_data_out[42] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_332 m_io_oeb[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3042_ sspi.req_data\[5\] m_arbiter.wb0_o_dat\[5\] _1402_ _1408_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinterconnect_outer_321 la_data_out[53] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_343 m_io_out[33] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_365 mgt_wb_dat_o[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_354 mgt_wb_dat_o[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_376 mgt_wb_dat_o[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_387 m_io_out[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_58_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2826_ net126 _1245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2940__I _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2757_ sspi.state\[1\] sspi.state\[6\] _1190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2923__A3 _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1708_ wb_cross_clk.m_wb_i_dat\[15\] _0414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2688_ wb_cross_clk.m_s_sync.d_data\[29\] net493 _1033_ _1131_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3771__I net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1639_ _1523_ net25 _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2136__A1 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2687__A2 net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3309_ _0089_ clknet_4_11_0_net196 wb_cross_clk.m_s_sync.d_data\[17\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2611__A2 wb_compressor.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1667__S _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2678__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2850__A2 _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1990_ _0657_ _0658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_55_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2602__A2 wb_compressor.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3591_ _0356_ clknet_leaf_21_user_clock2 m_arbiter.wb0_adr\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2611_ wb_compressor.state\[1\] wb_compressor.state\[6\] _0665_ _0666_ _1063_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_51_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2905__A3 _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2542_ _0553_ _0678_ _0206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2473_ wb_cross_clk.m_s_sync.s_data_ff\[42\] _1579_ _0964_ _0975_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3243__D net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3248__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3025_ m_arbiter.wb0_we _1397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3032__S _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2841__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3766__I net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2809_ sspi.res_data\[3\] _1224_ _0641_ _1234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input60_I iram_o_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2845__I net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1924__I sspi.bit_cnt\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2520__A1 _0676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3540__CLK clknet_leaf_9_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ _0647_ net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_31_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3574_ _0339_ clknet_leaf_44_user_clock2 clk_div.cnt\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2525_ wb_cross_clk.s_burst_cnt\[0\] _1009_ _1010_ _1011_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2456_ _0966_ _0175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold18 _0796_ net405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold29 wb_cross_clk.m_s_sync.s_data_ff\[7\] net416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2387_ _0779_ _0925_ _0928_ _0144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_39_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3008_ net251 _1380_ sspi.req_addr\[19\] _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_19_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3413__CLK clknet_leaf_5_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2750__A1 _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap207 net208 net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap229 _0425_ net229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2592__I1 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3290_ _0071_ clknet_leaf_43_user_clock2 clk_div.curr_div\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2310_ _0876_ net459 _0549_ _0118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2741__A1 _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2741__B2 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2241_ _0828_ net441 _0817_ _0096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2172_ _0781_ net427 _0544_ _0075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_64_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1956_ _0635_ _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1783__A2 _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3436__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2980__A1 _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1887_ _0569_ _0570_ _0571_ _0572_ _0573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3626_ rst_soc_sync.reset_sync_ff\[1\] _0017_ clknet_leaf_50_user_clock2 rst_soc_sync.reset_sync_ff\[2\]
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_3_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3557_ _0322_ clknet_leaf_13_user_clock2 m_arbiter.wb0_o_dat\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2732__A1 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2508_ _0923_ _0994_ _0995_ _0928_ _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3488_ _0253_ clknet_leaf_12_user_clock2 sspi.bit_cnt\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__2596__S net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2439_ _0957_ _0167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input23_I inner_wb_adr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2395__I _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2799__A1 _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3212__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1774__A2 _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2723__A1 _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3309__CLK clknet_4_11_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_24_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_9_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2254__B _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1649__I net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1810_ wb_compressor.wb_i_dat\[2\] wb_cross_clk.m_wb_i_dat\[2\] _0458_ _0503_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_41_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3459__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2790_ _0600_ _1210_ _1218_ net243 _1219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_26_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1741_ _0428_ wb_compressor.wb_i_dat\[11\] _0412_ _0442_ _0443_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_53_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1672_ _1588_ net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xwire260 net261 net260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3411_ _0191_ clknet_leaf_21_user_clock2 wb_cross_clk.s_m_sync.d_xfer_xor_sync\[1\]
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3342_ _0122_ clknet_4_3_0_net196 wb_cross_clk.m_s_sync.d_xfer_xor_sync\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2190__A2 _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3273_ _0054_ clknet_leaf_30_user_clock2 iram_latched\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_2_0__f_user_clock2_I clknet_0_user_clock2 vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_2224_ net483 _0772_ _0819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_49_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2155_ wb_cross_clk.m_s_sync.d_xfer_xor_sync\[1\] _0769_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2086_ _0699_ iram_latched\[8\] _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3040__S _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2650__B1 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2988_ _1369_ _1370_ _1335_ _0303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3774__I net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1939_ _0622_ _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3609_ _0374_ clknet_leaf_28_user_clock2 net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput90 m_io_in[33] net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2705__A1 _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2181__A2 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3130__A1 sspi.bit_cnt\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2339__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2641__B1 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Right_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_27_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1747__A2 _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2944__A1 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_Right_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3121__B2 sspi.res_data\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3121__A1 sspi.res_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Left_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2911_ _1295_ _1309_ _1310_ sspi.req_data\[12\] _1311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1986__A2 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2842_ net116 _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3188__A1 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2773_ _1189_ _1203_ _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1738__A2 _0440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1724_ wb_cross_clk.m_wb_i_dat\[14\] _0429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_44_Left_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold104 _0530_ net491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold126 _1144_ net513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold115 _1138_ net502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold148 irq_s_ff\[0\] net535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1655_ m_arbiter.wb0_adr\[21\] net16 _1523_ _1572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold137 _1561_ net524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_1_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3325_ _0105_ clknet_4_8_0_net196 wb_cross_clk.m_s_sync.d_data\[33\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3256_ _0037_ clknet_4_13_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1910__A2 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2207_ wb_cross_clk.m_s_sync.d_data\[14\] _0806_ _0807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3187_ net151 _1499_ _1500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_53_Left_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3769__I net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2138_ clk_div.next_div_val _0756_ _0757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2069_ _0703_ net56 _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input90_I m_io_in[33] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Left_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output177_I net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_15_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2848__I net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap223_I net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1901__A2 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2701__I1 net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__S _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3185__A4 _0658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3110_ _1419_ _1449_ _0346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinterconnect_outer_300 la_data_out[32] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_311 la_data_out[43] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_333 m_io_oeb[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3041_ _1407_ _0319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinterconnect_outer_322 la_data_out[54] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_344 m_io_out[34] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2694__S _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_366 mgt_wb_dat_o[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_355 mgt_wb_dat_o[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_377 mgt_wb_dat_o[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1656__A1 _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2707__B _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2825_ _1243_ _1229_ _1244_ _0917_ _0266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_6_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold120_I _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2908__A1 _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2756_ _1188_ _1189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2161__C _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1707_ _0412_ _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__2384__A2 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2687_ _1073_ net237 _1129_ _1130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1638_ m_arbiter.wb0_adr\[8\] _1555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2136__A2 _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3308_ _0088_ clknet_4_11_0_net196 wb_cross_clk.m_s_sync.d_data\[16\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3239_ net89 clknet_leaf_3_user_clock2 disable_s_ff\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2617__B net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_28_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2375__A2 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2602__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2610_ _0634_ _0581_ _0233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3590_ _0355_ clknet_leaf_7_user_clock2 m_arbiter.wb0_adr\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2366__A2 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2541_ _0553_ _0680_ _0205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2472_ _0974_ _0183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2488__I _0982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2118__A2 _0740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1877__A1 _0560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3024_ _0580_ _1396_ _0313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_54_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1801__A1 _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2172__B _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2808_ _0498_ _0502_ _1227_ _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_6_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2900__B _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2739_ _1554_ net140 _1174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input53_I iram_o_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_16_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3342__CLK clknet_4_3_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1678__S _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1643__I1 net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2082__B _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2257__B _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1972_ m_arbiter.wb0_o_dat\[10\] net29 _1526_ _0647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_31_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_49_Right_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3573_ _0338_ clknet_leaf_44_user_clock2 clk_div.cnt\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2524_ wb_cross_clk.s_burst_cnt\[0\] net240 _1010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2455_ wb_cross_clk.m_s_sync.s_data_ff\[33\] _1581_ _0964_ _0966_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold19 wb_cross_clk.m_s_sync.s_data_ff\[39\] net406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2386_ _1527_ net1 net210 _0928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_39_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_58_Right_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3007_ _1382_ _1383_ _1384_ _0308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2814__A3 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3777__I net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_Right_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1760__I _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_23_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_23_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2805__A3 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2018__A1 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap208 _1071_ net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2032__S _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1935__I net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2240_ net440 _0829_ _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2171_ net426 _0777_ _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_64_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1955_ _0608_ _0611_ _0635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1886_ wb_cross_clk.m_s_sync.d_data\[43\] net521 _0559_ _0572_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3038__S _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2980__A2 _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3625_ rst_soc_sync.reset_sync_ff\[0\] _0016_ clknet_leaf_50_user_clock2 rst_soc_sync.reset_sync_ff\[1\]
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3556_ _0321_ clknet_leaf_14_user_clock2 m_arbiter.wb0_o_dat\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2732__A2 _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2507_ _0933_ _0926_ _0995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3487_ _0252_ clknet_leaf_5_user_clock2 sspi.resp_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2438_ wb_cross_clk.m_s_sync.s_data_ff\[25\] net130 _0949_ _0957_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2369_ _0441_ _0889_ _0916_ _0917_ _0137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input16_I inner_wb_adr[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2360__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2971__A2 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2487__A1 _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3203__A3 net233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1740_ _0441_ _0415_ _0442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwire261 _0593_ net261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2270__B _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1671_ m_arbiter.wb0_adr\[1\] net14 net388 _1588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3410_ _0190_ clknet_leaf_47_user_clock2 wb_cross_clk.s_m_sync.d_xfer_xor_sync\[0\]
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3341_ _0121_ clknet_4_0_0_net196 wb_cross_clk.m_s_sync.d_xfer_xor_sync\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2714__A2 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I inner_wb_adr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3272_ _0053_ clknet_leaf_30_user_clock2 iram_latched\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2223_ wb_cross_clk.m_s_sync.d_data\[19\] _0818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_49_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2154_ wb_cross_clk.m_s_sync.d_data\[0\] _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2085_ _0717_ _0718_ _0631_ _0052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3403__CLK clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2987_ _1312_ _1351_ sspi.req_addr\[13\] _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2402__A1 _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1938_ _0524_ _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_1869_ _0555_ _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3608_ _0373_ clknet_leaf_28_user_clock2 net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput80 m_io_in[22] net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput91 m_io_in[34] net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3539_ _0304_ clknet_leaf_11_user_clock2 sspi.req_addr\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output122_I net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3030__I _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1995__A3 _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3197__A2 _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3121__A2 net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_7_0_net196 clknet_0_net196 clknet_4_7_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__2880__A1 _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3426__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2910_ _1208_ _1202_ net259 _1294_ _1310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_9_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2632__A1 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2841_ _1254_ _1229_ _1255_ _1253_ _0271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3188__A2 _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2772_ _1202_ net243 _0603_ _1203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3096__B _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1723_ _1553_ _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xhold116 net536 net511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_13_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold105 net108 net503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold149 net508 net536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold138 _1176_ net525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1654_ m_arbiter.wb0_adr\[22\] net17 _1523_ _1571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold127 wb_cross_clk.m_s_sync.s_data_ff\[20\] net523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_0_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2699__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3324_ _0104_ clknet_4_8_0_net196 wb_cross_clk.m_s_sync.d_data\[32\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3255_ _0036_ clknet_4_15_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2206_ _0770_ _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3186_ _1498_ _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2871__A1 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2137_ _0747_ _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_48_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2068_ _0700_ iram_latched\[2\] _0707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input83_I m_io_in[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3449__CLK clknet_4_6_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2862__A1 _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2085__B _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2090__A2 iram_latched\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3136__S _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_301 la_data_out[33] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3040_ sspi.req_data\[4\] m_arbiter.wb0_o_dat\[4\] _1402_ _1407_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinterconnect_outer_312 la_data_out[44] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_323 la_data_out[55] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_334 m_io_oeb[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_345 m_io_out[35] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_367 mgt_wb_dat_o[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_356 mgt_wb_dat_o[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_378 mgt_wb_dat_o[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1656__A2 _1571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2824_ sspi.res_data\[8\] _1224_ _1244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2755_ sspi.state\[6\] _0639_ _1187_ _1188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_14_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1706_ _0411_ _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2686_ wb_cross_clk.m_s_sync.d_data\[13\] _1074_ _1129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3046__S _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1853__I _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1637_ _1553_ _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_18_Left_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3307_ _0087_ clknet_4_11_0_net196 wb_cross_clk.m_s_sync.d_data\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3238_ net529 clknet_leaf_13_user_clock2 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3169_ m_arbiter.wb0_adr\[16\] sspi.req_addr\[16\] _1399_ _1490_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_1_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2633__B _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3021__A1 _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2127__A3 _0409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2438__I1 net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2063__A2 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1938__I _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1874__S _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2540_ _0553_ _1021_ _0204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_51_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2471_ wb_cross_clk.m_s_sync.s_data_ff\[41\] _1583_ _0964_ _0974_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3079__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3023_ _1356_ _1380_ _1395_ sspi.req_addr\[23\] _1396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1801__A2 _0495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2807_ _1231_ _1232_ _0260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3294__CLK clknet_4_1_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2738_ _1072_ net216 _1173_ _0660_ _0250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_41_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2669_ _1093_ _1111_ _1114_ _1115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input46_I inner_wb_stb vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_22_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_22_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2293__A2 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output202_I net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2538__B _0676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2808__A1 _0498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2284__A2 _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1971_ _0646_ net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_31_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3233__A1 m_arbiter.i_wb0_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3572_ _0337_ clknet_leaf_41_user_clock2 clk_div.cnt\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2523_ net240 _1006_ _1009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2454_ _0965_ _0174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2385_ _0925_ _0926_ _0927_ _0143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput1 inner_wb_4_burst net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_39_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2275__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3006_ _0629_ _1383_ _0622_ _1384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_19_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2266__A2 _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2821__B _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xmax_cap209 net210 net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3144__S _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2170_ wb_cross_clk.m_s_sync.d_data\[3\] _0771_ _0781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1701__A1 _0405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3099__B _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3206__A1 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1954_ _0579_ _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_29_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3624_ net263 _0015_ clknet_leaf_50_user_clock2 rst_soc_sync.reset_sync_ff\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_1885_ wb_cross_clk.m_s_sync.d_data\[44\] _1571_ _0558_ _0571_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2980__A3 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3555_ _0320_ clknet_leaf_15_user_clock2 m_arbiter.wb0_o_dat\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2193__A1 wb_cross_clk.m_s_sync.d_data\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2506_ wb_cross_clk.m_burst_cnt\[2\] _0992_ _0994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3486_ _0009_ clknet_leaf_2_user_clock2 sspi.state\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2437_ _0956_ _0166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3332__CLK clknet_4_6_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3054__S _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1861__I _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2368_ _0579_ _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2496__A2 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2299_ wb_cross_clk.m_s_sync.d_data\[43\] _0772_ _0870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1972__S _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3028__I _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput190 net190 m_io_out[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2487__A2 wb_cross_clk.s_m_sync.d_xfer_xor_sync\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3203__A4 _0658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2043__S _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwire240 _1003_ net240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2411__A2 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xwire251 _1341_ net251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1670_ _1569_ _1586_ net90 _1587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xwire262 _0584_ net262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3340_ _0120_ clknet_leaf_50_user_clock2 wb_cross_clk.m_s_sync.s_xfer_xor_flag vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3271_ _0052_ clknet_leaf_30_user_clock2 iram_latched\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2222_ _0815_ net425 _0817_ _0090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_49_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2153_ _0741_ _0759_ _0767_ _0071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2084_ _0703_ net61 _0718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2650__A2 _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2017__I _0676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2986_ _1313_ _1331_ _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2402__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1937_ sspi.state\[0\] _0621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1868_ wb_compressor.state\[3\] _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_32_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput70 m_io_in[13] net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput81 m_io_in[23] net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3607_ _0372_ clknet_leaf_6_user_clock2 m_arbiter.wb0_adr\[23\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1799_ net171 net226 net222 net198 _0494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3538_ _0303_ clknet_leaf_8_user_clock2 sspi.req_addr\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput92 m_io_in[35] net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_40_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1913__A1 _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3469_ _0249_ clknet_4_12_0_net196 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_66_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2641__A2 _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1904__A1 _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_9_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_9_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_46_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2840_ sspi.res_data\[13\] _1227_ _1255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2632__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2771_ sspi.bit_cnt\[2\] _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_14_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1722_ _0417_ _0427_ net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1653_ m_arbiter.wb0_adr\[12\] net6 _1523_ _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
Xhold117 _1564_ net504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold106 _1563_ net493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_9_Right_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold128 _1581_ net515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2699__A2 net512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3323_ _0103_ clknet_4_8_0_net196 wb_cross_clk.m_s_sync.d_data\[31\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3254_ _0035_ clknet_4_13_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2205_ _0804_ net451 _0794_ _0085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3185_ net241 net232 _0466_ _0658_ _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__2871__A2 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2136_ _1539_ _0751_ _0755_ _0066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2067_ _0705_ _0706_ _0631_ _0046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2969_ _1331_ _1356_ _1357_ sspi.req_addr\[7\] _1358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input76_I m_io_in[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2139__A1 _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2862__A2 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1976__I1 net31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2550__A1 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_302 la_data_out[34] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_313 la_data_out[45] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_324 la_data_out[56] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_335 m_io_oeb[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2853__A2 _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_368 mgt_wb_dat_o[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_357 mgt_wb_dat_o[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_346 mgt_wb_ack_o vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1656__A3 _1572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_379 m_io_oeb[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_58_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2823_ net125 _1243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2754_ sspi.state\[1\] sspi.state\[3\] _1187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_hold106_I _1563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1705_ _1587_ _0402_ _0410_ _0411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
X_2685_ _1072_ net505 _1128_ _0660_ _0242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_30_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1636_ net490 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2541__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2392__I1 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3306_ _0086_ clknet_4_11_0_net196 wb_cross_clk.m_s_sync.d_data\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3062__S _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_21_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_21_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3237_ net90 clknet_leaf_3_user_clock2 embed_s_ff\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2844__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3168_ _1489_ _0364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2119_ clk_div.cnt\[4\] clk_div.cnt\[5\] clk_div.cnt\[6\] clk_div.cnt\[7\] _0737_
+ clk_div.curr_div\[1\] _0743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_1_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3099_ clk_div.cnt\[11\] _1440_ _0756_ _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output182_I net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2780__A1 _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1980__S _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_41_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire231_I net233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3012__A2 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3147__S _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1954__I _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2051__S _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2470_ _0973_ _0182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3022_ net230 _1326_ _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3439__CLK clknet_4_13_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2806_ sspi.res_data\[2\] _1229_ _0641_ _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2737_ net191 _1093_ _1173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2762__A1 _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2668_ net487 _1079_ _1113_ _1086_ _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1619_ _1539_ net143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2599_ wb_compressor.state\[1\] wb_compressor.state\[6\] _0543_ _1056_ _1057_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2514__A1 _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input39_I inner_wb_o_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3194__C _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1949__I _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1970_ m_arbiter.wb0_o_dat\[9\] net43 _1540_ _0646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2116__S0 _0737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1885__S _0558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2992__A1 _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ _0336_ clknet_leaf_41_user_clock2 clk_div.cnt\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_24_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2522_ wb_cross_clk.m_s_sync.d_data\[2\] wb_cross_clk.m_s_sync.d_data\[1\] _1004_
+ _1007_ _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_12_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2453_ wb_cross_clk.m_s_sync.s_data_ff\[32\] _1582_ _0964_ _0965_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2384_ wb_cross_clk.m_s_sync.s_data_ff\[1\] _0925_ _0927_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput2 net486 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3005_ _1337_ _1380_ _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3261__CLK clknet_4_7_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2983__A1 _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3769_ net249 net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2586__I1 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1710__A2 _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3215__A2 _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2974__A1 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1777__A2 _0403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2726__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_64_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3206__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ _0578_ _0632_ _0633_ _0003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2965__A1 _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1884_ wb_cross_clk.m_s_sync.d_data\[36\] net518 _0558_ _0570_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3623_ _0388_ clknet_leaf_27_user_clock2 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3554_ _0319_ clknet_leaf_13_user_clock2 m_arbiter.wb0_o_dat\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2193__A2 _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2505_ _0992_ _0993_ _0579_ _0925_ _0197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3485_ _0008_ clknet_leaf_3_user_clock2 sspi.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2436_ wb_cross_clk.m_s_sync.s_data_ff\[24\] net129 _0949_ _0956_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2367_ wb_cross_clk.s_m_sync.s_data_ff\[13\] _0888_ _0916_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_22_Left_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2298_ net461 _0869_ _0549_ _0114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2922__B _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_8_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2184__A2 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput180 net180 m_io_out[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput191 net191 m_io_out[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3133__A1 sspi.state\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1695__A1 _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_user_clock2_I clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire241 _1594_ net241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_53_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2175__A2 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1962__I _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3155__S _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3270_ _0051_ clknet_leaf_31_user_clock2 iram_latched\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2221_ _0543_ _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2152_ clk_div.next_div_buff\[3\] _0759_ _0763_ _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_49_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2083_ _0699_ iram_latched\[7\] _0717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1989__A2 _0656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2985_ _0580_ _1368_ _0302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2938__A1 _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1936_ _0619_ _0618_ _0620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1867_ net84 _0554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1798_ net94 _0471_ _0493_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput71 m_io_in[14] net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput82 m_io_in[24] net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3606_ _0371_ clknet_leaf_7_user_clock2 m_arbiter.wb0_adr\[22\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput60 iram_o_data[6] net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput93 m_io_in[3] net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3537_ _0302_ clknet_leaf_19_user_clock2 sspi.req_addr\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1913__A2 _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2189__B _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3468_ _0248_ clknet_4_12_0_net196 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3399_ _0179_ clknet_leaf_46_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[37\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2419_ wb_cross_clk.m_s_sync.s_data_ff\[16\] net135 _0923_ _0947_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input21_I inner_wb_adr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2917__B _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2636__C _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output108_I net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2929__A1 sspi.req_addr\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2371__C _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1668__A1 _1581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1731__B _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1840__A1 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2770_ _1199_ _1201_ _0895_ _0254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1721_ iram_latched\[15\] _0426_ _0427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2396__A2 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3472__CLK clknet_4_2_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1652_ _1559_ _1562_ _1565_ _1568_ _1569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xhold107 _1132_ net494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2148__A2 _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold118 _1127_ net505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold129 _1156_ net516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_0_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3322_ _0102_ clknet_4_9_0_net196 wb_cross_clk.m_s_sync.d_data\[30\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3253_ _0034_ clknet_4_13_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2204_ net450 _0800_ _0805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3184_ _1577_ _1400_ _1497_ _0372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_20_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_20_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2320__A2 _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2135_ clk_div.next_div_buff\[3\] _0751_ _0755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2066_ _0703_ net55 _0706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1867__I net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2968_ _1210_ _0612_ _1336_ _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_60_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1919_ sspi.bit_cnt\[1\] sspi.bit_cnt\[0\] _0604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2387__A2 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2899_ _1261_ _1301_ sspi.req_data\[9\] _1302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input69_I m_io_in[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_8_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1898__A1 _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_39_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_39_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2366__C _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1978__S _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1822__A1 _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1673__I1 net3 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1726__B _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2550__A2 _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_303 la_data_out[35] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_314 la_data_out[46] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_325 la_data_out[57] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2302__A2 _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2049__S _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinterconnect_outer_336 m_io_oeb[36] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_369 mgt_wb_dat_o[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_358 mgt_wb_dat_o[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_347 mgt_wb_dat_o[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_58_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1664__I1 net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2292__B _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2822_ _1241_ _1242_ _0265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2369__A2 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2753_ _1184_ _1185_ _1186_ _0917_ _0252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_27_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ _0403_ _0404_ _0407_ _0409_ _0410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_2
X_2684_ net182 _1084_ _1128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3169__I1 sspi.req_addr\[16\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1635_ _1552_ net134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_39_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3305_ _0085_ clknet_4_11_0_net196 wb_cross_clk.m_s_sync.d_data\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3236_ _0025_ clknet_4_0_0_net196 wb_compressor.burst_cnt\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3167_ m_arbiter.wb0_adr\[15\] sspi.req_addr\[15\] _1478_ _1489_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3098_ clk_div.cnt\[11\] _1440_ _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2118_ clk_div.curr_div\[2\] _0740_ _0741_ _0742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2049_ wb_compressor.wb_i_dat\[12\] wb_cross_clk.s_m_sync.s_data_ff\[14\] _0688_
+ _0695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_1_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1804__B2 _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1655__I1 net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2221__I _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2891__I _1294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1646__I1 net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2599__A2 wb_compressor.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3163__S _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3021_ _0988_ _1393_ _1394_ _0312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_clkbuf_4_14_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1885__I1 _1571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2805_ _0504_ _0508_ _1227_ _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_41_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2736_ _0556_ _0570_ _0571_ _1079_ _1171_ _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2667_ _1074_ net234 _1112_ _1113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1618_ _1538_ _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2598_ wb_compressor.wb_err _0662_ _0669_ net85 _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_6_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3219_ net201 _1508_ _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2817__A3 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2417__S _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3533__CLK clknet_leaf_8_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2808__A3 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2116__S1 clk_div.curr_div\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2441__A1 _1593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3570_ _0335_ clknet_leaf_43_user_clock2 clk_div.cnt\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_23_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2521_ net240 _1006_ _1007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2796__I _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2452_ net211 _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2383_ _1540_ net2 _0926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XPHY_EDGE_ROW_18_Right_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_67_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput3 inner_wb_adr[0] net3 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3004_ sspi.req_addr\[18\] _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_39_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3406__CLK clknet_leaf_5_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_27_Right_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2036__I _0676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2983__A2 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3768_ net249 net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2719_ _0774_ _1157_ _0247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2735__A2 _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_7_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_7_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input51_I iram_o_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_36_Right_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2499__A1 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output138_I net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2671__A1 _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2974__A2 _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2726__A2 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Right_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1701__A3 _1593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3429__CLK clknet_4_2_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Right_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_64_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2662__A1 net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2414__A1 net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1952_ sspi.state\[6\] _0615_ _0633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1883_ wb_cross_clk.m_s_sync.d_data\[39\] _1584_ _0558_ _0569_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3622_ _0387_ clknet_leaf_27_user_clock2 net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3553_ _0318_ clknet_leaf_14_user_clock2 m_arbiter.wb0_o_dat\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3484_ _0007_ clknet_leaf_2_user_clock2 sspi.state\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2504_ wb_cross_clk.m_burst_cnt\[0\] _0878_ wb_cross_clk.m_burst_cnt\[1\] _0993_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2435_ _0408_ _0925_ _0955_ _0165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2366_ _0445_ _0889_ _0915_ _0580_ _0136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2297_ wb_cross_clk.m_s_sync.d_data\[42\] _0771_ _0869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2653__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2430__S _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput170 net170 m_io_oeb[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput181 net181 m_io_out[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2369__C _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput192 net192 m_io_out[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2892__A1 _0609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire220 _1035_ net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xwire231 net233 net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xwire242 _1458_ net242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3251__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3124__A2 _0603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2220_ net424 _0800_ _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2151_ _0765_ _0759_ _0766_ _0761_ _0070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3171__S _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2295__B _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2082_ _0715_ _0716_ _0631_ _0051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_49_user_clock2_I clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2635__A1 net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2984_ _1309_ _1331_ _1367_ sspi.req_addr\[12\] _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1935_ net92 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_56_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_12_0_net196 clknet_0_net196 clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_4_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1866_ _0542_ _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_31_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput72 m_io_in[15] net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1797_ iram_latched\[4\] _0457_ _0491_ _0413_ _0492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xinput50 iram_o_data[11] net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3605_ _0370_ clknet_leaf_6_user_clock2 m_arbiter.wb0_adr\[21\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput61 iram_o_data[7] net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput94 m_io_in[4] net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput83 m_io_in[25] net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3536_ _0301_ clknet_leaf_19_user_clock2 sspi.req_addr\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3467_ _0247_ clknet_4_12_0_net196 net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_0_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_38_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_38_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3398_ _0178_ clknet_leaf_46_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[36\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2418_ _0946_ _0157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2349_ wb_cross_clk.m_wb_i_dat\[4\] _0896_ _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input14_I inner_wb_adr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2477__I1 _1571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2626__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_0_Right_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1668__A2 _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2093__A2 iram_latched\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1840__A2 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1720_ _0425_ _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xhold108 net538 net506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_1651_ _1566_ _1567_ _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold119 wb_cross_clk.m_s_sync.s_data_ff\[0\] net514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_clkbuf_leaf_37_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3321_ _0101_ clknet_4_9_0_net196 wb_cross_clk.m_s_sync.d_data\[29\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3252_ _0033_ clknet_4_15_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input6_I inner_wb_adr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2856__A1 _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2203_ wb_cross_clk.m_s_sync.d_data\[13\] _0783_ _0804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3183_ sspi.req_addr\[23\] _1400_ _1497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2134_ _1544_ _0751_ _0754_ _0065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2065_ _0700_ iram_latched\[1\] _0705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2608__A1 _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2459__I1 _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2967_ _0606_ _0636_ _1332_ _1356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3297__CLK clknet_4_8_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1918_ _0601_ _0602_ _0603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_2898_ _1208_ _1266_ _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1849_ wb_compressor.burst_end\[2\] wb_compressor.burst_cnt\[2\] _0539_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_8_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3519_ _0284_ clknet_leaf_18_user_clock2 sspi.req_data\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1898__A2 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output120_I net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2862__A4 _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1822__A2 _0513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3024__A1 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinterconnect_outer_304 la_data_out[36] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_315 la_data_out[47] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_326 la_data_out[58] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_59_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinterconnect_outer_337 m_io_oeb[37] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_359 mgt_wb_dat_o[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_348 mgt_wb_dat_o[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2066__A2 net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_25_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout249_I net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2821_ sspi.res_data\[7\] _1224_ _0763_ _1242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2752_ sspi.resp_err _1184_ _1186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1703_ _0408_ net127 _0409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_2683_ _1086_ _1125_ _1126_ _0556_ _1127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1634_ _1551_ _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3304_ _0084_ clknet_4_10_0_net196 wb_cross_clk.m_s_sync.d_data\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3235_ _0024_ clknet_4_0_0_net196 wb_compressor.burst_cnt\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3166_ _1488_ _0363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3097_ _1440_ _1441_ _0341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2117_ clk_div.curr_div\[3\] _0741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2048_ _0694_ _0039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1804__A2 _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3006__A1 _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input81_I m_io_in[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output168_I net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3312__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2377__C _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2296__A2 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2599__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2220__A2 _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1731__A1 _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_50_Left_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3020_ _0619_ _1289_ _1391_ _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2287__A2 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_8_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2804_ _1228_ _1230_ _0259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_0_0_net196 clknet_0_net196 clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_42_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2211__A2 _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2735_ _0820_ _1074_ _1158_ _1170_ _1171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_41_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2666_ wb_cross_clk.m_s_sync.d_data\[10\] _0428_ _1112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3335__CLK clknet_4_4_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_6_user_clock2 clknet_2_0__leaf_user_clock2 clknet_leaf_6_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1617_ _1536_ _1537_ _1538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2597_ _1055_ _0227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3218_ net236 _1509_ _1516_ _0988_ _0387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2278__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3149_ m_arbiter.wb0_adr\[6\] sspi.req_addr\[6\] _1478_ _1480_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3102__B _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2941__B _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1961__A1 _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1713__A1 _0391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2269__A2 _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3218__A1 net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2851__B _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2441__A2 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2992__A3 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2520_ _0676_ _1005_ _1006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1952__A1 sspi.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2451_ _0963_ _0173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2382_ _0885_ _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2298__B _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1704__A1 _0403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput4 inner_wb_adr[10] net4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3003_ _1379_ _1381_ _1335_ _0307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_39_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2680__A2 _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2432__A2 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2983__A3 net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3767_ net249 net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2196__A1 wb_cross_clk.m_s_sync.d_data\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2718_ net188 _1084_ net516 _1157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2649_ wb_cross_clk.m_s_sync.d_data\[24\] net534 _0559_ _1097_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input44_I inner_wb_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2499__A2 net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1840__B _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2428__S _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3500__CLK clknet_leaf_16_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1777__A4 _0409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2111__A1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2662__A2 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2414__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1951_ _0622_ _0598_ _0632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3169__S _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2965__A3 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1882_ _0564_ _0565_ _0566_ _0567_ _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3621_ _0386_ clknet_leaf_27_user_clock2 net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3552_ _0317_ clknet_leaf_13_user_clock2 m_arbiter.wb0_o_dat\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2503_ wb_cross_clk.m_burst_cnt\[1\] wb_cross_clk.m_burst_cnt\[0\] _0878_ _0992_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_11_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3483_ _0006_ clknet_leaf_3_user_clock2 sspi.state\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2434_ wb_cross_clk.m_s_sync.s_data_ff\[23\] _0937_ _0955_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_37_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_37_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2365_ wb_cross_clk.s_m_sync.s_data_ff\[12\] _0888_ _0915_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2296_ net460 _0776_ _0868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3523__CLK clknet_leaf_16_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2405__A2 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1835__B _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput160 net160 m_io_oeb[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3118__B1 _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput171 net171 m_io_oeb[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput182 net182 m_io_out[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput193 net193 m_io_out[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2892__A2 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire210 _0884_ net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xwire243 _1193_ net243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1907__B2 _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2150_ clk_div.curr_div\[2\] _0759_ _0766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2081_ _0703_ net60 _0716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2635__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2983_ _1208_ _1202_ net259 _1336_ _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_8_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2938__A3 _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2399__A1 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1934_ _0581_ sspi.sy_clk\[3\] _0618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
Xinput40 inner_wb_o_dat[6] net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1865_ _0549_ net205 _0012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput73 m_io_in[16] net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1796_ wb_compressor.wb_i_dat\[4\] wb_cross_clk.m_wb_i_dat\[4\] _0458_ _0491_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput51 iram_o_data[12] net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput62 iram_o_data[8] net62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3604_ _0369_ clknet_leaf_4_user_clock2 m_arbiter.wb0_adr\[20\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput95 m_io_in[5] net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3535_ _0300_ clknet_leaf_19_user_clock2 sspi.req_addr\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput84 m_io_in[26] net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_3_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3466_ _0246_ clknet_4_12_0_net196 net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2417_ wb_cross_clk.m_s_sync.s_data_ff\[15\] net149 _0923_ _0946_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3397_ _0177_ clknet_leaf_46_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[35\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2348_ _0903_ _0904_ _0895_ _0129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2279_ net446 _0852_ _0857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2314__A1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1650_ m_arbiter.wb0_adr\[13\] net7 _1522_ _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold109 _1570_ net496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_34_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2553__A1 _1027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3320_ _0100_ clknet_4_11_0_net196 wb_cross_clk.m_s_sync.d_data\[28\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3251_ _0032_ clknet_4_15_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2202_ _0802_ net453 _0794_ _0084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3182_ _1496_ _0371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2133_ clk_div.next_div_buff\[2\] _0751_ _0754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2064_ _0702_ _0704_ _0631_ _0045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_0__f_user_clock2 clknet_0_user_clock2 clknet_2_0__leaf_user_clock2 vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2753__C _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold141_I net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2966_ _1353_ _1355_ _1335_ _0296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_60_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1917_ sspi.bit_cnt\[0\] _0602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_2897_ _0619_ _0636_ _1295_ _1266_ _1300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_44_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1848_ wb_compressor.burst_end\[0\] _0537_ _0538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_12_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1779_ _0472_ _0476_ _0477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2060__I _0701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3518_ _0283_ clknet_leaf_8_user_clock2 sspi.req_data\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3449_ _0229_ clknet_4_6_0_net196 wb_compressor.wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__2847__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3105__B _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2436__S _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1658__I0 m_arbiter.wb0_adr\[18\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2783__A1 _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2535__A1 wb_compressor.wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2838__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2838__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_305 la_data_out[37] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_316 la_data_out[48] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_59_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinterconnect_outer_338 m_io_out[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_349 mgt_wb_dat_o[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_327 la_data_out[59] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_58_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2145__I clk_div.curr_div\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2820_ _0460_ _0478_ _1223_ _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_26_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3015__A2 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2751_ _1527_ _0590_ _1185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3177__S _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_5_user_clock2 clknet_2_0__leaf_user_clock2 clknet_leaf_5_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1702_ net128 _0408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2682_ wb_cross_clk.m_s_sync.d_data\[28\] net504 _1033_ _1126_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1633_ _1549_ _1550_ _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3303_ _0083_ clknet_4_10_0_net196 wb_cross_clk.m_s_sync.d_data\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3234_ _0023_ clknet_4_2_0_net196 wb_compressor.burst_cnt\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3165_ m_arbiter.wb0_adr\[14\] sspi.req_addr\[14\] _1478_ _1488_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3096_ clk_div.cnt\[10\] _1438_ _0756_ _1441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2116_ clk_div.cnt\[12\] clk_div.cnt\[13\] clk_div.cnt\[14\] clk_div.cnt\[15\] _0737_
+ clk_div.curr_div\[1\] _0740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_2047_ wb_compressor.wb_i_dat\[11\] wb_cross_clk.s_m_sync.s_data_ff\[13\] _0688_
+ _0694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1894__I _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2949_ _1336_ net251 sspi.req_addr\[3\] _1342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input74_I m_io_in[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2517__A1 wb_compressor.wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3190__A1 _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1740__A2 _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2508__A1 _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1731__A2 wb_compressor.wb_i_dat\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2119__S0 _0737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1798__A2 _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2995__A1 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2047__I0 wb_compressor.wb_i_dat\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2803_ sspi.res_data\[1\] _1229_ _0641_ _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2747__A1 sspi.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2734_ _1554_ net139 _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2665_ wb_cross_clk.m_s_sync.d_data\[26\] _1080_ _0555_ _1110_ _1111_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_30_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1616_ _1525_ m_arbiter.wb0_o_dat\[3\] _1537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2596_ wb_compressor.wb_i_dat\[15\] net83 net214 _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout249 net250 net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3217_ net200 _1508_ _1516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3148_ _1479_ _0354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3079_ _1419_ _1428_ _0336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2738__A1 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output180_I net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2910__A1 _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1713__A2 _1579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3218__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2977__A1 _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2729__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2450_ wb_cross_clk.m_s_sync.s_data_ff\[31\] _1558_ _0949_ _0963_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_36_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_36_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2381_ _0924_ _0142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput5 inner_wb_adr[11] net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3002_ _1333_ _1380_ _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3209__A2 _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3302__CLK clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2983__A4 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3766_ net249 net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2196__A2 _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2717_ _1152_ _1153_ _1155_ _1071_ _1156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_30_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2648_ net142 _1086_ _1079_ _0931_ _1096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2579_ _1046_ _0218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input37_I inner_wb_o_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2444__S _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1631__A1 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2974__A4 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2187__A2 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1698__A1 _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2111__A2 _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3325__CLK clknet_4_8_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1950_ _0628_ _0630_ _0631_ _0008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1622__A1 _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1881_ wb_cross_clk.m_s_sync.d_data\[45\] _0391_ _0559_ _0567_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3620_ _0385_ clknet_leaf_27_user_clock2 net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3475__CLK clknet_4_3_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3551_ _0316_ clknet_leaf_13_user_clock2 m_arbiter.wb0_o_dat\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1992__I _0659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2178__A2 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2502_ _0986_ _0987_ _0988_ _0991_ _0196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3482_ _0005_ clknet_leaf_2_user_clock2 sspi.state\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2433_ _0463_ _0934_ _0954_ _0164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2364_ _0449_ _0889_ _0914_ _0580_ _0135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1689__A1 _0396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2350__A2 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2295_ net395 _0867_ _0549_ _0113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2638__B1 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2102__A2 iram_latched\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2772__B _0603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2169__A2 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput161 net161 m_io_oeb[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput150 net150 iram_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput194 net194 m_io_out[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput172 net172 m_io_oeb[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput183 net183 m_io_out[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2341__A2 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2947__B _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2892__A3 _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire211 _0884_ net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xwire233 _0470_ net233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3018__B _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2332__A2 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2080_ _0700_ iram_latched\[6\] _0715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1843__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2982_ _0580_ _1366_ _0301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3200__C _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2938__A4 _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2399__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1933_ sspi.state\[5\] _0617_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_26_Left_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput30 inner_wb_o_dat[11] net30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1864_ wb_compressor.state\[4\] _0533_ _0547_ wb_compressor.l_we _0551_ _0552_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3603_ _0368_ clknet_leaf_5_user_clock2 m_arbiter.wb0_adr\[19\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput41 inner_wb_o_dat[7] net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 iram_o_data[13] net52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1795_ _0486_ _0490_ net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput63 iram_o_data[9] net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput96 m_io_in[6] net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput74 m_io_in[17] net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2020__A1 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3534_ _0299_ clknet_leaf_8_user_clock2 sspi.req_addr\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput85 m_io_in[27] net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3465_ _0245_ clknet_4_14_0_net196 net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_10_Left_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2416_ _0945_ _0156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3396_ _0176_ clknet_leaf_46_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[34\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2347_ wb_cross_clk.s_m_sync.s_data_ff\[5\] _0891_ _0904_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2278_ wb_cross_clk.m_s_sync.d_data\[36\] _0835_ _0856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2314__A2 m_arbiter.i_wb0_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1825__B2 _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1825__A1 iram_latched\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1676__I1 net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1600__I _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1756__B _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_4_user_clock2 clknet_2_0__leaf_user_clock2 clknet_leaf_4_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3050__I0 sspi.req_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2002__A1 _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2553__A2 _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3250_ _0031_ clknet_4_11_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_50_user_clock2_I clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2201_ net452 _0800_ _0803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2305__A2 _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3181_ m_arbiter.wb0_adr\[22\] sspi.req_addr\[22\] _1399_ _1496_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2856__A3 net253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2132_ _1548_ _0751_ _0753_ _0064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _0703_ net48 _0704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1816__A1 _0504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1667__I1 net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold134_I _1572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2965_ _0629_ _1354_ _1331_ _1355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_17_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2896_ _0988_ _1297_ _1299_ _0282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1916_ sspi.bit_cnt\[1\] _0601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_17_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1847_ wb_compressor.burst_cnt\[0\] wb_compressor.burst_cnt\[1\] _0537_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1778_ net174 net228 net224 net201 _0476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3517_ _0282_ clknet_leaf_16_user_clock2 sspi.req_data\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3448_ _0228_ clknet_4_6_0_net196 wb_compressor.wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__2497__B _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3379_ _0159_ clknet_leaf_37_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[17\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1658__I1 net12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2535__A2 wb_compressor.wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_306 la_data_out[38] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_317 la_data_out[49] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_59_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinterconnect_outer_328 la_data_out[60] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_339 m_io_out[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_3_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3031__B _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2870__B _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2750_ _0597_ _1183_ _1184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_27_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2681_ _1073_ net236 _1124_ _1125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1701_ _0405_ _0406_ _1593_ _0407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_1632_ _1525_ net531 _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3302_ _0082_ clknet_4_10_0_net196 wb_cross_clk.m_s_sync.d_data\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2110__B _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3233_ m_arbiter.i_wb0_cyc _0523_ _1521_ _0988_ _0389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_55_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3164_ _1487_ _0362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2115_ _0736_ _0738_ _0739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3095_ clk_div.cnt\[10\] _1438_ _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3409__CLK clknet_4_1_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2046_ _0693_ _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2336__I _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2948_ sspi.bit_cnt\[3\] _1200_ _0605_ _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_60_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2879_ sspi.req_data\[5\] _1285_ _0763_ _1286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input67_I m_io_in[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2517__A2 wb_compressor.wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3190__A2 _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1879__I1 _1579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_35_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_35_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2865__B _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2692__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2119__S1 clk_div.curr_div\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_7_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2802_ _1223_ _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_26_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2733_ _1072_ net217 _1169_ _0660_ _0249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_27_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2664_ _1033_ _1593_ _1110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1615_ _1527_ net37 _1536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2595_ _1054_ _0226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1663__C _1579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3216_ net235 _1509_ _1515_ _1253_ _0386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3147_ m_arbiter.wb0_adr\[5\] sspi.req_addr\[5\] _1478_ _1479_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2683__A1 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2683__B2 _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3381__CLK clknet_leaf_31_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3078_ clk_div.cnt\[5\] _1427_ _1428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2029_ _0684_ _0030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2986__A2 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2910__A2 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2674__A1 wb_cross_clk.m_s_sync.d_data\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2977__A2 _1271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2729__A2 net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3254__CLK clknet_4_13_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3154__A2 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2380_ wb_cross_clk.m_s_sync.s_data_ff\[0\] _0922_ _0923_ _0924_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput6 inner_wb_adr[12] net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3001_ _1323_ _1350_ _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_59_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3765_ net249 net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2716_ _0560_ _1078_ _1154_ _1077_ _1155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2647_ _0553_ _1095_ _0237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2578_ wb_compressor.wb_i_dat\[6\] net73 _1039_ _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2656__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2408__A1 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2959__A2 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_13_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2895__A1 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2647__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Left_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Right_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1880_ wb_cross_clk.m_s_sync.d_data\[40\] _1575_ _0558_ _0566_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3550_ _0315_ clknet_leaf_14_user_clock2 m_arbiter.wb0_o_dat\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2501_ _0926_ _0989_ _0990_ _0991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3127__A2 _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Left_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3481_ _0004_ clknet_leaf_3_user_clock2 sspi.state\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_41_Right_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2432_ wb_cross_clk.m_s_sync.s_data_ff\[22\] _0937_ _0954_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2363_ wb_cross_clk.s_m_sync.s_data_ff\[11\] _0896_ _0914_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1689__A2 _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2294_ wb_cross_clk.m_s_sync.d_data\[41\] _0771_ _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2638__A1 net141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2638__B2 _0929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_56_Left_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_50_Right_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_65_Left_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput140 net140 iram_i_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput151 net151 m_io_oeb[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3118__A2 _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput173 net173 m_io_oeb[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput184 net184 m_io_out[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput162 net162 m_io_oeb[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput195 net195 m_io_out[36] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA_output136_I net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2455__S _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2801__A1 _0510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_user_clock2 clknet_2_0__leaf_user_clock2 clknet_leaf_3_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xwire234 _1535_ net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_18_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire245 _0680_ net245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2096__A2 iram_latched\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3442__CLK clknet_4_5_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1843__A2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2981_ _1306_ _1331_ _1365_ sspi.req_addr\[11\] _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2164__I _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1932_ _0578_ _0580_ _0598_ _0616_ _0007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_56_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1863_ _0550_ _0531_ _0551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput31 inner_wb_o_dat[12] net31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 inner_wb_adr[3] net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3602_ _0367_ clknet_leaf_4_user_clock2 m_arbiter.wb0_adr\[18\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput53 iram_o_data[14] net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 inner_wb_o_dat[8] net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1794_ _0462_ _0489_ _0490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput64 la_data_in[0] net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput86 m_io_in[2] net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput97 m_io_in[7] net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput75 m_io_in[18] net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3533_ _0298_ clknet_leaf_8_user_clock2 sspi.req_addr\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3464_ _0244_ clknet_4_14_0_net196 net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2415_ wb_cross_clk.m_s_sync.s_data_ff\[14\] net148 _0923_ _0945_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3395_ _0175_ clknet_leaf_45_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[33\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2346_ wb_cross_clk.m_wb_i_dat\[3\] _0896_ _0903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2277_ _0854_ net439 _0846_ _0107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input97_I m_io_in[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2802__I _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3315__CLK clknet_4_8_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1770__A1 _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3465__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2693__B _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1825__A2 _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2250__A2 _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2200_ wb_cross_clk.m_s_sync.d_data\[12\] _0783_ _0802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3180_ _1495_ _0370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2131_ clk_div.next_div_buff\[1\] _0751_ _0753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2062_ iram_wb_ack _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2069__A2 net56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2964_ net257 _0636_ _1270_ _1354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_57_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1915_ sspi.bit_cnt\[4\] _0600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_60_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2895_ _0619_ _1261_ _1298_ _1299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_8_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1846_ wb_compressor.burst_cnt\[0\] wb_compressor.burst_cnt\[1\] _0536_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3338__CLK clknet_4_1_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1777_ _0473_ _0403_ _0404_ _0409_ _0475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3516_ _0281_ clknet_leaf_10_user_clock2 sspi.req_data\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1752__A1 iram_latched\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Right_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3447_ _0227_ clknet_4_12_0_net196 wb_compressor.wb_i_dat\[15\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3378_ _0158_ clknet_leaf_37_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[16\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2329_ wb_cross_clk.s_m_sync.d_xfer_xor_sync\[2\] wb_cross_clk.s_m_sync.d_xfer_xor_sync\[1\]
+ _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_4
XANTENNA_input12_I inner_wb_adr[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3009__A1 _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2232__A2 _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1991__A1 _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2299__A2 _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_307 la_data_out[39] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_59_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinterconnect_outer_318 la_data_out[50] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_329 la_data_out[61] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_3_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1611__I net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2680_ wb_cross_clk.m_s_sync.d_data\[12\] _1074_ _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1700_ net132 _0406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_30_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1631_ _1527_ net28 _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3630__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3301_ _0081_ clknet_4_10_0_net196 wb_cross_clk.m_s_sync.d_data\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3206__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3232_ _1527_ net27 _1521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input4_I inner_wb_adr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3163_ m_arbiter.wb0_adr\[13\] sspi.req_addr\[13\] _1478_ _1487_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2114_ clk_div.cnt\[8\] clk_div.cnt\[9\] clk_div.cnt\[10\] clk_div.cnt\[11\] _0737_
+ clk_div.curr_div\[1\] _0738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3094_ net244 _1438_ _1439_ _0340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2045_ wb_compressor.wb_i_dat\[10\] wb_cross_clk.s_m_sync.s_data_ff\[12\] _0688_
+ _0693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2214__A2 _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2947_ _1339_ _1340_ _1335_ _0292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2878_ _1261_ _1284_ _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1829_ _0462_ _0519_ _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_25_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2301__B _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2971__B sspi.req_addr\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2463__S _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1716__A1 _0391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_2_3__f_user_clock2_I clknet_0_user_clock2 vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2801_ _0510_ _0514_ _1227_ _1228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_41_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2732_ net190 _1093_ _1169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2663_ _0553_ _1109_ _0239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2594_ wb_compressor.wb_i_dat\[14\] net82 net214 _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1614_ net234 net144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3215_ net199 _1508_ _1515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2132__A1 _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3526__CLK clknet_leaf_9_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3146_ _1399_ _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3077_ clk_div.cnt\[4\] _1423_ _1427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2028_ wb_compressor.wb_i_dat\[2\] wb_cross_clk.s_m_sync.s_data_ff\[4\] _0677_ _0684_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2435__A2 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1946__A1 sspi.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3127__B _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2910__A3 net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2966__B _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1870__B _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap212_I net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2685__C _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2674__A2 _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2977__A3 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2901__A3 _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1704__A4 _0409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput7 inner_wb_adr[13] net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3000_ _1327_ _1350_ sspi.req_addr\[17\] _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2665__A2 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2968__A3 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer2_I _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3764_ clknet_leaf_40_user_clock2 net133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2715_ wb_cross_clk.m_s_sync.d_data\[17\] net136 _0559_ _1154_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_15_0_net196 clknet_0_net196 clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__2630__I _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2646_ net177 _1072_ _1094_ _1095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2577_ _1045_ _0217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_66_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3129_ _1465_ _1466_ sspi.bit_cnt\[3\] _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2408__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_2_user_clock2 clknet_2_0__leaf_user_clock2 clknet_leaf_2_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2895__A2 _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2500_ _0933_ net210 _0990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3480_ _0003_ clknet_leaf_2_user_clock2 sspi.state\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2431_ _0953_ _0163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2362_ _0453_ _0889_ _0913_ _0580_ _0134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_20_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1689__A3 _1581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2293_ net394 _0776_ _0866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3214__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2638__A2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput152 net152 m_io_oeb[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput141 net141 iram_i_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput130 net130 iram_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_clkbuf_leaf_46_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2629_ _1078_ _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput174 net174 m_io_oeb[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput185 net185 m_io_out[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input42_I inner_wb_o_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput163 net163 m_io_oeb[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput196 clknet_4_0_0_net196 m_io_out[37] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output129_I net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2471__S _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xwire235 _1533_ net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xwire224 _0475_ net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2868__A2 _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1614__I net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2980_ _1208_ _1275_ _1336_ _1365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1931_ sspi.state\[5\] _0599_ _0615_ sspi.state\[7\] _0616_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1862_ wb_compressor.state\[6\] _0550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
Xinput10 inner_wb_adr[16] net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 inner_wb_adr[4] net21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3601_ _0366_ clknet_leaf_6_user_clock2 m_arbiter.wb0_adr\[17\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput54 iram_o_data[15] net54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1793_ _0487_ _0488_ _0489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput32 inner_wb_o_dat[13] net32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 inner_wb_o_dat[9] net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2556__A1 _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput76 m_io_in[19] net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3532_ _0297_ clknet_leaf_11_user_clock2 sspi.req_addr\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput98 mgt_wb_rst_i net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput65 la_oenb[0] net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput87 m_io_in[30] net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3463_ _0243_ clknet_4_9_0_net196 net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2414_ net237 _0934_ _0944_ _0155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3394_ _0174_ clknet_leaf_33_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[32\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2345_ _0901_ _0902_ _0895_ _0128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2276_ net438 _0852_ _0855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2795__A1 _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3186__I _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2547__A1 wb_compressor.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2304__B _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_33_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_33_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1770__A2 net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2570__I1 net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2786__A1 sspi.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2389__I1 _0929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2130_ _1552_ _0751_ _0752_ _0063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2061_ _0700_ iram_latched\[0\] _0702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2963_ _1289_ _1351_ sspi.req_addr\[6\] _1353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1914_ _0524_ _0582_ _0599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2894_ sspi.bit_cnt\[3\] _0610_ net259 _1298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1845_ wb_compressor.burst_end\[0\] _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_25_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_3_0_net196 clknet_0_net196 clknet_4_3_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_13_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1776_ _0473_ _0403_ _0404_ _0465_ _0474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3515_ _0280_ clknet_leaf_16_user_clock2 sspi.req_data\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1752__A2 _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3446_ _0226_ clknet_4_7_0_net196 wb_compressor.wb_i_dat\[14\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_22_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3377_ _0157_ clknet_leaf_31_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2328_ wb_cross_clk.msy_xor_ack _0889_ _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2259_ net396 _0829_ _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output196_I clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1991__A2 _0658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1743__A2 _0444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3432__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_308 la_data_out[40] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_59_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinterconnect_outer_319 la_data_out[51] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3582__CLK clknet_leaf_5_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2209__B _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1630_ _1548_ net141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__2879__B _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3300_ _0080_ clknet_4_10_0_net196 wb_cross_clk.m_s_sync.d_data\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2931__A1 _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3231_ _1518_ _1519_ _1520_ _0022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3162_ _1486_ _0361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2113_ clk_div.curr_div\[0\] _0737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3093_ clk_div.cnt\[9\] _1436_ _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2044_ _0692_ _0037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2998__B2 sspi.req_addr\[16\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3305__CLK clknet_4_11_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2946_ _0629_ _1331_ _1337_ _1340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2877_ _1282_ _1283_ _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_10_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1828_ _0518_ _0517_ _0519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3455__CLK clknet_4_3_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1725__A2 _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1759_ _0426_ _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3429_ _0209_ clknet_4_2_0_net196 wb_compressor.l_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2150__A2 _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_5_user_clock2_I clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output111_I net111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1661__A1 _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1716__A2 _1579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3328__CLK clknet_4_6_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3780_ net250 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2800_ _1223_ _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3478__CLK clknet_4_3_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2731_ _0556_ _0561_ _0572_ _1079_ _1167_ _1168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_27_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1955__A2 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2662_ net179 _1072_ _1108_ _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1613_ _1525_ net38 _1534_ _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2593_ _1053_ _0225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2904__A1 _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3214_ net234 _1509_ _1514_ _1253_ _0385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_5_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2132__A2 _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3145_ _1477_ _0353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3076_ _1426_ _0335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2027_ _0683_ _0029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_1_user_clock2 clknet_2_0__leaf_user_clock2 clknet_leaf_1_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_33_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2929_ sspi.req_addr\[0\] _1324_ _0622_ _1325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input72_I m_io_in[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1707__I _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2371__A2 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2910__A4 _1294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3171__I1 sspi.req_addr\[17\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1882__A1 _0564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2222__B _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2362__A2 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2649__S _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 inner_wb_adr[14] net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3763_ clknet_leaf_13_user_clock2 net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ wb_cross_clk.m_s_sync.d_data\[33\] _1080_ _0555_ _1153_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2645_ _1073_ _1087_ _1092_ _1093_ _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_11_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2576_ wb_compressor.wb_i_dat\[5\] net72 _1039_ _1045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2353__A2 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2105__A2 iram_latched\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3128_ sspi.res_data\[15\] _1200_ _0607_ sspi.res_data\[12\] _1265_ sspi.res_data\[13\]
+ _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai222_2
XTAP_TAPCELL_ROW_38_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3059_ _1416_ _0328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2307__B _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2344__A2 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2469__S _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2696__C _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2430_ wb_cross_clk.m_s_sync.s_data_ff\[21\] net140 _0949_ _0953_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2361_ wb_cross_clk.s_m_sync.s_data_ff\[10\] _0896_ _0913_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2292_ _0864_ net403 _0846_ _0112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1689__A4 _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_32_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_32_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2023__A1 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput120 net120 inner_wb_i_dat[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput142 net142 iram_i_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2628_ _0555_ _1077_ _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xoutput131 net131 iram_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput186 net186 m_io_out[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput153 net153 m_io_oeb[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput175 net175 m_io_out[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput164 net164 m_io_oeb[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_11_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2559_ _1033_ _0989_ _1032_ _1034_ _1035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xoutput197 net197 m_io_out[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input35_I inner_wb_o_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2088__I _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1688__I1 net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1837__A1 _0525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2801__A3 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwire214 _1038_ net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwire236 _1531_ net236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_33_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1630__I _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1930_ _0524_ _0614_ _0615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1861_ _0543_ _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput11 inner_wb_adr[17] net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 inner_wb_adr[5] net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3600_ _0365_ clknet_leaf_6_user_clock2 m_arbiter.wb0_adr\[16\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput33 inner_wb_o_dat[14] net33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput44 inner_wb_sel[0] net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1792_ net172 net227 net223 net199 _0488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3531_ _0296_ clknet_leaf_8_user_clock2 sspi.req_addr\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput55 iram_o_data[1] net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2556__A2 _0926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput77 m_io_in[1] net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput66 m_io_in[0] net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput88 m_io_in[31] net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3462_ _0242_ clknet_4_9_0_net196 net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2308__A2 _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2413_ wb_cross_clk.m_s_sync.s_data_ff\[13\] _0937_ _0944_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3393_ _0173_ clknet_leaf_33_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[31\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2344_ wb_cross_clk.s_m_sync.s_data_ff\[4\] _0891_ _0902_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2275_ wb_cross_clk.m_s_sync.d_data\[35\] _0835_ _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2572__S _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2795__A2 _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output141_I net141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2990__B sspi.req_addr\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1625__I _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2060_ _0701_ _0044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2392__S _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2962_ _1349_ _1352_ _1335_ _0295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1913_ _0582_ _0597_ _0598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2893_ _1295_ _1296_ sspi.req_data\[8\] _1297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1844_ _0533_ _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1775_ _0405_ _0406_ net131 _0473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3514_ _0279_ clknet_leaf_16_user_clock2 sspi.req_data\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3445_ _0225_ clknet_4_5_0_net196 wb_compressor.wb_i_dat\[13\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3234__CLK clknet_4_2_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3376_ _0156_ clknet_leaf_31_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2327_ _0888_ _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2258_ wb_cross_clk.m_s_sync.d_data\[30\] _0835_ _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2189_ _0792_ net419 _0794_ _0080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3009__A3 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output189_I net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1646__S _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3193__A2 _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2477__S _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_309 la_data_out[41] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_clkbuf_0_user_clock2_I user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3257__CLK clknet_4_5_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3184__A2 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3230_ _1518_ _1519_ _1520_ _0021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2695__A1 _0564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3161_ m_arbiter.wb0_adr\[12\] sspi.req_addr\[12\] _1478_ _1486_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2112_ clk_div.curr_div\[2\] _0736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2695__B2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3092_ clk_div.cnt\[9\] _1436_ _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2043_ wb_compressor.wb_i_dat\[9\] wb_cross_clk.s_m_sync.s_data_ff\[11\] _0688_ _0692_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_0_user_clock2 clknet_2_0__leaf_user_clock2 clknet_leaf_0_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2945_ sspi.req_addr\[2\] _1338_ _1339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2876_ _1209_ _0635_ _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ net151 net225 net221 net175 _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1758_ _0455_ _0456_ net125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1689_ _0396_ _1558_ _1581_ _1582_ _0397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3428_ _0208_ clknet_4_0_0_net196 wb_cross_clk.prev_xor_newreq vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3359_ _0139_ clknet_leaf_17_user_clock2 wb_cross_clk.m_wb_i_dat\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2989__A2 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1661__A2 net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2610__A1 _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2461__I1 _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2913__A2 _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2677__A1 _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2601__B2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2601__A1 wb_compressor.wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2730_ _0818_ _1074_ _1158_ _1166_ _1167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2661_ _1103_ _1104_ _1107_ _1093_ _1108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_26_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1612_ _1527_ m_arbiter.wb0_o_dat\[4\] _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2592_ wb_compressor.wb_i_dat\[13\] net81 net212 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3213_ net198 _1508_ _1514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2668__A1 net487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__B2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3233__C _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3144_ m_arbiter.wb0_adr\[4\] sspi.req_addr\[4\] _1400_ _1477_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3075_ _0756_ _1425_ _1426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1891__A2 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2026_ wb_compressor.wb_i_dat\[1\] wb_cross_clk.s_m_sync.s_data_ff\[3\] _0677_ _0683_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3422__CLK clknet_4_1_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2580__S _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_17_Left_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2928_ sspi.bit_cnt\[4\] _0611_ _1323_ _1324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_60_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2859_ _1267_ _1269_ _1207_ _0275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input65_I la_oenb[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2659__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1723__I _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1882__A2 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2682__I1 net504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2898__A1 _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 inner_wb_adr[15] net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3445__CLK clknet_4_5_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3075__A1 _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3762_ clknet_leaf_24_user_clock2 net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_31_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_31_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2713_ _1073_ net515 _1152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2644_ net207 _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2575_ _1044_ _0216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2889__A1 _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3127_ sspi.res_data\[14\] _1270_ _1202_ _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3058_ sspi.req_data\[13\] m_arbiter.wb0_o_dat\[13\] _1401_ _1416_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2009_ _0668_ _0670_ _0671_ _0023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3318__CLK clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_6_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3468__CLK clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2993__B sspi.req_addr\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2360_ _0911_ _0912_ _0895_ _0133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2291_ net402 _0852_ _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2099__A2 iram_latched\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Right_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2271__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3220__A1 net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2023__A2 net245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput110 net110 inner_wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_3_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput121 net121 inner_wb_i_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2627_ _0550_ _1025_ _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xoutput143 net143 iram_i_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput132 net132 iram_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput154 net154 m_io_oeb[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput176 net176 m_io_out[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput165 net165 m_io_oeb[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_56_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2558_ wb_cross_clk.m_s_sync.d_data\[2\] _1033_ _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_34_Left_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput198 net198 m_io_out[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput187 net187 m_io_out[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2489_ _0623_ wb_cross_clk.s_m_sync.d_xfer_xor_sync\[1\] _0983_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2731__B1 _0572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input28_I inner_wb_o_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1837__A2 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2318__B _0880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Left_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2262__A2 _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire237 _1529_ net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3062__I1 m_arbiter.wb0_o_dat\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xwire248 _0390_ net248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xwire215 net525 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2988__B _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_52_Left_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_18_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2253__A2 _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1860_ _0545_ _0548_ _0544_ _0013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput12 inner_wb_adr[18] net12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1791_ net95 _0471_ _0487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3202__A1 net237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput34 inner_wb_o_dat[15] net34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput45 inner_wb_sel[1] net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 inner_wb_adr[6] net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3530_ _0295_ clknet_leaf_7_user_clock2 sspi.req_addr\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput78 m_io_in[20] net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput67 m_io_in[10] net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput56 iram_o_data[2] net56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput89 m_io_in[32] net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3461_ _0241_ clknet_4_12_0_net196 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2412_ net236 _0934_ _0943_ _0154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3392_ _0172_ clknet_2_2__leaf_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[30\]
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2343_ wb_cross_clk.m_wb_i_dat\[2\] _0896_ _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2274_ _0851_ net437 _0846_ _0106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1819__A2 _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_12_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2492__A2 _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1989_ _0591_ _0656_ _0657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2483__A2 _0676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2235__A2 _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1746__A1 _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2961_ _1284_ _1351_ sspi.req_addr\[5\] _1352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1912_ _0590_ _0596_ _0522_ _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2892_ _0609_ _1202_ _0607_ _1296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_4_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1843_ net85 net84 _0411_ _0530_ _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_25_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1774_ net97 _0471_ _0472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1737__A1 iram_latched\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3513_ _0278_ clknet_leaf_12_user_clock2 sspi.req_data\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3444_ _0224_ clknet_4_5_0_net196 wb_compressor.wb_i_dat\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3375_ _0155_ clknet_leaf_37_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2326_ wb_cross_clk.s_m_sync.d_xfer_xor_sync\[2\] wb_cross_clk.s_m_sync.d_xfer_xor_sync\[1\]
+ _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__3529__CLK clknet_leaf_9_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2257_ _0840_ net473 _0817_ _0101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2188_ _0543_ _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2217__A2 _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2382__I _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input95_I m_io_in[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2331__B _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1900__A1 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2557__I _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2208__A2 _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2225__C _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2241__B _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3160_ _1485_ _0360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3091_ _1419_ _1436_ _1437_ _0339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2695__A2 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2111_ _0700_ _0631_ _0061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2042_ _0691_ _0036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1958__A1 _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2944_ _1336_ _1337_ _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_hold125_I _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2875_ sspi.bit_cnt\[1\] _0602_ _1282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_44_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ net66 _0471_ _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2383__A1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1757_ iram_latched\[8\] _0426_ _0456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1688_ m_arbiter.wb0_adr\[8\] net25 _1557_ _0396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2578__S _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3427_ _0207_ clknet_leaf_32_user_clock2 wb_cross_clk.prev_xor_ack vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_39_Right_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3358_ _0138_ clknet_leaf_17_user_clock2 wb_cross_clk.m_wb_i_dat\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2309_ net458 _0852_ _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2686__A2 _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3289_ _0070_ clknet_leaf_42_user_clock2 clk_div.curr_div\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input10_I inner_wb_adr[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1657__S _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Right_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2126__A1 _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_Right_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_30_user_clock2 clknet_2_3__leaf_user_clock2 clknet_leaf_30_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2660_ _1029_ _1079_ _1106_ _1086_ _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1611_ net235 net145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2591_ _1052_ _0224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3212_ _1539_ _1509_ _1513_ _1253_ _0384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_5_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2197__I _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__A2 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3143_ _1476_ _0352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3074_ clk_div.cnt\[4\] _1423_ _1425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2025_ _0682_ _0028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2840__A2 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_49_user_clock2 clknet_2_0__leaf_user_clock2 clknet_leaf_49_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2927_ _0639_ _1180_ _1323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_17_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2858_ sspi.req_data\[1\] _1268_ _1269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1809_ _0498_ _0502_ net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2789_ _0600_ _0613_ _1218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input58_I iram_o_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2108__A1 iram_latched\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2659__A2 _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3247__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1882__A3 _0566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2831__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3761_ clknet_leaf_13_user_clock2 net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2712_ _0774_ _1151_ _0246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2643_ _0555_ _1089_ _1091_ _1074_ _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2574_ wb_compressor.wb_i_dat\[4\] net71 _1039_ _1044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_10_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3126_ _1462_ _1463_ _1202_ _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_38_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3057_ _1415_ _0327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2008_ wb_compressor.burst_cnt\[0\] _0668_ _0671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_46_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2121__S0 _0737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__A1 _0926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2565__I net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1791__A2 _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2290_ wb_cross_clk.m_s_sync.d_data\[40\] _0772_ _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_63_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2559__A1 _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3220__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput100 net100 c1_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2626_ _1073_ _0463_ _1075_ _1076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput111 net111 inner_wb_i_dat[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput122 net122 inner_wb_i_dat[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput133 net133 iram_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput177 net177 m_io_out[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput155 net155 m_io_oeb[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput166 net166 m_io_oeb[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2557_ _0559_ _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__2731__A1 _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput144 net144 iram_i_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput199 net199 m_io_out[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput188 net188 m_io_out[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2488_ _0982_ _0191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2731__B2 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2586__S net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3109_ clk_div.cnt\[14\] _1446_ clk_div.cnt\[15\] _1449_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2318__C _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_290 la_data_out[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2798__A1 _0516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xwire205 _0552_ net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3211__A2 _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwire216 net519 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3435__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1665__S _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2970__A1 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3585__CLK clknet_leaf_9_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2228__C _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2244__B _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 inner_wb_adr[19] net13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3202__A2 _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1790_ iram_latched\[5\] _0457_ _0485_ _0413_ _0486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_40_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput24 inner_wb_adr[7] net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput35 inner_wb_o_dat[1] net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 inner_wb_stb net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput68 m_io_in[11] net68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput79 m_io_in[21] net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput57 iram_o_data[3] net57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3460_ _0240_ clknet_4_14_0_net196 net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2411_ wb_cross_clk.m_s_sync.s_data_ff\[12\] _0937_ _0943_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3391_ _0171_ clknet_leaf_36_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[29\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2342_ _0899_ _0900_ _0895_ _0127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2713__A1 _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2273_ net436 _0852_ _0853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3308__CLK clknet_4_11_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3458__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1988_ _0654_ _0655_ _0656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1755__A2 _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2952__A1 sspi.bit_cnt\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2609_ _1062_ _0232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3589_ _0354_ clknet_leaf_20_user_clock2 m_arbiter.wb0_adr\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2704__A1 net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input40_I inner_wb_o_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2180__A2 _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output127_I net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2064__B _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3196__A1 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2943__A1 sspi.bit_cnt\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2171__A2 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3120__A1 _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2960_ _1326_ _1350_ _1351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2891_ _1294_ _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1911_ net218 _0595_ _0412_ _0596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1842_ wb_compressor.state\[6\] _0531_ _0532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1737__A2 _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1773_ _0464_ _0466_ net231 net241 _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3512_ _0277_ clknet_leaf_13_user_clock2 sspi.req_data\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3443_ _0223_ clknet_4_5_0_net196 wb_compressor.wb_i_dat\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2162__A2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3374_ _0154_ clknet_leaf_37_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2325_ _0553_ _0769_ _0123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2256_ net472 _0829_ _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3111__A1 m_arbiter.i_wb0_cyc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2187_ net418 _0777_ _0793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_0_user_clock2 user_clock2 clknet_0_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input88_I m_io_in[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2153__A2 _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2916__A1 _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2144__A2 _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2110_ _0734_ _0735_ _0721_ _0060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3090_ clk_div.cnt\[8\] _1433_ _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2041_ wb_compressor.wb_i_dat\[8\] wb_cross_clk.s_m_sync.s_data_ff\[10\] _0688_ _0691_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2943_ sspi.bit_cnt\[3\] _0605_ _1270_ _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_18_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2874_ _1279_ _1281_ _1207_ _0278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2080__A1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1825_ iram_latched\[0\] _0457_ _0515_ _0413_ _0516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_5_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1756_ _0428_ wb_compressor.wb_i_dat\[8\] _0412_ _0454_ _0455_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_53_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2907__A1 _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2151__C _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1687_ _1560_ _1561_ _1567_ _0395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_0_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3426_ _0206_ clknet_4_14_0_net196 wb_cross_clk.ack_xor_flag vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3357_ _0137_ clknet_leaf_17_user_clock2 wb_cross_clk.m_wb_i_dat\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2135__A2 _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2308_ wb_cross_clk.m_s_sync.d_data\[46\] _0772_ _0876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2594__S net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3288_ _0069_ clknet_leaf_43_user_clock2 clk_div.curr_div\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_56_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2239_ _0776_ _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_67_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2071__A1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2342__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2374__A2 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1610_ _1525_ net39 _1532_ _1533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_2_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2365__A2 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2590_ wb_compressor.wb_i_dat\[12\] net80 net212 _1052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3211_ net197 _1508_ _1513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3165__I1 sspi.req_addr\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3142_ m_arbiter.wb0_adr\[3\] sspi.req_addr\[3\] _1400_ _1476_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3073_ _1419_ _1423_ _1424_ _0334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2024_ wb_compressor.wb_i_dat\[0\] wb_cross_clk.s_m_sync.s_data_ff\[2\] _0677_ _0682_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2926_ _1320_ _1322_ _1207_ _0289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2857_ net239 net253 _1268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1808_ _0462_ _0501_ _0502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2356__A2 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2788_ _1195_ _1216_ sspi.bit_cnt\[4\] _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1739_ wb_cross_clk.m_wb_i_dat\[11\] _0441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3772__I net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2108__A2 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3409_ _0189_ clknet_4_1_0_net196 wb_cross_clk.s_m_sync.s_xfer_xor_flag vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2347__A2 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3147__I1 sspi.req_addr\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1858__A1 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2247__B _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3341__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1881__I1 _0391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3760_ clknet_leaf_24_user_clock2 net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2711_ net187 _1084_ net510 _1151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2642_ _1090_ _1091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2573_ _1043_ _0215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2338__A2 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3125_ sspi.res_data\[8\] net259 _1282_ sspi.res_data\[9\] _1463_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_38_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3056_ sspi.req_data\[12\] m_arbiter.wb0_o_dat\[12\] _1401_ _1415_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2007_ _0540_ _0669_ _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_18_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3767__I net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2121__S1 clk_div.curr_div\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2909_ _0609_ _0610_ _1260_ _0607_ _1309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA_input70_I m_io_in[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2067__B _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_43_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2740__A2 _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput101 net101 dcache_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2625_ wb_cross_clk.m_s_sync.d_data\[22\] _1074_ _1075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput112 net112 inner_wb_i_dat[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput123 net123 inner_wb_i_dat[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput134 net134 iram_i_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_23_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_6_0_net196 clknet_0_net196 clknet_4_6_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xoutput156 net156 m_io_oeb[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput167 net167 m_io_oeb[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_11_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2556_ _0415_ _0926_ _1031_ _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput145 net145 iram_i_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput178 net178 m_io_out[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput189 net189 m_io_out[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_11_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2487_ _0623_ wb_cross_clk.s_m_sync.d_xfer_xor_sync\[0\] _0982_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3387__CLK clknet_leaf_38_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2495__A1 _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3108_ _1419_ _1448_ _0345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinterconnect_outer_280 la_data_out[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3039_ _1406_ _0318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinterconnect_outer_291 la_data_out[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2798__A2 _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2615__B _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwire228 _0474_ net228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwire217 net522 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2722__A2 _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_31_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput25 inner_wb_adr[8] net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput36 inner_wb_o_dat[2] net36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput14 inner_wb_adr[1] net14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2410__A1 net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput47 inner_wb_we net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput69 m_io_in[12] net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput58 iram_o_data[4] net58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2410_ net235 _0934_ _0942_ _0153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2260__B _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3390_ _0170_ clknet_leaf_36_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[28\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2341_ wb_cross_clk.s_m_sync.s_data_ff\[3\] _0891_ _0900_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2713__A2 net515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2272_ _0776_ _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_48_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1987_ _1524_ net499 _0655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2952__A2 _0610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2608_ _0641_ sspi.sy_clk\[1\] _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3588_ _0353_ clknet_leaf_3_user_clock2 m_arbiter.wb0_adr\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3780__I net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2539_ net240 _1020_ _1021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2704__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input33_I inner_wb_o_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2345__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2640__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3196__A2 _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1676__S _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3342__D _0122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_47_user_clock2 clknet_2_0__leaf_user_clock2 clknet_leaf_47_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2890_ sspi.state\[6\] _0582_ _1221_ _1294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1910_ wb_compressor.wb_ack _1553_ _0594_ _0595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1841_ _0521_ _0412_ net491 _0531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__3187__A2 _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1772_ _0468_ _0403_ _0418_ _0469_ _0470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3511_ _0276_ clknet_leaf_12_user_clock2 sspi.req_data\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3442_ _0222_ clknet_4_5_0_net196 wb_compressor.wb_i_dat\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2698__A1 _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3373_ _0153_ clknet_leaf_38_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2324_ _0553_ _0887_ _0122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2255_ wb_cross_clk.m_s_sync.d_data\[29\] _0835_ _0840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2186_ wb_cross_clk.m_s_sync.d_data\[8\] _0783_ _0792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3425__CLK clknet_4_3_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2473__I1 _1579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3775__I net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2689__A1 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2689__B2 _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2613__A1 net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2803__B _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_2_user_clock2_I clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2030__S _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold3 net511 net390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3448__CLK clknet_4_6_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2040_ _0690_ _0035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2852__A1 _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2604__A1 _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2455__I1 _1581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2942_ _1330_ _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_57_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2873_ sspi.req_data\[4\] _1280_ _1281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2080__A2 iram_latched\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1824_ wb_compressor.wb_i_dat\[0\] wb_cross_clk.m_wb_i_dat\[0\] _0415_ _0515_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1755_ _0453_ _0415_ _0454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1686_ _0390_ _0392_ _0393_ _0394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_40_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3036__S _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3425_ _0205_ clknet_4_3_0_net196 wb_cross_clk.err_xor_flag vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3356_ _0136_ clknet_leaf_17_user_clock2 wb_cross_clk.m_wb_i_dat\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3287_ _0068_ clknet_leaf_41_user_clock2 clk_div.curr_div\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2307_ _0874_ net471 _0549_ _0117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2238_ wb_cross_clk.m_s_sync.d_data\[24\] _0806_ _0828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_56_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2169_ net481 _0777_ _0780_ _0774_ _0074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2694__I1 net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2446__I1 _1563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output187_I net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3020__A1 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_wire236_I _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3087__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_3__f_user_clock2 clknet_0_user_clock2 clknet_2_3__leaf_user_clock2 vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3270__CLK clknet_leaf_31_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3210_ _1544_ _1509_ _1512_ _1253_ _0383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_66_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3141_ _1475_ _0351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3072_ clk_div.cnt\[3\] _1421_ _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2023_ _0677_ net245 _0681_ _0027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2428__I1 net139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2925_ sspi.req_data\[15\] _1321_ _1322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2856_ _0629_ net239 net253 _1267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_14_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1807_ _0499_ _0500_ _0501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2787_ _1215_ _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1738_ _0439_ _0440_ net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1669_ _1573_ _1576_ _1580_ _1585_ _1586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_0_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3408_ _0188_ clknet_leaf_5_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[46\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3339_ _0119_ clknet_leaf_5_user_clock2 wb_cross_clk.prev_ack vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2419__I1 net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3293__CLK clknet_4_1_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3232__A1 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2710_ _1146_ _1147_ _1149_ net208 _1150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_30_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1794__A1 _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2641_ wb_cross_clk.m_s_sync.d_data\[7\] _1077_ _1078_ wb_cross_clk.m_s_sync.d_data\[3\]
+ _1090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2572_ wb_compressor.wb_i_dat\[3\] net70 _1039_ _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_10_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3124_ sspi.res_data\[11\] _0603_ _1288_ sspi.res_data\[10\] _1462_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_66_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3055_ _1414_ _0326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2006_ _0533_ _0662_ _0669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2649__I1 net534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2908_ _0634_ _1308_ _0285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2839_ net115 _1254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input63_I iram_o_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire1 net495 net492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2348__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2265__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3214__A1 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2256__A2 _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1767__A1 net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2624_ _0458_ _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput113 net113 inner_wb_i_dat[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput124 net124 inner_wb_i_dat[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput102 net102 ic0_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2716__B1 _1154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput157 net157 m_io_oeb[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput135 net135 iram_i_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput168 net250 m_io_oeb[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2555_ wb_cross_clk.m_s_sync.d_data\[1\] _1553_ _1031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput146 net146 iram_i_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput179 net179 m_io_out[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2486_ _0981_ _0190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3044__S _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3107_ clk_div.cnt\[14\] _1446_ _1448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xinterconnect_outer_270 la_data_out[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3038_ sspi.req_data\[3\] m_arbiter.wb0_o_dat\[3\] _1402_ _1406_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3778__I net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_281 la_data_out[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_292 la_data_out[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_66_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2798__A3 _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwire218 _0592_ net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2631__B _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3331__CLK clknet_4_6_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1930__A1 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2806__B _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2238__A2 _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_46_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_29_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1997__A1 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput15 inner_wb_adr[20] net15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 inner_wb_adr[9] net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput37 inner_wb_o_dat[3] net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2410__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput48 iram_o_data[0] net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput59 iram_o_data[5] net59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2340_ wb_cross_clk.m_wb_i_dat\[1\] _0896_ _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1921__A1 _0603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2271_ wb_cross_clk.m_s_sync.d_data\[34\] _0835_ _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_48_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_5_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1986_ _1526_ net47 _0654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2401__A2 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2952__A3 _0607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1782__S _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2607_ _1061_ _0231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3587_ _0352_ clknet_leaf_8_user_clock2 m_arbiter.wb0_adr\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2538_ _0528_ _1005_ _0676_ _1020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1912__A1 _0590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2469_ wb_cross_clk.m_s_sync.s_data_ff\[40\] _1575_ _0964_ _0973_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input26_I inner_wb_adr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2943__A3 _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1903__A1 _0403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2028__S _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2631__A2 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1840_ _1553_ _0527_ _0529_ _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_53_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3377__CLK clknet_leaf_31_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3510_ _0275_ clknet_leaf_12_user_clock2 sspi.req_data\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1771_ net130 net129 _0469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_25_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3441_ _0221_ clknet_4_13_0_net196 wb_compressor.wb_i_dat\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3372_ _0152_ clknet_leaf_39_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2323_ wb_cross_clk.m_s_sync.d_xfer_xor_sync\[0\] _0887_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2254_ _0838_ net421 _0817_ _0100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2185_ _0790_ net417 _0544_ _0079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ _0645_ net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2386__A1 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output132_I net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2861__A2 _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Left_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold4 net391 inner_ext_irq vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3142__S _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2941_ _1329_ _1334_ _1335_ _0291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2872_ _1202_ _0604_ net239 _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1823_ _0510_ _0514_ net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_44_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1754_ wb_cross_clk.m_wb_i_dat\[8\] _0453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3424_ _0204_ clknet_4_1_0_net196 wb_cross_clk.ack_next_hold vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1685_ _1571_ _1572_ _0393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3355_ _0135_ clknet_leaf_24_user_clock2 wb_cross_clk.m_wb_i_dat\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3286_ _0067_ clknet_leaf_43_user_clock2 clk_div.next_div_val vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2540__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2306_ net470 _0852_ _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2237_ _0826_ net431 _0817_ _0095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_56_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3052__S _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2843__A2 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2176__B _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2168_ wb_cross_clk.m_s_sync.d_data\[2\] _0776_ _0780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3542__CLK clknet_leaf_8_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2099_ _0699_ iram_latched\[12\] _0728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input93_I m_io_in[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1970__S _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Right_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2834__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2598__B2 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2598__A1 wb_compressor.wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2041__S _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1880__S _0558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3140_ m_arbiter.wb0_adr\[2\] sspi.req_addr\[2\] _1400_ _1475_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3071_ clk_div.cnt\[0\] clk_div.cnt\[1\] clk_div.cnt\[2\] clk_div.cnt\[3\] _1423_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__2825__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2022_ wb_cross_clk.s_m_sync.s_data_ff\[1\] _0677_ _0681_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_59_Left_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_39_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Right_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2724__B _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2924_ _0613_ _1295_ _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2855_ _0605_ _1265_ _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_5_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1806_ net170 net226 net222 net197 _0500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2786_ sspi.state\[6\] _1187_ _1214_ _1215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3002__A2 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1737_ iram_latched\[12\] _0426_ _0440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1854__I _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_62_Right_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1668_ _1581_ _1582_ _1583_ _1584_ _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_40_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3407_ _0187_ clknet_leaf_47_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[45\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2513__A1 _0926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2513__B2 _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3338_ _0118_ clknet_4_1_0_net196 wb_cross_clk.m_s_sync.d_data\[46\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1599_ _1523_ _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
X_3269_ _0050_ clknet_leaf_31_user_clock2 iram_latched\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3438__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2809__B _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__I _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3232__A2 net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1794__A2 _0489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2640_ _1554_ _0408_ _1088_ _1089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1875__S _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2571_ _1042_ _0214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2594__I1 net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2743__A1 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_27_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3123_ _1459_ _1460_ _0610_ _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_66_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3054_ sspi.req_data\[11\] m_arbiter.wb0_o_dat\[11\] _1401_ _1414_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_38_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2005_ _0667_ _0668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2907_ _1295_ _1306_ _1307_ sspi.req_data\[11\] _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_18_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2982__A1 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2838_ _1251_ _1229_ _1252_ _1253_ _0270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_5_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2769_ _1200_ _0607_ _1197_ _1201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_41_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2734__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xwire2 _1468_ net495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input56_I iram_o_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_45_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_45_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1759__I _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3260__CLK clknet_4_4_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3214__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2973__A1 _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1776__A2 _0403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2725__A1 _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3603__CLK clknet_leaf_5_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2274__B _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_15_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3205__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2623_ _1554_ _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput114 net114 inner_wb_i_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput125 net125 inner_wb_i_dat[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput103 net103 ic1_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2554_ _0546_ _1027_ _1030_ _0209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2716__B2 _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2716__A1 _0560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput158 net158 m_io_oeb[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput136 net136 iram_i_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput147 net147 iram_i_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput169 net169 m_io_oeb[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2485_ wb_cross_clk.s_m_sync.s_xfer_xor_flag _0623_ _0981_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3106_ _1446_ _1447_ _0344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinterconnect_outer_271 la_data_out[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_3037_ _1405_ _0317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3060__S _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinterconnect_outer_282 la_data_out[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_293 la_data_out[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_19_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwire219 _0589_ net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2955__A1 _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2183__A2 _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1694__A1 net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire211_I _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput16 inner_wb_adr[21] net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput27 inner_wb_cyc net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2946__A1 _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput38 inner_wb_o_dat[4] net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput49 iram_o_data[10] net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2174__A2 _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2270_ _0849_ net449 _0846_ _0105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_48_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1685__A1 _1571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1985_ _0653_ net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2606_ _0641_ sspi.sy_clk\[0\] _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2165__A2 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3586_ _0351_ clknet_leaf_4_user_clock2 m_arbiter.wb0_adr\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1862__I wb_compressor.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2537_ _1018_ _1007_ _1019_ _0660_ _0203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2179__B _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2468_ _0972_ _0181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1912__A2 _0596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2399_ _1552_ _0934_ _0936_ _0148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input19_I inner_wb_adr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3192__C _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2089__B _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1947__I _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1690__I1 net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1770_ _1524_ net6 _0467_ _0468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_8_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1883__S _0558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3440_ _0220_ clknet_4_13_0_net196 wb_compressor.wb_i_dat\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2778__I sspi.bit_cnt\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3371_ _0151_ clknet_leaf_40_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2147__A2 _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2322_ net401 _0544_ _0121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2253_ net420 _0829_ _0839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2184_ net416 _0777_ _0791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_25_Left_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_40_Left_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1830__A1 _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1968_ m_arbiter.wb0_o_dat\[8\] net42 _1540_ _0645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2386__A2 net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3471__CLK clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1899_ wb_cross_clk.msy_xor_err wb_cross_clk.prev_xor_err _0584_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_31_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2138__A2 _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3569_ _0334_ clknet_leaf_41_user_clock2 clk_div.cnt\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output125_I net125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1968__S _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2074__A1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2377__A2 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2129__A2 _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold5 net506 net392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__2039__S _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1878__S _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2940_ _0579_ _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2065__A1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2871_ _1202_ _0619_ _0604_ _1264_ _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_45_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1822_ _0462_ _0513_ _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1753_ _0451_ _0452_ net126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1684_ _0391_ _1579_ _0392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_40_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3423_ _0203_ clknet_4_3_0_net196 wb_cross_clk.s_burst_cnt\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3354_ _0134_ clknet_leaf_24_user_clock2 wb_cross_clk.m_wb_i_dat\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3285_ _0066_ clknet_leaf_43_user_clock2 clk_div.next_div_buff\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2305_ wb_cross_clk.m_s_sync.d_data\[45\] _0772_ _0874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2236_ net430 _0800_ _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2167_ net480 _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2098_ _0726_ _0727_ _0721_ _0056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2192__B _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1654__I1 net17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input86_I m_io_in[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2359__A2 _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_2_1__f_user_clock2_I clknet_0_user_clock2 vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3070_ _1419_ _1421_ _1422_ _0333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2021_ wb_compressor.wb_err wb_cross_clk.err_xor_flag _0680_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2277__B _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2923_ _0629_ _0613_ _1295_ _1320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_33_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2854_ _0601_ sspi.bit_cnt\[0\] _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_17_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1805_ net93 _0471_ _0499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2785_ _0639_ _0636_ _1210_ _1214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2740__B _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1736_ _0428_ wb_compressor.wb_i_dat\[12\] _0412_ _0438_ _0439_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_53_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1667_ m_arbiter.wb0_adr\[17\] net11 _1557_ _1584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3406_ _0186_ clknet_leaf_5_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[44\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1598_ _1522_ _1523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_5_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3337_ _0117_ clknet_4_4_0_net196 wb_cross_clk.m_s_sync.d_data\[45\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3268_ _0049_ clknet_leaf_31_user_clock2 iram_latched\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3199_ net173 _1498_ _1506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_44_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_44_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2219_ wb_cross_clk.m_s_sync.d_data\[18\] _0806_ _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output192_I net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Left_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2504__A2 _0878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire241_I _1594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2560__B _1027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2570_ wb_compressor.wb_i_dat\[2\] net69 _1039_ _1042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_10_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3122_ sspi.res_data\[7\] _0603_ _1288_ sspi.res_data\[6\] _1460_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3053_ _1413_ _0325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2004_ _0577_ _0664_ _0665_ _0666_ _0667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2735__B _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2906_ _1208_ _1294_ _1275_ _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_46_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3058__S _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2837_ _0579_ _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2768_ sspi.bit_cnt\[1\] sspi.bit_cnt\[0\] _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_5_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2699_ _1073_ net512 _1140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1719_ _0418_ _0420_ _0422_ _0423_ _0424_ _0425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__2734__A2 net139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I iram_o_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_11_0_net196 clknet_0_net196 clknet_4_11_0_net196 vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__2364__C _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2670__A1 net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3405__CLK clknet_leaf_5_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1976__S _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_net196 net196 clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2489__A1 _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2047__S _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1886__S _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2964__A2 _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2622_ net206 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput115 net115 inner_wb_i_dat[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput104 net104 inner_clock vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2553_ _1027_ _1029_ _1030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2716__A2 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput126 net126 inner_wb_i_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput159 net159 m_io_oeb[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput137 net137 iram_i_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput148 net148 iram_i_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_10_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2484_ _0553_ _0980_ _0189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3428__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3105_ clk_div.cnt\[13\] _1444_ _0756_ _1447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3036_ sspi.req_data\[2\] m_arbiter.wb0_o_dat\[2\] _1402_ _1405_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinterconnect_outer_272 la_data_out[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_283 la_data_out[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_294 la_data_out[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2652__B2 _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2652__A1 _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1796__S _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2404__A1 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2707__A2 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1694__A2 net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2643__B2 _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2643__A1 _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3199__A2 _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput17 inner_wb_adr[22] net17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 inner_wb_o_dat[0] net28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2946__A2 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput39 inner_wb_o_dat[5] net39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1685__A2 _1572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3161__S _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1984_ clknet_leaf_50_user_clock2 clk_div.res_clk clk_div.clock_sel_r _0653_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2937__A2 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2605_ _1060_ _0230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3585_ _0350_ clknet_leaf_9_user_clock2 m_arbiter.wb0_adr\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2536_ wb_cross_clk.s_burst_cnt\[3\] _1019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3250__CLK clknet_4_11_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2467_ wb_cross_clk.m_s_sync.s_data_ff\[39\] _1584_ _0964_ _0972_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2398_ wb_cross_clk.m_s_sync.s_data_ff\[6\] _0925_ _0936_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2195__B _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3019_ _1354_ _1380_ sspi.req_addr\[22\] _1393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2415__S _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2928__A2 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2616__A1 _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1978__I0 m_arbiter.wb0_o_dat\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3370_ _0150_ clknet_leaf_39_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2321_ _0634_ _0886_ _0120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2252_ wb_cross_clk.m_s_sync.d_data\[28\] _0835_ _0838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2183_ wb_cross_clk.m_s_sync.d_data\[7\] _0783_ _0790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2083__A2 iram_latched\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1830__A2 _0516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1967_ _0638_ _0643_ _0644_ _0004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1898_ _0426_ _0527_ _0583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1873__I _0558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3568_ _0333_ clknet_leaf_41_user_clock2 clk_div.cnt\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2519_ wb_cross_clk.m_s_sync.d_data\[0\] wb_cross_clk.prev_xor_newreq _1005_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3499_ _0264_ clknet_leaf_23_user_clock2 sspi.res_data\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input31_I inner_wb_o_dat[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output118_I net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2074__A2 iram_latched\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3296__CLK clknet_4_8_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3023__B2 sspi.req_addr\[23\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold6 net393 inner_reset vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_58_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2065__A2 iram_latched\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1812__A2 _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2870_ _1276_ _1278_ _1207_ _0277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2055__S _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1821_ _0512_ _0511_ _0513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1752_ iram_latched\[9\] _0426_ _0452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ m_arbiter.wb0_adr\[23\] net18 _1523_ _0391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3422_ _0202_ clknet_4_1_0_net196 wb_cross_clk.s_burst_cnt\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3353_ _0133_ clknet_leaf_26_user_clock2 wb_cross_clk.m_wb_i_dat\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3284_ _0065_ clknet_leaf_42_user_clock2 clk_div.next_div_buff\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2304_ _0872_ net469 _0549_ _0116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_43_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_43_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2235_ wb_cross_clk.m_s_sync.d_data\[23\] _0806_ _0826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2166_ _0775_ net413 _0544_ _0073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2097_ iram_wb_ack net50 _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_3_Right_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2999_ _0580_ _1378_ _0306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input79_I m_io_in[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3198__C _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3311__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2020_ _0677_ _0678_ _0679_ _0026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3461__CLK clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2922_ _1318_ _1319_ _1207_ _0288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1797__A1 iram_latched\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1797__B2 _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2853_ _0635_ _1261_ _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1804_ iram_latched\[3\] _0457_ _0497_ _0413_ _0498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2784_ _0634_ _1213_ _0256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1735_ _0437_ _0415_ _0438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold109_I _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2210__A2 _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1666_ m_arbiter.wb0_adr\[19\] net13 _1557_ _1583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_9_0_net196 clknet_0_net196 clknet_4_9_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_0_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3405_ _0185_ clknet_leaf_5_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[43\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1597_ m_arbiter.o_sel_sig _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_5_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3336_ _0116_ clknet_4_1_0_net196 wb_cross_clk.m_s_sync.d_data\[44\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1721__A1 iram_latched\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3267_ _0048_ clknet_leaf_30_user_clock2 iram_latched\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3198_ net235 _1499_ _1505_ _0761_ _0378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2218_ _0813_ net455 _0794_ _0089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2149_ clk_div.next_div_buff\[2\] _0765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1598__I _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output185_I net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2588__I0 wb_compressor.wb_i_dat\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2201__A2 _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3334__CLK clknet_4_4_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1960__B2 _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire234_I _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2268__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2825__C _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2440__A2 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1951__A1 _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3121_ sspi.res_data\[4\] net259 _1282_ sspi.res_data\[5\] _1459_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3052_ sspi.req_data\[10\] m_arbiter.wb0_o_dat\[10\] _1401_ _1413_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_40_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2259__A2 _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2003_ wb_compressor.state\[6\] wb_compressor.state\[2\] _0555_ _0666_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3208__A1 _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2905_ _0619_ _0636_ _1275_ _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_45_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2836_ sspi.res_data\[12\] _1227_ _1252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2767_ sspi.bit_cnt\[1\] net204 _1199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2698_ _0774_ _1139_ _0244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1718_ _1559_ _1562_ _1565_ _1568_ _0424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
X_1649_ net90 _1566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3319_ _0099_ clknet_4_8_0_net196 wb_cross_clk.m_s_sync.d_data\[27\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2926__B _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2645__C _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2670__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2725__A3 _1160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2413__A2 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3159__S _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2964__A3 _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2621_ wb_compressor.state\[6\] _0531_ _0575_ _1070_ _1023_ _1071_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_35_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput116 net116 inner_wb_i_dat[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput105 net105 inner_disable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_51_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2552_ _1554_ _0933_ _1028_ _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_23_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput138 net138 iram_i_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput149 net149 iram_i_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput127 net127 iram_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_11_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2483_ wb_cross_clk.s_m_sync.s_xfer_xor_flag _0676_ _0980_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3104_ clk_div.cnt\[13\] _1444_ _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3035_ _1404_ _0316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinterconnect_outer_273 la_data_out[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_284 la_data_out[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_295 la_data_out[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_53_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2404__A2 _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2819_ _1239_ _1240_ _0264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2701__S _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input61_I iram_o_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output148_I net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2375__C _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3522__CLK clknet_leaf_16_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput18 inner_wb_adr[23] net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput29 inner_wb_o_dat[10] net29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_20_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2954__I0 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1906__A1 _0525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_net196_I net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1983_ _0652_ net140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_55_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2604_ _0641_ net91 _1060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3584_ _0349_ clknet_leaf_7_user_clock2 m_arbiter.wb0_adr\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2535_ wb_compressor.wb_ack wb_compressor.wb_err _1002_ _1018_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2466_ _0971_ _0180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2397_ _0933_ _0934_ _0935_ _0147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3018_ _1390_ _1392_ _1335_ _0311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2625__A2 _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1903__A4 _0409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2320_ _0879_ _0885_ _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2552__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2251_ _0836_ net463 _0817_ _0099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_42_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_42_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2855__A2 _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2182_ _0788_ net433 _0544_ _0078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2743__C _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1966_ sspi.state\[2\] _0599_ _0644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2791__A1 _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1897_ _0581_ sspi.sy_clk\[3\] _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_12_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3567_ _0332_ clknet_leaf_41_user_clock2 clk_div.cnt\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3146__I _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ _0933_ net240 _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3498_ _0263_ clknet_leaf_26_user_clock2 sspi.res_data\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2449_ _0962_ _0172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input24_I inner_wb_adr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2846__A2 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2426__S _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2653__C _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3023__A2 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2782__A1 _0609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2782__B2 _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_4_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2534__A1 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2828__C _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold7 net527 net394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_58_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ net162 net225 net221 net186 _0512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1751_ _0428_ wb_compressor.wb_i_dat\[9\] _0412_ _0450_ _0451_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3167__S _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1682_ _1574_ _1575_ _1583_ _1584_ _0390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3421_ _0201_ clknet_4_0_0_net196 wb_cross_clk.s_burst_cnt\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3352_ _0132_ clknet_leaf_26_user_clock2 wb_cross_clk.m_wb_i_dat\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1923__B sspi.bit_cnt\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2303_ net468 _0852_ _0873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2738__C _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3283_ _0064_ clknet_leaf_43_user_clock2 clk_div.next_div_buff\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2828__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2234_ _0824_ net423 _0817_ _0094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1642__C _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2165_ net412 _0777_ _0778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2096_ _0699_ iram_latched\[11\] _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3005__A2 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2998_ _1375_ _1376_ _1377_ sspi.req_addr\[16\] _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1949_ _0579_ _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3619_ _0384_ clknet_leaf_27_user_clock2 net197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2929__B _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output130_I net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3263__CLK clknet_leaf_31_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2755__A1 sspi.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2507__A1 _0933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1730__A2 _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2921_ _1261_ _1316_ sspi.req_data\[14\] _1319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1797__A2 _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2852_ _1260_ _1262_ _1263_ _0274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1803_ wb_compressor.wb_i_dat\[3\] wb_cross_clk.m_wb_i_dat\[3\] _0458_ _0497_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2783_ _1208_ net204 _1211_ _1212_ _1213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_22_Right_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_1734_ wb_cross_clk.m_wb_i_dat\[12\] _0437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1665_ m_arbiter.wb0_adr\[10\] net4 _1557_ _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3404_ _0184_ clknet_leaf_47_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[42\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3335_ _0115_ clknet_4_4_0_net196 wb_cross_clk.m_s_sync.d_data\[43\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_37_Left_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1721__A2 _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3266_ _0047_ clknet_leaf_30_user_clock2 iram_latched\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_31_Right_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2217_ net454 _0800_ _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3197_ net172 _1498_ _1505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_4_10_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2148_ _0762_ _0759_ _0764_ _0069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2079_ _0713_ _0714_ _0631_ _0050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_46_Left_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2985__A1 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input91_I m_io_in[34] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2588__I1 net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2737__A1 net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output178_I net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_64_Left_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3217__A2 _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2841__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2728__A1 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3153__A1 sspi.req_addr\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3120_ _1202_ _1456_ _1457_ _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1703__A2 net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3051_ _1412_ _0324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2002_ _0575_ _0662_ _0665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3208__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2904_ _0634_ _1305_ _0284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2835_ net114 _1251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2719__A1 _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2766_ _1196_ _1198_ _0253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2697_ net184 _1084_ net502 _1139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1717_ _1573_ _1576_ _1580_ _1585_ _0423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
X_1648_ _1563_ _1564_ _1565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_67_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3318_ _0098_ clknet_4_10_0_net196 wb_cross_clk.m_s_sync.d_data\[26\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3249_ _0030_ clknet_4_15_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2958__A1 _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2661__C _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3301__CLK clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2186__A2 _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3135__A1 _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3064__I net244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3013__B _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2949__A1 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1621__A1 _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2620_ _1026_ _1070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2143__I _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput106 net106 inner_embed_mode vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2177__A2 _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2551_ wb_cross_clk.m_s_sync.d_data\[5\] _0458_ _1028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3175__S _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput117 net117 inner_wb_i_dat[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput139 net139 iram_i_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_50_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput128 net128 iram_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2482_ _0979_ _0188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3103_ _1444_ _1445_ _0343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3034_ sspi.req_data\[1\] m_arbiter.wb0_o_dat\[1\] _1402_ _1404_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinterconnect_outer_274 la_data_out[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_285 la_data_out[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_296 la_data_out[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3324__CLK clknet_4_8_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1612__A1 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3474__CLK clknet_4_3_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2818_ sspi.res_data\[6\] _1224_ _0763_ _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2168__A2 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2749_ net254 _1182_ _1183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input54_I iram_o_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3117__A1 _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2937__B net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2715__I1 net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2340__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1603__A1 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput19 inner_wb_adr[2] net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2159__A2 _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1906__A2 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3108__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_41_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_41_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1751__B _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1842__A1 wb_compressor.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1982_ m_arbiter.wb0_o_dat\[15\] net34 _1540_ _0652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2398__A2 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2603_ _1059_ _0229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3583_ _0348_ clknet_leaf_2_user_clock2 net195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2534_ _0543_ _1016_ _1017_ _0202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_2_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2465_ wb_cross_clk.m_s_sync.s_data_ff\[38\] _1574_ _0964_ _0971_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2396_ wb_cross_clk.m_s_sync.s_data_ff\[5\] _0925_ _0935_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2322__A2 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3017_ _1284_ _1391_ sspi.req_addr\[21\] _1392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1833__A1 _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2561__A2 _1027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2077__A1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1746__B _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2552__A2 _0933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2250_ net462 _0829_ _0837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2181_ net432 _0777_ _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2068__A1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1815__A1 _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__I1 net13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1965_ _0641_ _0639_ _0643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1896_ sspi.sy_clk\[2\] _0581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_12_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3566_ _0331_ clknet_leaf_41_user_clock2 clk_div.cnt\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3497_ _0262_ clknet_leaf_22_user_clock2 sspi.res_data\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2543__A2 _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2517_ wb_compressor.wb_ack wb_compressor.wb_err wb_cross_clk.s_burst_cnt\[3\] _1002_
+ _1003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2448_ wb_cross_clk.m_s_sync.s_data_ff\[30\] _0396_ _0949_ _0962_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2379_ net209 _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_input17_I inner_wb_adr[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2059__A1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3111__B _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1657__I1 net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold8 _0866_ net395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_58_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2844__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1750_ _0449_ _0415_ _0450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_29_Left_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_1681_ _1565_ net132 _1593_ _1594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_52_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3420_ _0200_ clknet_4_0_0_net196 wb_cross_clk.s_burst_cnt\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3351_ _0131_ clknet_leaf_26_user_clock2 wb_cross_clk.m_wb_i_dat\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2302_ wb_cross_clk.m_s_sync.d_data\[44\] _0772_ _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input9_I inner_wb_adr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3282_ _0063_ clknet_leaf_42_user_clock2 clk_div.next_div_buff\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2233_ net422 _0800_ _0825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2164_ _0776_ _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2095_ _0724_ _0725_ _0721_ _0055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2770__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2997_ sspi.bit_cnt\[4\] _1375_ _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1948_ sspi.state\[2\] _0629_ _0582_ _0630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1879_ wb_cross_clk.m_s_sync.d_data\[42\] _1579_ _0558_ _0565_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3618_ _0383_ clknet_leaf_29_user_clock2 net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2996__I _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3549_ _0314_ clknet_leaf_6_user_clock2 m_arbiter.wb0_we vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_36_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output123_I net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3408__CLK clknet_leaf_5_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3558__CLK clknet_leaf_16_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2755__A2 _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2507__A2 _0926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2691__A1 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2920_ _1295_ _1317_ _1318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2146__I _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2851_ sspi.req_data\[0\] _1262_ _0763_ _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1802_ _0492_ _0496_ net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2782_ _0609_ _0606_ _0637_ _0639_ _1188_ _1212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_25_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1733_ _0435_ _0436_ net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1664_ m_arbiter.wb0_adr\[11\] net5 _1557_ _1581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_3403_ _0183_ clknet_2_0__leaf_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[41\]
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3334_ _0114_ clknet_4_4_0_net196 wb_cross_clk.m_s_sync.d_data\[42\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3265_ _0046_ clknet_leaf_30_user_clock2 iram_latched\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2216_ wb_cross_clk.m_s_sync.d_data\[17\] _0806_ _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3196_ net234 _1499_ _1504_ _0761_ _0377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2765__B _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2147_ clk_div.next_div_buff\[1\] _0759_ _0763_ _0764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2078_ _0703_ net59 _0714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1895__I _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_24_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input84_I m_io_in[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2737__A2 _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3380__CLK clknet_leaf_31_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_30_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3153__A2 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3050_ sspi.req_data\[9\] m_arbiter.wb0_o_dat\[9\] _1401_ _1412_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2001_ wb_compressor.state\[5\] wb_compressor.state\[4\] _0533_ _0664_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2664__A1 _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2903_ _1295_ _1303_ _1304_ sspi.req_data\[10\] _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2967__A2 _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2834_ _1249_ _1229_ _1250_ _0917_ _0269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_45_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold114_I _0396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2765_ sspi.bit_cnt\[0\] _1197_ _0641_ _1198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2696_ _1134_ _1135_ _1137_ _1093_ _1138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1716_ _0391_ _1579_ _0390_ _0421_ _0422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__3253__CLK clknet_4_13_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1647_ m_arbiter.wb0_adr\[6\] net23 _1523_ _1564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3317_ _0097_ clknet_4_10_0_net196 wb_cross_clk.m_s_sync.d_data\[25\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_12_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3248_ _0029_ clknet_4_15_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_16_Left_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3179_ m_arbiter.wb0_adr\[21\] sspi.req_addr\[21\] _1399_ _1495_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2655__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2715__S _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output190_I net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2450__S _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_7_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2430__I1 net140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_40_user_clock2 clknet_2_2__leaf_user_clock2 clknet_leaf_40_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2894__A1 sspi.bit_cnt\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2646__A1 net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput107 net537 net391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2550_ _0542_ _0575_ _1026_ _1027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__2421__I1 net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput118 net118 inner_wb_i_dat[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_2_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput129 net129 iram_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2481_ wb_cross_clk.m_s_sync.s_data_ff\[46\] _0525_ _0885_ _0979_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3102_ clk_div.cnt\[12\] _1442_ _0756_ _1445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3033_ _1403_ _0315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinterconnect_outer_275 la_data_out[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_286 la_data_out[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_297 la_data_out[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_58_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2334__I _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2817_ _0480_ _0484_ _1227_ _1239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_42_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2748_ _1180_ _1181_ _1182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2679_ _0774_ _1123_ _0241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input47_I inner_wb_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2628__A1 _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2479__I1 _0391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3299__CLK clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2847__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2867__A1 _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2619__A1 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1981_ _0651_ net139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_55_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1993__I _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2602_ wb_compressor.state\[1\] wb_compressor.state\[6\] _0543_ _1058_ _1059_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_24_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3582_ _0347_ clknet_leaf_5_user_clock2 m_arbiter.i_wb0_cyc vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2533_ wb_cross_clk.s_burst_cnt\[2\] _1007_ _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2464_ _0970_ _0179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2395_ _0885_ _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2086__A2 iram_latched\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3016_ _1326_ net252 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3441__CLK clknet_4_13_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1833__A2 net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2849__A1 sspi.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2239__I _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2077__A2 iram_latched\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3026__A1 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3314__CLK clknet_4_11_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2180_ wb_cross_clk.m_s_sync.d_data\[6\] _0783_ _0788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3464__CLK clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1815__A2 _0507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ _0624_ _0632_ _0642_ _0005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2240__A2 _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1895_ _0579_ _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3565_ _0330_ clknet_leaf_14_user_clock2 m_arbiter.wb0_o_dat\[15\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3496_ _0261_ clknet_leaf_23_user_clock2 sspi.res_data\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2516_ wb_cross_clk.s_burst_cnt\[2\] wb_cross_clk.s_burst_cnt\[1\] wb_cross_clk.s_burst_cnt\[0\]
+ _1002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1751__A1 _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2447_ _0961_ _0171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2378_ wb_cross_clk.m_new_req_flag _0922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2059__A2 _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2231__A2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3337__CLK clknet_4_4_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2678__B _1122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1742__A1 iram_latched\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3487__CLK clknet_leaf_5_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold9 net533 net396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_58_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1680_ net131 _1593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_40_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3350_ _0130_ clknet_leaf_29_user_clock2 wb_cross_clk.m_wb_i_dat\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2301_ _0870_ net479 _0549_ _0115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3281_ _0062_ clknet_leaf_50_user_clock2 clk_div.res_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2232_ wb_cross_clk.m_s_sync.d_data\[22\] _0806_ _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2163_ wb_cross_clk.m_s_sync.d_xfer_xor_sync\[2\] wb_cross_clk.m_s_sync.d_xfer_xor_sync\[1\]
+ _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_2094_ iram_wb_ack net49 _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2996_ _1332_ _1376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2213__A2 _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1947_ _0619_ _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_1878_ wb_cross_clk.m_s_sync.d_data\[38\] _1574_ _0559_ _0564_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3617_ _0382_ clknet_leaf_28_user_clock2 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3548_ _0313_ clknet_leaf_9_user_clock2 sspi.req_addr\[23\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3479_ _0002_ clknet_leaf_5_user_clock2 sspi.state\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_55_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_14_0_net196 clknet_0_net196 clknet_4_14_0_net196 vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__2961__B sspi.req_addr\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2453__S _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2204__A2 _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_30_Left_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1963__A1 _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3502__CLK clknet_leaf_16_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2443__A2 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2850_ _0611_ _1261_ _1262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1801_ _0462_ _0495_ _0496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2781_ _1208_ net243 _1210_ _1211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1732_ iram_latched\[13\] _0426_ _0436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1663_ _1526_ _1577_ _1578_ _1579_ _1580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_0_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3402_ _0182_ clknet_leaf_47_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[40\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3333_ _0113_ clknet_4_6_0_net196 wb_cross_clk.m_s_sync.d_data\[41\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3264_ _0045_ clknet_leaf_30_user_clock2 iram_latched\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_7_Right_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2215_ _0811_ net475 _0794_ _0088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1950__B _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3195_ net171 _1498_ _1504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2146_ _0622_ _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_2077_ _0700_ iram_latched\[5\] _0713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2434__A2 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2979_ _0580_ _1364_ _0300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input77_I m_io_in[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2800__I _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1860__B _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2448__S _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2673__A2 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3525__CLK clknet_leaf_9_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1936__A1 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2000_ _1525_ _0590_ net110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_38_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2664__A2 _1593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2902_ _1208_ _1295_ _1271_ _1304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_46_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2967__A3 _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2833_ sspi.res_data\[11\] _1224_ _1250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2764_ net243 _1188_ _1197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1715_ _1566_ _1570_ _0421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2695_ _0564_ _1078_ _1136_ _1086_ _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1646_ m_arbiter.wb0_adr\[7\] net24 _1557_ _1563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3316_ _0096_ clknet_4_10_0_net196 wb_cross_clk.m_s_sync.d_data\[24\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3548__CLK clknet_leaf_9_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3247_ _0028_ clknet_4_14_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3178_ _1494_ _0369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_65_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2129_ clk_div.next_div_buff\[0\] _0751_ _0752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2407__A2 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output183_I net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1855__B _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2894__A2 _0610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2646__A2 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1810__S _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1909__A1 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput119 net119 inner_wb_i_dat[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput108 net392 net393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2480_ _0978_ _0187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3101_ clk_div.cnt\[12\] _1442_ _1444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3032_ sspi.req_data\[0\] m_arbiter.wb0_o_dat\[0\] _1402_ _1403_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinterconnect_outer_265 irq[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_276 la_data_out[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_287 la_data_out[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_59_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_outer_298 la_data_out[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
X_2816_ _1237_ _1238_ _0263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2747_ sspi.state\[6\] sspi.state\[2\] sspi.state\[4\] _1181_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2678_ net181 _1084_ _1122_ _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1629_ _1547_ _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2325__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2628__A2 _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_2_0_net196 clknet_0_net196 clknet_4_2_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_49_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2461__S _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2564__A1 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1980_ m_arbiter.wb0_o_dat\[14\] net33 _1540_ _0651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3581_ _0346_ clknet_leaf_49_user_clock2 clk_div.cnt\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2601_ wb_compressor.wb_ack _0662_ _0669_ net84 _1058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xrebuffer1 _1522_ net388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2532_ wb_cross_clk.m_s_sync.d_data\[1\] _1004_ _1009_ _1015_ _1016_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_24_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2463_ wb_cross_clk.m_s_sync.s_data_ff\[37\] _1561_ _0964_ _0970_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2394_ _0654_ _0655_ _0933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_48_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3015_ _1348_ _1380_ _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3779_ net250 net167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2849__A2 _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2785__A1 _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2874__B _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1963_ _0641_ sspi.state\[2\] _0620_ _0642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_50_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1894_ _0524_ _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_55_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3564_ _0329_ clknet_leaf_15_user_clock2 m_arbiter.wb0_o_dat\[14\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3495_ _0260_ clknet_leaf_23_user_clock2 sspi.res_data\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2515_ _1001_ _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2446_ wb_cross_clk.m_s_sync.s_data_ff\[29\] _1563_ _0949_ _0961_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2377_ _0414_ _0889_ _0921_ _0917_ _0141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3008__A2 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3192__A1 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1742__A2 _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3183__A1 sspi.req_addr\[23\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1733__A2 _0436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3431__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2300_ net478 _0852_ _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3280_ _0061_ clknet_leaf_33_user_clock2 iram_wb_ack_del vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2930__A1 _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2231_ _0822_ _0771_ _0823_ _0660_ _0093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2162_ wb_cross_clk.m_s_sync.d_data\[1\] _0771_ _0775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2093_ _0699_ iram_latched\[10\] _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3212__C _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2623__I _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2995_ _0611_ _1323_ _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1946_ sspi.state\[6\] _0614_ _0628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1877_ _0560_ _0561_ _0562_ _0563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3616_ _0381_ clknet_leaf_28_user_clock2 net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3547_ _0312_ clknet_leaf_8_user_clock2 sspi.req_addr\[22\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2921__A1 _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3478_ _0014_ clknet_4_3_0_net196 wb_compressor.state\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_2429_ _0952_ _0162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input22_I inner_wb_adr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1702__I net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3304__CLK clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3454__CLK clknet_4_3_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2912__A1 _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1715__A2 _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2979__A1 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ _0493_ _0494_ _0495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2780_ _1200_ net256 _1210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_14_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1731_ _0428_ wb_compressor.wb_i_dat\[13\] _0412_ _0434_ _0435_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_26_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1662_ m_arbiter.wb0_adr\[20\] net15 _1523_ _1579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_3401_ _0181_ clknet_leaf_47_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[39\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2903__A1 _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3332_ _0112_ clknet_4_6_0_net196 wb_cross_clk.m_s_sync.d_data\[40\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3263_ _0044_ clknet_leaf_31_user_clock2 iram_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3194_ _1539_ _1499_ _1503_ _0761_ _0376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_56_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2214_ net474 _0800_ _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2131__A2 _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2145_ clk_div.curr_div\[1\] _0762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_3_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3327__CLK clknet_4_6_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2076_ _0711_ _0712_ _0631_ _0049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1642__A1 _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3477__CLK clknet_4_2_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2978_ _1303_ _1331_ _1363_ sspi.req_addr\[10\] _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1929_ _0600_ _0582_ _0613_ _0614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2198__A2 _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2370__A2 _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2691__C _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2263__I _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_33_Left_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2212__B _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2361__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Left_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold90 _0859_ net477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2901_ _0605_ _0608_ _1270_ _1287_ _1303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_9_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2832_ net113 _1249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2763_ _0602_ net204 _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1927__A2 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1714_ _0405_ _0393_ _0419_ _0420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2694_ wb_cross_clk.m_s_sync.d_data\[14\] net148 _1033_ _1136_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1645_ _1560_ _1561_ _1562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2352__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3315_ _0095_ clknet_4_8_0_net196 wb_cross_clk.m_s_sync.d_data\[23\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3246_ _0027_ clknet_4_12_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3177_ m_arbiter.wb0_adr\[20\] sspi.req_addr\[20\] _1399_ _1494_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_65_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2792__B _1207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2128_ _0750_ _0525_ _0656_ _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_2059_ _0700_ _0457_ _0591_ _0596_ _0701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1615__A1 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output176_I net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2343__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2459__S _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2894__A3 net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1606__A1 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput109 net109 inner_wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3100_ _1442_ _1443_ _0342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3031_ _1397_ _1400_ _1402_ _0314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinterconnect_outer_266 irq[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_277 la_data_out[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_62_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinterconnect_outer_288 la_data_out[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_299 la_data_out[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_58_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3220__C _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2815_ sspi.res_data\[5\] _1224_ _0763_ _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2746_ sspi.state\[0\] _0618_ _1180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3515__CLK clknet_leaf_16_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2677_ _1093_ _1118_ _1121_ _1122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1628_ _1545_ _1546_ _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3229_ _1518_ _1519_ _1520_ _0020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1911__S _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1836__A1 _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2867__A3 _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1678__I1 net21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1620__I _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3538__CLK clknet_leaf_8_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer2 _1522_ net389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3580_ _0345_ clknet_leaf_49_user_clock2 clk_div.cnt\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2600_ _1057_ _0228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2531_ _1002_ _1014_ net240 _1015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2555__A2 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2462_ _0969_ _0178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2393_ _0932_ _0146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1818__A1 iram_latched\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3014_ _1387_ _1388_ _1389_ _0310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1818__B2 _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2491__A1 _0634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2562__S _1027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3778_ net250 net166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2729_ _1554_ net138 _1166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input52_I iram_o_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2310__B _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output139_I net139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1641__S _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1809__A1 _0498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2785__A2 _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_38_Right_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Right_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Right_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1962_ _0622_ _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_1893_ sspi.state\[1\] _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3632_ _0389_ clknet_leaf_4_user_clock2 m_arbiter.o_sel_sig vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3563_ _0328_ clknet_leaf_15_user_clock2 m_arbiter.wb0_o_dat\[13\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3494_ _0259_ clknet_leaf_23_user_clock2 sspi.res_data\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2514_ _0623_ _1000_ _1001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_65_Right_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2445_ _0960_ _0170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2376_ wb_cross_clk.s_m_sync.s_data_ff\[17\] _0888_ _0921_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2700__A2 _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2059__A4 _0596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3192__A2 _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2467__S _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3383__CLK clknet_leaf_31_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2215__B _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3183__A2 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2230_ net485 _0772_ _0823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2885__B _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2161_ _0768_ _0771_ _0773_ _0774_ _0072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2092_ _0722_ _0723_ _0721_ _0054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2994_ _1373_ _1374_ _1335_ _0305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1945_ _0627_ _0009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1876_ wb_cross_clk.m_s_sync.d_data\[37\] net524 _0559_ _0562_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3615_ _0380_ clknet_leaf_25_user_clock2 net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3256__CLK clknet_4_13_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3546_ _0311_ clknet_leaf_7_user_clock2 sspi.req_addr\[21\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1980__I0 m_arbiter.wb0_o_dat\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3477_ _0013_ clknet_4_2_0_net196 wb_compressor.state\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2428_ wb_cross_clk.m_s_sync.s_data_ff\[20\] net139 _0949_ _0952_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2359_ wb_cross_clk.s_m_sync.s_data_ff\[9\] _0891_ _0912_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2685__A1 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I inner_wb_adr[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2676__B2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2676__A1 net220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1651__A2 _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1730_ _0433_ _0415_ _0434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1661_ _1526_ net18 _1578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3400_ _0180_ clknet_leaf_6_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[38\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3331_ _0111_ clknet_4_6_0_net196 wb_cross_clk.m_s_sync.d_data\[39\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3262_ _0043_ clknet_4_13_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[17\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input7_I inner_wb_adr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3193_ net170 _1498_ _1503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2667__A1 _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2213_ wb_cross_clk.m_s_sync.d_data\[16\] _0806_ _0811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2144_ _0758_ _0759_ _0760_ _0761_ _0068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1890__A2 _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2075_ _0703_ net58 _0712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2570__S _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2977_ _1208_ _1271_ _1336_ _1363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1928_ _0606_ _0612_ _0613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_32_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1859_ _0546_ _0547_ _0548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3529_ _0294_ clknet_leaf_9_user_clock2 sspi.req_addr\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2658__A1 wb_cross_clk.m_s_sync.d_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output121_I net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3421__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2897__A1 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1824__S _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold91 wb_cross_clk.m_s_sync.s_data_ff\[43\] net478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold80 _0860_ net467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_58_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2900_ _1300_ _1302_ _1207_ _0283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2831_ _1247_ _1229_ _1248_ _0917_ _0268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_54_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2762_ _0597_ _1189_ _1194_ _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_5_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__I1 net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1713_ _0391_ _1579_ _0419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2693_ wb_cross_clk.m_s_sync.d_data\[30\] _1080_ _0556_ _1135_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3218__C _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1644_ m_arbiter.wb0_adr\[15\] net9 _1522_ _1561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3314_ _0094_ clknet_4_11_0_net196 wb_cross_clk.m_s_sync.d_data\[22\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3245_ _0026_ clknet_4_14_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2629__I _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3176_ _1493_ _0368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3444__CLK clknet_4_5_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2127_ _0469_ _0407_ _0409_ _0749_ _0750_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_49_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2058_ _0699_ _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_49_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2812__A1 sspi.res_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2415__I1 net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input82_I m_io_in[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1644__S _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2475__S _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1618__I _1538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1790__A1 iram_latched\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3317__CLK clknet_4_10_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1790__B2 _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3467__CLK clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3030_ _1401_ _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xinterconnect_outer_267 irq[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_278 la_data_out[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_62_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_outer_289 la_data_out[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_19_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2814_ _0486_ _0490_ _1227_ _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_26_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2022__A2 _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2745_ sspi.state\[1\] _1178_ _1179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2676_ net220 _1079_ _1120_ _1086_ _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1627_ _1524_ m_arbiter.wb0_o_dat\[1\] _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1781__A1 _0460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3228_ _1518_ _1519_ _1520_ _0019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_61_Left_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3159_ m_arbiter.wb0_adr\[11\] sspi.req_addr\[11\] _1478_ _1485_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1836__A2 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2261__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3210__A1 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1772__A1 _0468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3029__A1 sspi.state\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2218__B _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2252__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer3 _0404_ net500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_51_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2888__B _0622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2530_ wb_cross_clk.s_burst_cnt\[1\] wb_cross_clk.s_burst_cnt\[0\] wb_cross_clk.s_burst_cnt\[2\]
+ _1014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2461_ wb_cross_clk.m_s_sync.s_data_ff\[36\] _1560_ _0964_ _0969_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2392_ wb_cross_clk.m_s_sync.s_data_ff\[4\] _0931_ _0923_ _0932_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3013_ _0629_ _1388_ _0622_ _1389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1818__A2 _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2491__A2 _0880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2243__A2 _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3777_ net250 net165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2728_ _1072_ net498 _1165_ _0660_ _0248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_14_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2659_ _1554_ _1539_ _1105_ _1106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input45_I inner_wb_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_45_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1961_ _0634_ _0640_ _0006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2225__A2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1892_ _0576_ _0577_ _0010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ rst_cw_sync.reset_sync_ff\[2\] _0022_ clknet_4_0_0_net196 net193 vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3562_ _0327_ clknet_leaf_23_user_clock2 m_arbiter.wb0_o_dat\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1736__A1 _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2513_ _0926_ _0990_ _0999_ _0885_ _1000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_59_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3493_ _0258_ clknet_leaf_18_user_clock2 sspi.res_data\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2444_ wb_cross_clk.m_s_sync.s_data_ff\[28\] _1564_ _0949_ _0960_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2375_ _0429_ _0889_ _0920_ _0917_ _0140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2637__I _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2216__A2 _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1727__A1 iram_latched\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3528__CLK clknet_leaf_8_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2991__B _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2207__A2 _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_user_clock2_I clknet_2_2__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ _0542_ _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2091_ iram_wb_ack net63 _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2993_ _1218_ _1323_ sspi.req_addr\[15\] _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1944_ _0623_ _0626_ _0627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3614_ _0379_ clknet_leaf_25_user_clock2 net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1875_ wb_cross_clk.m_s_sync.d_data\[35\] net507 _0559_ _0561_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3545_ _0310_ clknet_leaf_4_user_clock2 sspi.req_addr\[20\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3476_ _0012_ clknet_4_2_0_net196 wb_compressor.state\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__2568__S _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2427_ _0951_ _0161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2134__A1 _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2358_ wb_cross_clk.m_wb_i_dat\[7\] _0896_ _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2289_ net407 _0863_ _0846_ _0111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_55_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Left_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3173__I0 m_arbiter.wb0_adr\[18\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2676__A2 _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_21_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ m_arbiter.wb0_adr\[23\] _1577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_1_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3330_ _0110_ clknet_4_7_0_net196 wb_cross_clk.m_s_sync.d_data\[38\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3261_ _0042_ clknet_4_7_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[16\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3192_ _1544_ _1499_ _1502_ _0761_ _0375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2667__A2 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2212_ _0809_ net435 _0794_ _0087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2143_ _0622_ _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_2074_ _0700_ iram_latched\[4\] _0711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2976_ _1361_ _1362_ _1335_ _0299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1927_ _0608_ _0611_ _0612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1858_ net84 wb_compressor.state\[2\] _0547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3373__CLK clknet_leaf_38_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1789_ wb_compressor.wb_i_dat\[5\] wb_cross_clk.m_wb_i_dat\[5\] _0458_ _0485_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3528_ _0293_ clknet_leaf_8_user_clock2 sspi.req_addr\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3459_ _0239_ clknet_4_14_0_net196 net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2658__A2 _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2830__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2897__A2 _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold81 wb_cross_clk.m_s_sync.s_data_ff\[44\] net468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold92 _0871_ net479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold70 _0845_ net457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_58_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3246__CLK clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_4_user_clock2_I clknet_2_0__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2830_ sspi.res_data\[10\] _1224_ _1248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2821__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2761_ net243 _1194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2692_ _1073_ net501 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1712_ net255 net247 _0418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1643_ m_arbiter.wb0_adr\[14\] net8 net389 _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3313_ _0093_ clknet_4_12_0_net196 wb_cross_clk.m_s_sync.d_data\[21\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3244_ net535 clknet_leaf_13_user_clock2 net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3175_ m_arbiter.wb0_adr\[19\] sspi.req_addr\[19\] _1399_ _1493_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_65_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2126_ _1570_ _0394_ net255 _0397_ _0749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_37_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2057_ iram_wb_ack _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__3065__A2 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2812__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2959_ sspi.bit_cnt\[4\] _0611_ _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_8_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input75_I m_io_in[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2500__A1 _0933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3269__CLK clknet_leaf_31_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap208_I _1071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2803__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1790__A2 _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1634__I _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2590__I1 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinterconnect_outer_268 la_data_out[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinterconnect_outer_279 la_data_out[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_62_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2813_ _1235_ _1236_ _0262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2744_ sspi.state\[5\] _0624_ _1178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2675_ _1554_ net235 _1119_ _1120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1626_ _1540_ net35 _1545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1781__A2 _0478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2576__S _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3227_ _1518_ _1519_ _1520_ _0018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3158_ _1484_ _0359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2109_ net54 _0703_ _0735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3089_ _1431_ _1435_ _1432_ _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_9_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3210__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output181_I net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1772__A2 _0403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2572__I1 net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2721__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2994__B _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3029__A2 _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1629__I _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2234__B _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3201__A2 _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Left_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3434__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2460_ _0968_ _0177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1763__A2 _1594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2391_ _1525_ net45 _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__2712__A1 _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_2__f_user_clock2 clknet_0_user_clock2 clknet_2_2__leaf_user_clock2 vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3012_ _1344_ _1380_ _1388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2779__A1 _0610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3776_ net250 net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2727_ net189 _1084_ _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2951__A1 _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2658_ wb_cross_clk.m_s_sync.d_data\[9\] _0428_ _1105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1609_ _1527_ m_arbiter.wb0_o_dat\[5\] _1532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2589_ _1051_ _0223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input38_I inner_wb_o_dat[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3307__CLK clknet_4_11_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1745__A2 _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2170__A2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1960_ sspi.state\[0\] _0620_ _0638_ _0639_ _0640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1891_ wb_compressor.state\[1\] _0542_ _0577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2899__B sspi.req_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3630_ rst_cw_sync.reset_sync_ff\[1\] _0021_ clknet_4_0_0_net196 rst_cw_sync.reset_sync_ff\[2\]
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_0_24_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3561_ _0326_ clknet_leaf_18_user_clock2 m_arbiter.wb0_o_dat\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2512_ wb_cross_clk.m_burst_cnt\[3\] _0998_ _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3492_ _0257_ clknet_leaf_10_user_clock2 sspi.bit_cnt\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_11_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2443_ _0406_ _0925_ _0959_ _0169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2374_ wb_cross_clk.s_m_sync.s_data_ff\[16\] _0888_ _0920_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2161__A2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2139__B _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3110__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2621__B1 _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3759_ clknet_leaf_24_user_clock2 net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1727__A2 _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2152__A2 _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1663__A1 _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2915__A1 _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2231__C _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ _0699_ iram_latched\[9\] _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2992_ _0629_ _0613_ _1336_ _1373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_28_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1943_ _0624_ _0598_ _0625_ _0626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3613_ _0378_ clknet_leaf_27_user_clock2 net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1874_ wb_cross_clk.m_s_sync.d_data\[41\] _1583_ _0559_ _0560_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2906__A1 _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3544_ _0309_ clknet_leaf_7_user_clock2 sspi.req_addr\[19\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3475_ _0001_ clknet_4_3_0_net196 wb_compressor.state\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_24_Left_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_2426_ wb_cross_clk.m_s_sync.s_data_ff\[19\] net138 _0949_ _0951_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2134__A2 _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2357_ _0909_ _0910_ _0895_ _0132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2288_ wb_cross_clk.m_s_sync.d_data\[39\] _0771_ _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2584__S _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1645__A1 _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1948__A2 _0629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2373__A2 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2061__A1 _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1637__I _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2364__A2 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3260_ _0041_ clknet_4_4_0_net196 wb_cross_clk.s_m_sync.s_data_ff\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3191_ net169 _1498_ _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2211_ net434 _0800_ _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2142_ _0737_ _0759_ _0760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2073_ _0709_ _0710_ _0631_ _0048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1627__A1 _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2975_ _1301_ _1351_ sspi.req_addr\[9\] _1362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3518__CLK clknet_leaf_8_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1926_ _0609_ _0610_ net259 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_44_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1650__I1 net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2152__B _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1857_ wb_compressor.l_we _0546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1788_ _0480_ _0484_ net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2355__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3527_ _0292_ clknet_leaf_9_user_clock2 sspi.req_addr\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_770 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3458_ _0238_ clknet_4_14_0_net196 net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3389_ _0169_ clknet_leaf_45_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[27\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2409_ wb_cross_clk.m_s_sync.s_data_ff\[11\] _0937_ _0942_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input20_I inner_wb_adr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_4_5_0_net196 clknet_0_net196 clknet_4_5_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_63_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1658__S _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1641__I1 net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2346__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2897__A3 _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_wire260_I net261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold71 wb_cross_clk.m_s_sync.s_data_ff\[46\] net458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold82 _0873_ net469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold60 _0857_ net447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_26_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold93 wb_cross_clk.m_s_sync.s_data_ff\[2\] net480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1609__A1 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2237__B _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2760_ _0639_ _1192_ _1180_ _1193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1711_ _1554_ wb_compressor.wb_i_dat\[15\] _0413_ _0416_ _0417_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2691_ _1072_ net494 _1133_ _0660_ _0243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_14_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1642_ _1526_ _1555_ _1556_ _1558_ _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__2337__A2 _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2700__B _0556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3312_ _0092_ clknet_4_14_0_net196 wb_cross_clk.m_s_sync.d_data\[20\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3243_ net87 clknet_leaf_13_user_clock2 irq_s_ff\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3174_ _1492_ _0367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_65_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2125_ _0748_ _0062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2056_ _0698_ _0043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2147__B _0763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2958_ _1331_ _1348_ _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1909_ _1553_ net260 _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2889_ _1260_ _1292_ _1293_ _0281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input68_I m_io_in[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2328__A2 _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2016__A1 wb_compressor.wb_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_2_0_net196_I clknet_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinterconnect_outer_269 la_data_out[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_59_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2682__S _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2812_ sspi.res_data\[4\] _1224_ _0763_ _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2558__A2 _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2743_ _1072_ net215 _1177_ _0660_ _0251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_41_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ wb_cross_clk.m_s_sync.d_data\[11\] _0428_ _1119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1625_ _1544_ net142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_10_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2730__A2 _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1761__S _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3226_ _1518_ _1519_ _1520_ _0017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3157_ m_arbiter.wb0_adr\[10\] sspi.req_addr\[10\] _1478_ _1484_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2108_ iram_latched\[15\] _0700_ _0734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3088_ clk_div.cnt\[8\] _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2039_ wb_compressor.wb_i_dat\[7\] wb_cross_clk.s_m_sync.s_data_ff\[9\] _0688_ _0690_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2797__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3236__CLK clknet_4_0_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2721__A2 net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3628__264 net264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_28_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2390_ _0930_ _0145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3011_ sspi.req_addr\[20\] _1387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2779__A2 net259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_29_user_clock2_I clknet_2_3__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2144__C _0761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3259__CLK clknet_4_5_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3775_ net250 net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2726_ _0565_ _1079_ net497 _1164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2657_ wb_cross_clk.m_s_sync.d_data\[25\] _1080_ _0556_ _1104_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1608_ net236 net146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2588_ wb_compressor.wb_i_dat\[11\] net79 net212 _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3770__I net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3209_ net194 _1508_ _1512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2335__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__S _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3195__A2 _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2070__B _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2458__A1 _0468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Right_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1681__A2 net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1890_ wb_compressor.state\[0\] _0575_ _0576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2481__I1 _0525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3560_ _0325_ clknet_leaf_18_user_clock2 m_arbiter.wb0_o_dat\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_25_Right_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2933__A2 _0611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2511_ wb_cross_clk.m_burst_cnt\[2\] _0992_ _0998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3491_ _0256_ clknet_leaf_10_user_clock2 sspi.bit_cnt\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_2442_ wb_cross_clk.m_s_sync.s_data_ff\[27\] _0923_ _0959_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2373_ _0433_ _0889_ _0919_ _0917_ _0139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2697__A1 net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_user_clock2_I clknet_2_1__leaf_user_clock2 vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_34_Right_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_49_Left_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2621__A1 wb_compressor.state\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3765__I net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_43_Right_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3758_ clknet_leaf_13_user_clock2 net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2924__A2 _1295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2709_ _0566_ _1078_ _1148_ _1086_ _1149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_30_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input50_I iram_o_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Left_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Right_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output137_I net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3424__CLK clknet_4_1_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Left_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Right_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2612__A1 net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2679__A1 _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2991_ _1371_ _1372_ _1335_ _0304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1942_ sspi.state\[7\] _0614_ _0625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1957__A3 _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1873_ _0558_ _0559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_28_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3612_ _0377_ clknet_leaf_27_user_clock2 net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2906__A2 _1294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3543_ _0308_ clknet_leaf_4_user_clock2 sspi.req_addr\[18\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3237__D net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3474_ _0011_ clknet_4_3_0_net196 wb_compressor.state\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_2425_ _0950_ _0160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2356_ wb_cross_clk.s_m_sync.s_data_ff\[8\] _0891_ _0910_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3447__CLK clknet_4_12_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2287_ net406 _0776_ _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input98_I mgt_wb_rst_i vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1948__A3 _0582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2436__I1 net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2061__A2 iram_latched\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3010__A1 _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2210_ wb_cross_clk.m_s_sync.d_data\[15\] _0806_ _0809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3190_ _1548_ _1499_ _1501_ _0761_ _0374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_56_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2141_ clk_div.next_div_val _0747_ _0759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2072_ _0703_ net57 _0710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2974_ _0619_ _0636_ _1266_ _1336_ _1361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_60_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1925_ sspi.bit_cnt\[2\] _0610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_44_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold128_I _1581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1856_ _0533_ _0540_ wb_compressor.state\[5\] _0545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1787_ _0462_ _0483_ _0484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3526_ _0291_ clknet_leaf_9_user_clock2 sspi.req_addr\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3457_ _0237_ clknet_4_9_0_net196 net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2408_ net234 _0934_ _0941_ _0152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3388_ _0168_ clknet_leaf_35_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[26\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2339_ _0897_ _0898_ _0895_ _0126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_2_Right_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I inner_wb_adr[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2815__A1 sspi.res_data\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2291__A2 _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold50 _0853_ net437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold72 _0877_ net459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold83 wb_cross_clk.m_s_sync.s_data_ff\[45\] net470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold61 wb_cross_clk.m_s_sync.s_data_ff\[33\] net448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold94 _0779_ net481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_58_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2282__A2 _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1710_ _0414_ _0415_ _0416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2690_ net183 _1084_ _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1641_ m_arbiter.wb0_adr\[9\] net26 _1557_ _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XANTENNA__3292__CLK clknet_4_1_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3311_ _0091_ clknet_4_14_0_net196 wb_cross_clk.m_s_sync.d_data\[19\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3242_ net532 clknet_leaf_0_user_clock2 clk_div.clock_sel vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input5_I inner_wb_adr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3173_ m_arbiter.wb0_adr\[18\] sspi.req_addr\[18\] _1399_ _1492_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2124_ clk_div.res_clk net244 _0748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_37_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2055_ wb_compressor.wb_i_dat\[15\] wb_cross_clk.s_m_sync.s_data_ff\[17\] _0688_
+ _0698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2273__A2 _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2957_ _1284_ _1332_ _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2888_ sspi.req_data\[7\] _1292_ _0622_ _1293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1908_ wb_cross_clk.msy_xor_ack wb_cross_clk.prev_xor_ack _0593_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_60_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1839_ _0528_ wb_cross_clk.m_s_sync.d_data\[46\] net490 _0529_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__3773__I net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3509_ _0274_ clknet_leaf_13_user_clock2 sspi.req_data\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2073__B _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2016__A2 wb_compressor.wb_err vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1775__A1 _0405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2255__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2811_ _0492_ _0496_ _1227_ _1235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_42_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2742_ net192 _1093_ _1177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1766__A1 net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2673_ wb_cross_clk.m_s_sync.d_data\[27\] _1080_ _0555_ _1117_ _1118_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1624_ _1543_ _1544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3225_ _1518_ _1519_ _1520_ _0016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3034__S _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3156_ _1483_ _0358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2107_ _0732_ _0733_ _0721_ _0059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3087_ _1419_ _1433_ _1434_ _0338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2038_ _0689_ _0034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3768__I net249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2246__A2 _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input80_I m_io_in[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1757__A1 iram_latched\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_max_cap213_I net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2485__A2 _0623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3330__CLK clknet_4_7_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3010_ _0988_ _1385_ _1386_ _0309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_47_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2228__A2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1987__A1 _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3774_ net249 net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2725_ _1158_ _1159_ _1160_ _1161_ _1162_ _1163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_14_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2656_ _1073_ net528 _1103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1607_ _1525_ net40 _1530_ _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2587_ _1050_ _0222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3208_ _1548_ _1509_ _1511_ _1253_ _0382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3139_ _1474_ _0350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2219__A2 _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2351__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2458__A2 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2526__B _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1681__A3 _1593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3490_ _0255_ clknet_leaf_12_user_clock2 sspi.bit_cnt\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_12_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2510_ _0997_ _0198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2441_ _1593_ _0925_ _0958_ _0168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2688__S _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2372_ wb_cross_clk.s_m_sync.s_data_ff\[15\] _0888_ _0919_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2697__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3376__CLK clknet_leaf_31_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2385__A1 _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2708_ wb_cross_clk.m_s_sync.d_data\[16\] net135 _0559_ _1148_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2639_ wb_cross_clk.m_s_sync.d_data\[23\] _0458_ _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input43_I inner_wb_o_dat[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3249__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2990_ _1316_ _1351_ sspi.req_addr\[14\] _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1941_ sspi.state\[3\] _0624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1872_ net490 _0558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_3611_ _0376_ clknet_leaf_28_user_clock2 net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2703__C _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2906__A3 _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3542_ _0307_ clknet_leaf_8_user_clock2 sspi.req_addr\[17\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3473_ _0000_ clknet_4_2_0_net196 wb_compressor.state\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2424_ wb_cross_clk.m_s_sync.s_data_ff\[18\] net137 _0949_ _0950_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2355_ wb_cross_clk.m_wb_i_dat\[6\] _0896_ _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2286_ net467 _0861_ _0846_ _0110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3042__S _1402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2166__B _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3776__I net250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_7_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2833__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3541__CLK clknet_leaf_9_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2076__B _0631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2140_ clk_div.next_div_buff\[0\] _0758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2071_ _0700_ iram_latched\[3\] _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_19_user_clock2 clknet_2_1__leaf_user_clock2 clknet_leaf_19_user_clock2
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2824__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2973_ _0988_ _1359_ _1360_ _0298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2714__B _0555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_1924_ sspi.bit_cnt\[3\] _0609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_44_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_1855_ _0532_ _0541_ _0544_ _0014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1786_ _0481_ _0482_ _0483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3525_ _0290_ clknet_leaf_9_user_clock2 sspi.req_addr\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2760__A1 _0639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3456_ _0236_ clknet_4_9_0_net196 net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2407_ wb_cross_clk.m_s_sync.s_data_ff\[10\] _0937_ _0941_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3387_ _0167_ clknet_leaf_38_user_clock2 wb_cross_clk.m_s_sync.s_data_ff\[25\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2338_ wb_cross_clk.s_m_sync.s_data_ff\[2\] _0891_ _0898_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2269_ net448 _0829_ _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2815__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2051__I0 wb_compressor.wb_i_dat\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2751__A1 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1690__S _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold40 _0782_ net427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold73 wb_cross_clk.m_s_sync.s_data_ff\[42\] net460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold51 wb_cross_clk.m_s_sync.s_data_ff\[35\] net438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold62 _0850_ net449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold95 net514 net482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold84 _0875_ net471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_58_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2806__A2 _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold99_I inner_wb_8_burst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2026__S _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2114__S0 _0737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3437__CLK clknet_4_15_0_net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1640_ _1522_ _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2742__A1 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3310_ _0090_ clknet_4_11_0_net196 wb_cross_clk.m_s_sync.d_data\[18\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3587__CLK clknet_leaf_8_user_clock2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3241_ net88 clknet_leaf_0_user_clock2 split_s_ff\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3172_ _1491_ _0366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2123_ _0739_ _0742_ _0744_ _0746_ _0747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_37_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_2054_ _0697_ _0042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_17_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2956_ _1347_ _0294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2887_ _0606_ _0636_ _1261_ _1292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_45_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1907_ iram_wb_ack_del net229 _0591_ _0462_ _0588_ _0592_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__1784__A2 _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1838_ wb_cross_clk.ack_next_hold _0528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1769_ _1526_ m_arbiter.wb0_adr\[12\] _0467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2733__A1 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3508_ _0273_ clknet_leaf_18_user_clock2 sspi.res_data\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3439_ _0219_ clknet_4_13_0_net196 wb_compressor.wb_i_dat\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2354__B _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3213__A2 _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2972__A1 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2529__B _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3204__I _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3140__S _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2264__B _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_2810_ _1233_ _1234_ _0261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_42_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2741_ _0556_ _0562_ _0567_ _1079_ _1175_ _1176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_54_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2672_ _1033_ _0406_ _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1623_ _1541_ _1542_ _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2191__A2 _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3224_ _1518_ _1519_ _1520_ _0015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
.ends

