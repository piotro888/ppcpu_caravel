magic
tech gf180mcuD
magscale 1 5
timestamp 1699380672
<< obsm1 >>
rect 672 911 119280 33585
<< metal2 >>
rect 3024 34600 3080 35000
rect 3920 34600 3976 35000
rect 4816 34600 4872 35000
rect 5712 34600 5768 35000
rect 6608 34600 6664 35000
rect 7504 34600 7560 35000
rect 8400 34600 8456 35000
rect 9296 34600 9352 35000
rect 10192 34600 10248 35000
rect 11088 34600 11144 35000
rect 11984 34600 12040 35000
rect 12880 34600 12936 35000
rect 13776 34600 13832 35000
rect 14672 34600 14728 35000
rect 15568 34600 15624 35000
rect 16464 34600 16520 35000
rect 17360 34600 17416 35000
rect 18256 34600 18312 35000
rect 19152 34600 19208 35000
rect 20048 34600 20104 35000
rect 20944 34600 21000 35000
rect 21840 34600 21896 35000
rect 22736 34600 22792 35000
rect 23632 34600 23688 35000
rect 24528 34600 24584 35000
rect 25424 34600 25480 35000
rect 26320 34600 26376 35000
rect 27216 34600 27272 35000
rect 28112 34600 28168 35000
rect 29008 34600 29064 35000
rect 29904 34600 29960 35000
rect 30800 34600 30856 35000
rect 31696 34600 31752 35000
rect 32592 34600 32648 35000
rect 33488 34600 33544 35000
rect 34384 34600 34440 35000
rect 35280 34600 35336 35000
rect 36176 34600 36232 35000
rect 37072 34600 37128 35000
rect 37968 34600 38024 35000
rect 38864 34600 38920 35000
rect 39760 34600 39816 35000
rect 40656 34600 40712 35000
rect 41552 34600 41608 35000
rect 42448 34600 42504 35000
rect 43344 34600 43400 35000
rect 44240 34600 44296 35000
rect 45136 34600 45192 35000
rect 46032 34600 46088 35000
rect 46928 34600 46984 35000
rect 47824 34600 47880 35000
rect 48720 34600 48776 35000
rect 49616 34600 49672 35000
rect 50512 34600 50568 35000
rect 51408 34600 51464 35000
rect 52304 34600 52360 35000
rect 53200 34600 53256 35000
rect 54096 34600 54152 35000
rect 54992 34600 55048 35000
rect 55888 34600 55944 35000
rect 56784 34600 56840 35000
rect 57680 34600 57736 35000
rect 58576 34600 58632 35000
rect 59472 34600 59528 35000
rect 60368 34600 60424 35000
rect 61264 34600 61320 35000
rect 62160 34600 62216 35000
rect 63056 34600 63112 35000
rect 63952 34600 64008 35000
rect 64848 34600 64904 35000
rect 65744 34600 65800 35000
rect 66640 34600 66696 35000
rect 67536 34600 67592 35000
rect 68432 34600 68488 35000
rect 69328 34600 69384 35000
rect 70224 34600 70280 35000
rect 71120 34600 71176 35000
rect 72016 34600 72072 35000
rect 72912 34600 72968 35000
rect 73808 34600 73864 35000
rect 74704 34600 74760 35000
rect 75600 34600 75656 35000
rect 76496 34600 76552 35000
rect 77392 34600 77448 35000
rect 78288 34600 78344 35000
rect 79184 34600 79240 35000
rect 80080 34600 80136 35000
rect 80976 34600 81032 35000
rect 81872 34600 81928 35000
rect 82768 34600 82824 35000
rect 83664 34600 83720 35000
rect 84560 34600 84616 35000
rect 85456 34600 85512 35000
rect 86352 34600 86408 35000
rect 87248 34600 87304 35000
rect 88144 34600 88200 35000
rect 89040 34600 89096 35000
rect 89936 34600 89992 35000
rect 90832 34600 90888 35000
rect 91728 34600 91784 35000
rect 92624 34600 92680 35000
rect 93520 34600 93576 35000
rect 94416 34600 94472 35000
rect 95312 34600 95368 35000
rect 96208 34600 96264 35000
rect 97104 34600 97160 35000
rect 98000 34600 98056 35000
rect 98896 34600 98952 35000
rect 99792 34600 99848 35000
rect 100688 34600 100744 35000
rect 101584 34600 101640 35000
rect 102480 34600 102536 35000
rect 103376 34600 103432 35000
rect 104272 34600 104328 35000
rect 105168 34600 105224 35000
rect 106064 34600 106120 35000
rect 106960 34600 107016 35000
rect 107856 34600 107912 35000
rect 108752 34600 108808 35000
rect 109648 34600 109704 35000
rect 110544 34600 110600 35000
rect 111440 34600 111496 35000
rect 112336 34600 112392 35000
rect 113232 34600 113288 35000
rect 114128 34600 114184 35000
rect 115024 34600 115080 35000
rect 115920 34600 115976 35000
rect 116816 34600 116872 35000
rect 4928 0 4984 400
rect 5152 0 5208 400
rect 5376 0 5432 400
rect 5600 0 5656 400
rect 5824 0 5880 400
rect 6048 0 6104 400
rect 6272 0 6328 400
rect 6496 0 6552 400
rect 6720 0 6776 400
rect 6944 0 7000 400
rect 7168 0 7224 400
rect 7392 0 7448 400
rect 7616 0 7672 400
rect 7840 0 7896 400
rect 8064 0 8120 400
rect 8288 0 8344 400
rect 8512 0 8568 400
rect 8736 0 8792 400
rect 8960 0 9016 400
rect 9184 0 9240 400
rect 9408 0 9464 400
rect 9632 0 9688 400
rect 9856 0 9912 400
rect 10080 0 10136 400
rect 10304 0 10360 400
rect 10528 0 10584 400
rect 10752 0 10808 400
rect 10976 0 11032 400
rect 11200 0 11256 400
rect 11424 0 11480 400
rect 11648 0 11704 400
rect 11872 0 11928 400
rect 12096 0 12152 400
rect 12320 0 12376 400
rect 12544 0 12600 400
rect 12768 0 12824 400
rect 12992 0 13048 400
rect 13216 0 13272 400
rect 13440 0 13496 400
rect 13664 0 13720 400
rect 13888 0 13944 400
rect 14112 0 14168 400
rect 14336 0 14392 400
rect 14560 0 14616 400
rect 14784 0 14840 400
rect 15008 0 15064 400
rect 15232 0 15288 400
rect 15456 0 15512 400
rect 15680 0 15736 400
rect 15904 0 15960 400
rect 16128 0 16184 400
rect 16352 0 16408 400
rect 16576 0 16632 400
rect 16800 0 16856 400
rect 17024 0 17080 400
rect 17248 0 17304 400
rect 17472 0 17528 400
rect 17696 0 17752 400
rect 17920 0 17976 400
rect 18144 0 18200 400
rect 18368 0 18424 400
rect 18592 0 18648 400
rect 18816 0 18872 400
rect 19040 0 19096 400
rect 19264 0 19320 400
rect 19488 0 19544 400
rect 19712 0 19768 400
rect 19936 0 19992 400
rect 20160 0 20216 400
rect 20384 0 20440 400
rect 20608 0 20664 400
rect 20832 0 20888 400
rect 21056 0 21112 400
rect 21280 0 21336 400
rect 21504 0 21560 400
rect 21728 0 21784 400
rect 21952 0 22008 400
rect 22176 0 22232 400
rect 22400 0 22456 400
rect 22624 0 22680 400
rect 22848 0 22904 400
rect 23072 0 23128 400
rect 23296 0 23352 400
rect 23520 0 23576 400
rect 23744 0 23800 400
rect 23968 0 24024 400
rect 24192 0 24248 400
rect 24416 0 24472 400
rect 24640 0 24696 400
rect 24864 0 24920 400
rect 25088 0 25144 400
rect 25312 0 25368 400
rect 25536 0 25592 400
rect 25760 0 25816 400
rect 25984 0 26040 400
rect 26208 0 26264 400
rect 26432 0 26488 400
rect 26656 0 26712 400
rect 26880 0 26936 400
rect 27104 0 27160 400
rect 27328 0 27384 400
rect 27552 0 27608 400
rect 27776 0 27832 400
rect 28000 0 28056 400
rect 28224 0 28280 400
rect 28448 0 28504 400
rect 28672 0 28728 400
rect 28896 0 28952 400
rect 29120 0 29176 400
rect 29344 0 29400 400
rect 29568 0 29624 400
rect 29792 0 29848 400
rect 30016 0 30072 400
rect 30240 0 30296 400
rect 30464 0 30520 400
rect 30688 0 30744 400
rect 30912 0 30968 400
rect 31136 0 31192 400
rect 31360 0 31416 400
rect 31584 0 31640 400
rect 31808 0 31864 400
rect 32032 0 32088 400
rect 32256 0 32312 400
rect 32480 0 32536 400
rect 32704 0 32760 400
rect 32928 0 32984 400
rect 33152 0 33208 400
rect 33376 0 33432 400
rect 33600 0 33656 400
rect 33824 0 33880 400
rect 34048 0 34104 400
rect 34272 0 34328 400
rect 34496 0 34552 400
rect 34720 0 34776 400
rect 34944 0 35000 400
rect 35168 0 35224 400
rect 35392 0 35448 400
rect 35616 0 35672 400
rect 35840 0 35896 400
rect 36064 0 36120 400
rect 36288 0 36344 400
rect 36512 0 36568 400
rect 36736 0 36792 400
rect 36960 0 37016 400
rect 37184 0 37240 400
rect 37408 0 37464 400
rect 37632 0 37688 400
rect 37856 0 37912 400
rect 38080 0 38136 400
rect 38304 0 38360 400
rect 38528 0 38584 400
rect 38752 0 38808 400
rect 38976 0 39032 400
rect 39200 0 39256 400
rect 39424 0 39480 400
rect 39648 0 39704 400
rect 39872 0 39928 400
rect 40096 0 40152 400
rect 40320 0 40376 400
rect 40544 0 40600 400
rect 40768 0 40824 400
rect 40992 0 41048 400
rect 41216 0 41272 400
rect 41440 0 41496 400
rect 41664 0 41720 400
rect 41888 0 41944 400
rect 42112 0 42168 400
rect 42336 0 42392 400
rect 42560 0 42616 400
rect 42784 0 42840 400
rect 43008 0 43064 400
rect 43232 0 43288 400
rect 43456 0 43512 400
rect 43680 0 43736 400
rect 43904 0 43960 400
rect 44128 0 44184 400
rect 44352 0 44408 400
rect 44576 0 44632 400
rect 44800 0 44856 400
rect 45024 0 45080 400
rect 45248 0 45304 400
rect 45472 0 45528 400
rect 45696 0 45752 400
rect 45920 0 45976 400
rect 46144 0 46200 400
rect 46368 0 46424 400
rect 46592 0 46648 400
rect 46816 0 46872 400
rect 47040 0 47096 400
rect 47264 0 47320 400
rect 47488 0 47544 400
rect 47712 0 47768 400
rect 47936 0 47992 400
rect 48160 0 48216 400
rect 48384 0 48440 400
rect 48608 0 48664 400
rect 48832 0 48888 400
rect 49056 0 49112 400
rect 49280 0 49336 400
rect 49504 0 49560 400
rect 49728 0 49784 400
rect 49952 0 50008 400
rect 50176 0 50232 400
rect 50400 0 50456 400
rect 50624 0 50680 400
rect 50848 0 50904 400
rect 51072 0 51128 400
rect 51296 0 51352 400
rect 51520 0 51576 400
rect 51744 0 51800 400
rect 51968 0 52024 400
rect 52192 0 52248 400
rect 52416 0 52472 400
rect 52640 0 52696 400
rect 52864 0 52920 400
rect 53088 0 53144 400
rect 53312 0 53368 400
rect 53536 0 53592 400
rect 53760 0 53816 400
rect 53984 0 54040 400
rect 54208 0 54264 400
rect 54432 0 54488 400
rect 54656 0 54712 400
rect 54880 0 54936 400
rect 55104 0 55160 400
rect 55328 0 55384 400
rect 55552 0 55608 400
rect 55776 0 55832 400
rect 56000 0 56056 400
rect 56224 0 56280 400
rect 56448 0 56504 400
rect 56672 0 56728 400
rect 56896 0 56952 400
rect 57120 0 57176 400
rect 57344 0 57400 400
rect 57568 0 57624 400
rect 57792 0 57848 400
rect 58016 0 58072 400
rect 58240 0 58296 400
rect 58464 0 58520 400
rect 58688 0 58744 400
rect 58912 0 58968 400
rect 59136 0 59192 400
rect 59360 0 59416 400
rect 59584 0 59640 400
rect 59808 0 59864 400
rect 60032 0 60088 400
rect 60256 0 60312 400
rect 60480 0 60536 400
rect 60704 0 60760 400
rect 60928 0 60984 400
rect 61152 0 61208 400
rect 61376 0 61432 400
rect 61600 0 61656 400
rect 61824 0 61880 400
rect 62048 0 62104 400
rect 62272 0 62328 400
rect 62496 0 62552 400
rect 62720 0 62776 400
rect 62944 0 63000 400
rect 63168 0 63224 400
rect 63392 0 63448 400
rect 63616 0 63672 400
rect 63840 0 63896 400
rect 64064 0 64120 400
rect 64288 0 64344 400
rect 64512 0 64568 400
rect 64736 0 64792 400
rect 64960 0 65016 400
rect 65184 0 65240 400
rect 65408 0 65464 400
rect 65632 0 65688 400
rect 65856 0 65912 400
rect 66080 0 66136 400
rect 66304 0 66360 400
rect 66528 0 66584 400
rect 66752 0 66808 400
rect 66976 0 67032 400
rect 67200 0 67256 400
rect 67424 0 67480 400
rect 67648 0 67704 400
rect 67872 0 67928 400
rect 68096 0 68152 400
rect 68320 0 68376 400
rect 68544 0 68600 400
rect 68768 0 68824 400
rect 68992 0 69048 400
rect 69216 0 69272 400
rect 69440 0 69496 400
rect 69664 0 69720 400
rect 69888 0 69944 400
rect 70112 0 70168 400
rect 70336 0 70392 400
rect 70560 0 70616 400
rect 70784 0 70840 400
rect 71008 0 71064 400
rect 71232 0 71288 400
rect 71456 0 71512 400
rect 71680 0 71736 400
rect 71904 0 71960 400
rect 72128 0 72184 400
rect 72352 0 72408 400
rect 72576 0 72632 400
rect 72800 0 72856 400
rect 73024 0 73080 400
rect 73248 0 73304 400
rect 73472 0 73528 400
rect 73696 0 73752 400
rect 73920 0 73976 400
rect 74144 0 74200 400
rect 74368 0 74424 400
rect 74592 0 74648 400
rect 74816 0 74872 400
rect 75040 0 75096 400
rect 75264 0 75320 400
rect 75488 0 75544 400
rect 75712 0 75768 400
rect 75936 0 75992 400
rect 76160 0 76216 400
rect 76384 0 76440 400
rect 76608 0 76664 400
rect 76832 0 76888 400
rect 77056 0 77112 400
rect 77280 0 77336 400
rect 77504 0 77560 400
rect 77728 0 77784 400
rect 77952 0 78008 400
rect 78176 0 78232 400
rect 78400 0 78456 400
rect 78624 0 78680 400
rect 78848 0 78904 400
rect 79072 0 79128 400
rect 79296 0 79352 400
rect 79520 0 79576 400
rect 79744 0 79800 400
rect 79968 0 80024 400
rect 80192 0 80248 400
rect 80416 0 80472 400
rect 80640 0 80696 400
rect 80864 0 80920 400
rect 81088 0 81144 400
rect 81312 0 81368 400
rect 81536 0 81592 400
rect 81760 0 81816 400
rect 81984 0 82040 400
rect 82208 0 82264 400
rect 82432 0 82488 400
rect 82656 0 82712 400
rect 82880 0 82936 400
rect 83104 0 83160 400
rect 83328 0 83384 400
rect 83552 0 83608 400
rect 83776 0 83832 400
rect 84000 0 84056 400
rect 84224 0 84280 400
rect 84448 0 84504 400
rect 84672 0 84728 400
rect 84896 0 84952 400
rect 85120 0 85176 400
rect 85344 0 85400 400
rect 85568 0 85624 400
rect 85792 0 85848 400
rect 86016 0 86072 400
rect 86240 0 86296 400
rect 86464 0 86520 400
rect 86688 0 86744 400
rect 86912 0 86968 400
rect 87136 0 87192 400
rect 87360 0 87416 400
rect 87584 0 87640 400
rect 87808 0 87864 400
rect 88032 0 88088 400
rect 88256 0 88312 400
rect 88480 0 88536 400
rect 88704 0 88760 400
rect 88928 0 88984 400
rect 89152 0 89208 400
rect 89376 0 89432 400
rect 89600 0 89656 400
rect 89824 0 89880 400
rect 90048 0 90104 400
rect 90272 0 90328 400
rect 90496 0 90552 400
rect 90720 0 90776 400
rect 90944 0 91000 400
rect 91168 0 91224 400
rect 91392 0 91448 400
rect 91616 0 91672 400
rect 91840 0 91896 400
rect 92064 0 92120 400
rect 92288 0 92344 400
rect 92512 0 92568 400
rect 92736 0 92792 400
rect 92960 0 93016 400
rect 93184 0 93240 400
rect 93408 0 93464 400
rect 93632 0 93688 400
rect 93856 0 93912 400
rect 94080 0 94136 400
rect 94304 0 94360 400
rect 94528 0 94584 400
rect 94752 0 94808 400
rect 94976 0 95032 400
rect 95200 0 95256 400
rect 95424 0 95480 400
rect 95648 0 95704 400
rect 95872 0 95928 400
rect 96096 0 96152 400
rect 96320 0 96376 400
rect 96544 0 96600 400
rect 96768 0 96824 400
rect 96992 0 97048 400
rect 97216 0 97272 400
rect 97440 0 97496 400
rect 97664 0 97720 400
rect 97888 0 97944 400
rect 98112 0 98168 400
rect 98336 0 98392 400
rect 98560 0 98616 400
rect 98784 0 98840 400
rect 99008 0 99064 400
rect 99232 0 99288 400
rect 99456 0 99512 400
rect 99680 0 99736 400
rect 99904 0 99960 400
rect 100128 0 100184 400
rect 100352 0 100408 400
rect 100576 0 100632 400
rect 100800 0 100856 400
rect 101024 0 101080 400
rect 101248 0 101304 400
rect 101472 0 101528 400
rect 101696 0 101752 400
rect 101920 0 101976 400
rect 102144 0 102200 400
rect 102368 0 102424 400
rect 102592 0 102648 400
rect 102816 0 102872 400
rect 103040 0 103096 400
rect 103264 0 103320 400
rect 103488 0 103544 400
rect 103712 0 103768 400
rect 103936 0 103992 400
rect 104160 0 104216 400
rect 104384 0 104440 400
rect 104608 0 104664 400
rect 104832 0 104888 400
rect 105056 0 105112 400
rect 105280 0 105336 400
rect 105504 0 105560 400
rect 105728 0 105784 400
rect 105952 0 106008 400
rect 106176 0 106232 400
rect 106400 0 106456 400
rect 106624 0 106680 400
rect 106848 0 106904 400
rect 107072 0 107128 400
rect 107296 0 107352 400
rect 107520 0 107576 400
rect 107744 0 107800 400
rect 107968 0 108024 400
rect 108192 0 108248 400
rect 108416 0 108472 400
rect 108640 0 108696 400
rect 108864 0 108920 400
rect 109088 0 109144 400
rect 109312 0 109368 400
rect 109536 0 109592 400
rect 109760 0 109816 400
rect 109984 0 110040 400
rect 110208 0 110264 400
rect 110432 0 110488 400
rect 110656 0 110712 400
rect 110880 0 110936 400
rect 111104 0 111160 400
rect 111328 0 111384 400
rect 111552 0 111608 400
rect 111776 0 111832 400
rect 112000 0 112056 400
rect 112224 0 112280 400
rect 112448 0 112504 400
rect 112672 0 112728 400
rect 112896 0 112952 400
rect 113120 0 113176 400
rect 113344 0 113400 400
rect 113568 0 113624 400
rect 113792 0 113848 400
rect 114016 0 114072 400
rect 114240 0 114296 400
rect 114464 0 114520 400
rect 114688 0 114744 400
rect 114912 0 114968 400
<< obsm2 >>
rect 630 34570 2994 34650
rect 3110 34570 3890 34650
rect 4006 34570 4786 34650
rect 4902 34570 5682 34650
rect 5798 34570 6578 34650
rect 6694 34570 7474 34650
rect 7590 34570 8370 34650
rect 8486 34570 9266 34650
rect 9382 34570 10162 34650
rect 10278 34570 11058 34650
rect 11174 34570 11954 34650
rect 12070 34570 12850 34650
rect 12966 34570 13746 34650
rect 13862 34570 14642 34650
rect 14758 34570 15538 34650
rect 15654 34570 16434 34650
rect 16550 34570 17330 34650
rect 17446 34570 18226 34650
rect 18342 34570 19122 34650
rect 19238 34570 20018 34650
rect 20134 34570 20914 34650
rect 21030 34570 21810 34650
rect 21926 34570 22706 34650
rect 22822 34570 23602 34650
rect 23718 34570 24498 34650
rect 24614 34570 25394 34650
rect 25510 34570 26290 34650
rect 26406 34570 27186 34650
rect 27302 34570 28082 34650
rect 28198 34570 28978 34650
rect 29094 34570 29874 34650
rect 29990 34570 30770 34650
rect 30886 34570 31666 34650
rect 31782 34570 32562 34650
rect 32678 34570 33458 34650
rect 33574 34570 34354 34650
rect 34470 34570 35250 34650
rect 35366 34570 36146 34650
rect 36262 34570 37042 34650
rect 37158 34570 37938 34650
rect 38054 34570 38834 34650
rect 38950 34570 39730 34650
rect 39846 34570 40626 34650
rect 40742 34570 41522 34650
rect 41638 34570 42418 34650
rect 42534 34570 43314 34650
rect 43430 34570 44210 34650
rect 44326 34570 45106 34650
rect 45222 34570 46002 34650
rect 46118 34570 46898 34650
rect 47014 34570 47794 34650
rect 47910 34570 48690 34650
rect 48806 34570 49586 34650
rect 49702 34570 50482 34650
rect 50598 34570 51378 34650
rect 51494 34570 52274 34650
rect 52390 34570 53170 34650
rect 53286 34570 54066 34650
rect 54182 34570 54962 34650
rect 55078 34570 55858 34650
rect 55974 34570 56754 34650
rect 56870 34570 57650 34650
rect 57766 34570 58546 34650
rect 58662 34570 59442 34650
rect 59558 34570 60338 34650
rect 60454 34570 61234 34650
rect 61350 34570 62130 34650
rect 62246 34570 63026 34650
rect 63142 34570 63922 34650
rect 64038 34570 64818 34650
rect 64934 34570 65714 34650
rect 65830 34570 66610 34650
rect 66726 34570 67506 34650
rect 67622 34570 68402 34650
rect 68518 34570 69298 34650
rect 69414 34570 70194 34650
rect 70310 34570 71090 34650
rect 71206 34570 71986 34650
rect 72102 34570 72882 34650
rect 72998 34570 73778 34650
rect 73894 34570 74674 34650
rect 74790 34570 75570 34650
rect 75686 34570 76466 34650
rect 76582 34570 77362 34650
rect 77478 34570 78258 34650
rect 78374 34570 79154 34650
rect 79270 34570 80050 34650
rect 80166 34570 80946 34650
rect 81062 34570 81842 34650
rect 81958 34570 82738 34650
rect 82854 34570 83634 34650
rect 83750 34570 84530 34650
rect 84646 34570 85426 34650
rect 85542 34570 86322 34650
rect 86438 34570 87218 34650
rect 87334 34570 88114 34650
rect 88230 34570 89010 34650
rect 89126 34570 89906 34650
rect 90022 34570 90802 34650
rect 90918 34570 91698 34650
rect 91814 34570 92594 34650
rect 92710 34570 93490 34650
rect 93606 34570 94386 34650
rect 94502 34570 95282 34650
rect 95398 34570 96178 34650
rect 96294 34570 97074 34650
rect 97190 34570 97970 34650
rect 98086 34570 98866 34650
rect 98982 34570 99762 34650
rect 99878 34570 100658 34650
rect 100774 34570 101554 34650
rect 101670 34570 102450 34650
rect 102566 34570 103346 34650
rect 103462 34570 104242 34650
rect 104358 34570 105138 34650
rect 105254 34570 106034 34650
rect 106150 34570 106930 34650
rect 107046 34570 107826 34650
rect 107942 34570 108722 34650
rect 108838 34570 109618 34650
rect 109734 34570 110514 34650
rect 110630 34570 111410 34650
rect 111526 34570 112306 34650
rect 112422 34570 113202 34650
rect 113318 34570 114098 34650
rect 114214 34570 114994 34650
rect 115110 34570 115890 34650
rect 116006 34570 116786 34650
rect 116902 34570 119322 34650
rect 630 430 119322 34570
rect 630 177 4898 430
rect 5014 177 5122 430
rect 5238 177 5346 430
rect 5462 177 5570 430
rect 5686 177 5794 430
rect 5910 177 6018 430
rect 6134 177 6242 430
rect 6358 177 6466 430
rect 6582 177 6690 430
rect 6806 177 6914 430
rect 7030 177 7138 430
rect 7254 177 7362 430
rect 7478 177 7586 430
rect 7702 177 7810 430
rect 7926 177 8034 430
rect 8150 177 8258 430
rect 8374 177 8482 430
rect 8598 177 8706 430
rect 8822 177 8930 430
rect 9046 177 9154 430
rect 9270 177 9378 430
rect 9494 177 9602 430
rect 9718 177 9826 430
rect 9942 177 10050 430
rect 10166 177 10274 430
rect 10390 177 10498 430
rect 10614 177 10722 430
rect 10838 177 10946 430
rect 11062 177 11170 430
rect 11286 177 11394 430
rect 11510 177 11618 430
rect 11734 177 11842 430
rect 11958 177 12066 430
rect 12182 177 12290 430
rect 12406 177 12514 430
rect 12630 177 12738 430
rect 12854 177 12962 430
rect 13078 177 13186 430
rect 13302 177 13410 430
rect 13526 177 13634 430
rect 13750 177 13858 430
rect 13974 177 14082 430
rect 14198 177 14306 430
rect 14422 177 14530 430
rect 14646 177 14754 430
rect 14870 177 14978 430
rect 15094 177 15202 430
rect 15318 177 15426 430
rect 15542 177 15650 430
rect 15766 177 15874 430
rect 15990 177 16098 430
rect 16214 177 16322 430
rect 16438 177 16546 430
rect 16662 177 16770 430
rect 16886 177 16994 430
rect 17110 177 17218 430
rect 17334 177 17442 430
rect 17558 177 17666 430
rect 17782 177 17890 430
rect 18006 177 18114 430
rect 18230 177 18338 430
rect 18454 177 18562 430
rect 18678 177 18786 430
rect 18902 177 19010 430
rect 19126 177 19234 430
rect 19350 177 19458 430
rect 19574 177 19682 430
rect 19798 177 19906 430
rect 20022 177 20130 430
rect 20246 177 20354 430
rect 20470 177 20578 430
rect 20694 177 20802 430
rect 20918 177 21026 430
rect 21142 177 21250 430
rect 21366 177 21474 430
rect 21590 177 21698 430
rect 21814 177 21922 430
rect 22038 177 22146 430
rect 22262 177 22370 430
rect 22486 177 22594 430
rect 22710 177 22818 430
rect 22934 177 23042 430
rect 23158 177 23266 430
rect 23382 177 23490 430
rect 23606 177 23714 430
rect 23830 177 23938 430
rect 24054 177 24162 430
rect 24278 177 24386 430
rect 24502 177 24610 430
rect 24726 177 24834 430
rect 24950 177 25058 430
rect 25174 177 25282 430
rect 25398 177 25506 430
rect 25622 177 25730 430
rect 25846 177 25954 430
rect 26070 177 26178 430
rect 26294 177 26402 430
rect 26518 177 26626 430
rect 26742 177 26850 430
rect 26966 177 27074 430
rect 27190 177 27298 430
rect 27414 177 27522 430
rect 27638 177 27746 430
rect 27862 177 27970 430
rect 28086 177 28194 430
rect 28310 177 28418 430
rect 28534 177 28642 430
rect 28758 177 28866 430
rect 28982 177 29090 430
rect 29206 177 29314 430
rect 29430 177 29538 430
rect 29654 177 29762 430
rect 29878 177 29986 430
rect 30102 177 30210 430
rect 30326 177 30434 430
rect 30550 177 30658 430
rect 30774 177 30882 430
rect 30998 177 31106 430
rect 31222 177 31330 430
rect 31446 177 31554 430
rect 31670 177 31778 430
rect 31894 177 32002 430
rect 32118 177 32226 430
rect 32342 177 32450 430
rect 32566 177 32674 430
rect 32790 177 32898 430
rect 33014 177 33122 430
rect 33238 177 33346 430
rect 33462 177 33570 430
rect 33686 177 33794 430
rect 33910 177 34018 430
rect 34134 177 34242 430
rect 34358 177 34466 430
rect 34582 177 34690 430
rect 34806 177 34914 430
rect 35030 177 35138 430
rect 35254 177 35362 430
rect 35478 177 35586 430
rect 35702 177 35810 430
rect 35926 177 36034 430
rect 36150 177 36258 430
rect 36374 177 36482 430
rect 36598 177 36706 430
rect 36822 177 36930 430
rect 37046 177 37154 430
rect 37270 177 37378 430
rect 37494 177 37602 430
rect 37718 177 37826 430
rect 37942 177 38050 430
rect 38166 177 38274 430
rect 38390 177 38498 430
rect 38614 177 38722 430
rect 38838 177 38946 430
rect 39062 177 39170 430
rect 39286 177 39394 430
rect 39510 177 39618 430
rect 39734 177 39842 430
rect 39958 177 40066 430
rect 40182 177 40290 430
rect 40406 177 40514 430
rect 40630 177 40738 430
rect 40854 177 40962 430
rect 41078 177 41186 430
rect 41302 177 41410 430
rect 41526 177 41634 430
rect 41750 177 41858 430
rect 41974 177 42082 430
rect 42198 177 42306 430
rect 42422 177 42530 430
rect 42646 177 42754 430
rect 42870 177 42978 430
rect 43094 177 43202 430
rect 43318 177 43426 430
rect 43542 177 43650 430
rect 43766 177 43874 430
rect 43990 177 44098 430
rect 44214 177 44322 430
rect 44438 177 44546 430
rect 44662 177 44770 430
rect 44886 177 44994 430
rect 45110 177 45218 430
rect 45334 177 45442 430
rect 45558 177 45666 430
rect 45782 177 45890 430
rect 46006 177 46114 430
rect 46230 177 46338 430
rect 46454 177 46562 430
rect 46678 177 46786 430
rect 46902 177 47010 430
rect 47126 177 47234 430
rect 47350 177 47458 430
rect 47574 177 47682 430
rect 47798 177 47906 430
rect 48022 177 48130 430
rect 48246 177 48354 430
rect 48470 177 48578 430
rect 48694 177 48802 430
rect 48918 177 49026 430
rect 49142 177 49250 430
rect 49366 177 49474 430
rect 49590 177 49698 430
rect 49814 177 49922 430
rect 50038 177 50146 430
rect 50262 177 50370 430
rect 50486 177 50594 430
rect 50710 177 50818 430
rect 50934 177 51042 430
rect 51158 177 51266 430
rect 51382 177 51490 430
rect 51606 177 51714 430
rect 51830 177 51938 430
rect 52054 177 52162 430
rect 52278 177 52386 430
rect 52502 177 52610 430
rect 52726 177 52834 430
rect 52950 177 53058 430
rect 53174 177 53282 430
rect 53398 177 53506 430
rect 53622 177 53730 430
rect 53846 177 53954 430
rect 54070 177 54178 430
rect 54294 177 54402 430
rect 54518 177 54626 430
rect 54742 177 54850 430
rect 54966 177 55074 430
rect 55190 177 55298 430
rect 55414 177 55522 430
rect 55638 177 55746 430
rect 55862 177 55970 430
rect 56086 177 56194 430
rect 56310 177 56418 430
rect 56534 177 56642 430
rect 56758 177 56866 430
rect 56982 177 57090 430
rect 57206 177 57314 430
rect 57430 177 57538 430
rect 57654 177 57762 430
rect 57878 177 57986 430
rect 58102 177 58210 430
rect 58326 177 58434 430
rect 58550 177 58658 430
rect 58774 177 58882 430
rect 58998 177 59106 430
rect 59222 177 59330 430
rect 59446 177 59554 430
rect 59670 177 59778 430
rect 59894 177 60002 430
rect 60118 177 60226 430
rect 60342 177 60450 430
rect 60566 177 60674 430
rect 60790 177 60898 430
rect 61014 177 61122 430
rect 61238 177 61346 430
rect 61462 177 61570 430
rect 61686 177 61794 430
rect 61910 177 62018 430
rect 62134 177 62242 430
rect 62358 177 62466 430
rect 62582 177 62690 430
rect 62806 177 62914 430
rect 63030 177 63138 430
rect 63254 177 63362 430
rect 63478 177 63586 430
rect 63702 177 63810 430
rect 63926 177 64034 430
rect 64150 177 64258 430
rect 64374 177 64482 430
rect 64598 177 64706 430
rect 64822 177 64930 430
rect 65046 177 65154 430
rect 65270 177 65378 430
rect 65494 177 65602 430
rect 65718 177 65826 430
rect 65942 177 66050 430
rect 66166 177 66274 430
rect 66390 177 66498 430
rect 66614 177 66722 430
rect 66838 177 66946 430
rect 67062 177 67170 430
rect 67286 177 67394 430
rect 67510 177 67618 430
rect 67734 177 67842 430
rect 67958 177 68066 430
rect 68182 177 68290 430
rect 68406 177 68514 430
rect 68630 177 68738 430
rect 68854 177 68962 430
rect 69078 177 69186 430
rect 69302 177 69410 430
rect 69526 177 69634 430
rect 69750 177 69858 430
rect 69974 177 70082 430
rect 70198 177 70306 430
rect 70422 177 70530 430
rect 70646 177 70754 430
rect 70870 177 70978 430
rect 71094 177 71202 430
rect 71318 177 71426 430
rect 71542 177 71650 430
rect 71766 177 71874 430
rect 71990 177 72098 430
rect 72214 177 72322 430
rect 72438 177 72546 430
rect 72662 177 72770 430
rect 72886 177 72994 430
rect 73110 177 73218 430
rect 73334 177 73442 430
rect 73558 177 73666 430
rect 73782 177 73890 430
rect 74006 177 74114 430
rect 74230 177 74338 430
rect 74454 177 74562 430
rect 74678 177 74786 430
rect 74902 177 75010 430
rect 75126 177 75234 430
rect 75350 177 75458 430
rect 75574 177 75682 430
rect 75798 177 75906 430
rect 76022 177 76130 430
rect 76246 177 76354 430
rect 76470 177 76578 430
rect 76694 177 76802 430
rect 76918 177 77026 430
rect 77142 177 77250 430
rect 77366 177 77474 430
rect 77590 177 77698 430
rect 77814 177 77922 430
rect 78038 177 78146 430
rect 78262 177 78370 430
rect 78486 177 78594 430
rect 78710 177 78818 430
rect 78934 177 79042 430
rect 79158 177 79266 430
rect 79382 177 79490 430
rect 79606 177 79714 430
rect 79830 177 79938 430
rect 80054 177 80162 430
rect 80278 177 80386 430
rect 80502 177 80610 430
rect 80726 177 80834 430
rect 80950 177 81058 430
rect 81174 177 81282 430
rect 81398 177 81506 430
rect 81622 177 81730 430
rect 81846 177 81954 430
rect 82070 177 82178 430
rect 82294 177 82402 430
rect 82518 177 82626 430
rect 82742 177 82850 430
rect 82966 177 83074 430
rect 83190 177 83298 430
rect 83414 177 83522 430
rect 83638 177 83746 430
rect 83862 177 83970 430
rect 84086 177 84194 430
rect 84310 177 84418 430
rect 84534 177 84642 430
rect 84758 177 84866 430
rect 84982 177 85090 430
rect 85206 177 85314 430
rect 85430 177 85538 430
rect 85654 177 85762 430
rect 85878 177 85986 430
rect 86102 177 86210 430
rect 86326 177 86434 430
rect 86550 177 86658 430
rect 86774 177 86882 430
rect 86998 177 87106 430
rect 87222 177 87330 430
rect 87446 177 87554 430
rect 87670 177 87778 430
rect 87894 177 88002 430
rect 88118 177 88226 430
rect 88342 177 88450 430
rect 88566 177 88674 430
rect 88790 177 88898 430
rect 89014 177 89122 430
rect 89238 177 89346 430
rect 89462 177 89570 430
rect 89686 177 89794 430
rect 89910 177 90018 430
rect 90134 177 90242 430
rect 90358 177 90466 430
rect 90582 177 90690 430
rect 90806 177 90914 430
rect 91030 177 91138 430
rect 91254 177 91362 430
rect 91478 177 91586 430
rect 91702 177 91810 430
rect 91926 177 92034 430
rect 92150 177 92258 430
rect 92374 177 92482 430
rect 92598 177 92706 430
rect 92822 177 92930 430
rect 93046 177 93154 430
rect 93270 177 93378 430
rect 93494 177 93602 430
rect 93718 177 93826 430
rect 93942 177 94050 430
rect 94166 177 94274 430
rect 94390 177 94498 430
rect 94614 177 94722 430
rect 94838 177 94946 430
rect 95062 177 95170 430
rect 95286 177 95394 430
rect 95510 177 95618 430
rect 95734 177 95842 430
rect 95958 177 96066 430
rect 96182 177 96290 430
rect 96406 177 96514 430
rect 96630 177 96738 430
rect 96854 177 96962 430
rect 97078 177 97186 430
rect 97302 177 97410 430
rect 97526 177 97634 430
rect 97750 177 97858 430
rect 97974 177 98082 430
rect 98198 177 98306 430
rect 98422 177 98530 430
rect 98646 177 98754 430
rect 98870 177 98978 430
rect 99094 177 99202 430
rect 99318 177 99426 430
rect 99542 177 99650 430
rect 99766 177 99874 430
rect 99990 177 100098 430
rect 100214 177 100322 430
rect 100438 177 100546 430
rect 100662 177 100770 430
rect 100886 177 100994 430
rect 101110 177 101218 430
rect 101334 177 101442 430
rect 101558 177 101666 430
rect 101782 177 101890 430
rect 102006 177 102114 430
rect 102230 177 102338 430
rect 102454 177 102562 430
rect 102678 177 102786 430
rect 102902 177 103010 430
rect 103126 177 103234 430
rect 103350 177 103458 430
rect 103574 177 103682 430
rect 103798 177 103906 430
rect 104022 177 104130 430
rect 104246 177 104354 430
rect 104470 177 104578 430
rect 104694 177 104802 430
rect 104918 177 105026 430
rect 105142 177 105250 430
rect 105366 177 105474 430
rect 105590 177 105698 430
rect 105814 177 105922 430
rect 106038 177 106146 430
rect 106262 177 106370 430
rect 106486 177 106594 430
rect 106710 177 106818 430
rect 106934 177 107042 430
rect 107158 177 107266 430
rect 107382 177 107490 430
rect 107606 177 107714 430
rect 107830 177 107938 430
rect 108054 177 108162 430
rect 108278 177 108386 430
rect 108502 177 108610 430
rect 108726 177 108834 430
rect 108950 177 109058 430
rect 109174 177 109282 430
rect 109398 177 109506 430
rect 109622 177 109730 430
rect 109846 177 109954 430
rect 110070 177 110178 430
rect 110294 177 110402 430
rect 110518 177 110626 430
rect 110742 177 110850 430
rect 110966 177 111074 430
rect 111190 177 111298 430
rect 111414 177 111522 430
rect 111638 177 111746 430
rect 111862 177 111970 430
rect 112086 177 112194 430
rect 112310 177 112418 430
rect 112534 177 112642 430
rect 112758 177 112866 430
rect 112982 177 113090 430
rect 113206 177 113314 430
rect 113430 177 113538 430
rect 113654 177 113762 430
rect 113878 177 113986 430
rect 114102 177 114210 430
rect 114326 177 114434 430
rect 114550 177 114658 430
rect 114774 177 114882 430
rect 114998 177 119322 430
<< metal3 >>
rect 0 32704 400 32760
rect 119600 32704 120000 32760
rect 0 32368 400 32424
rect 119600 32368 120000 32424
rect 0 32032 400 32088
rect 119600 32032 120000 32088
rect 0 31696 400 31752
rect 119600 31696 120000 31752
rect 0 31360 400 31416
rect 119600 31360 120000 31416
rect 0 31024 400 31080
rect 119600 31024 120000 31080
rect 0 30688 400 30744
rect 119600 30688 120000 30744
rect 0 30352 400 30408
rect 119600 30352 120000 30408
rect 0 30016 400 30072
rect 119600 30016 120000 30072
rect 0 29680 400 29736
rect 119600 29680 120000 29736
rect 0 29344 400 29400
rect 119600 29344 120000 29400
rect 0 29008 400 29064
rect 119600 29008 120000 29064
rect 0 28672 400 28728
rect 119600 28672 120000 28728
rect 0 28336 400 28392
rect 119600 28336 120000 28392
rect 0 28000 400 28056
rect 119600 28000 120000 28056
rect 0 27664 400 27720
rect 119600 27664 120000 27720
rect 0 27328 400 27384
rect 119600 27328 120000 27384
rect 0 26992 400 27048
rect 119600 26992 120000 27048
rect 0 26656 400 26712
rect 119600 26656 120000 26712
rect 0 26320 400 26376
rect 119600 26320 120000 26376
rect 0 25984 400 26040
rect 119600 25984 120000 26040
rect 0 25648 400 25704
rect 119600 25648 120000 25704
rect 0 25312 400 25368
rect 119600 25312 120000 25368
rect 0 24976 400 25032
rect 119600 24976 120000 25032
rect 0 24640 400 24696
rect 119600 24640 120000 24696
rect 0 24304 400 24360
rect 119600 24304 120000 24360
rect 0 23968 400 24024
rect 119600 23968 120000 24024
rect 0 23632 400 23688
rect 119600 23632 120000 23688
rect 0 23296 400 23352
rect 119600 23296 120000 23352
rect 0 22960 400 23016
rect 119600 22960 120000 23016
rect 0 22624 400 22680
rect 119600 22624 120000 22680
rect 0 22288 400 22344
rect 119600 22288 120000 22344
rect 0 21952 400 22008
rect 119600 21952 120000 22008
rect 0 21616 400 21672
rect 119600 21616 120000 21672
rect 0 21280 400 21336
rect 119600 21280 120000 21336
rect 0 20944 400 21000
rect 119600 20944 120000 21000
rect 0 20608 400 20664
rect 119600 20608 120000 20664
rect 0 20272 400 20328
rect 119600 20272 120000 20328
rect 0 19936 400 19992
rect 119600 19936 120000 19992
rect 0 19600 400 19656
rect 119600 19600 120000 19656
rect 0 19264 400 19320
rect 119600 19264 120000 19320
rect 0 18928 400 18984
rect 119600 18928 120000 18984
rect 0 18592 400 18648
rect 119600 18592 120000 18648
rect 0 18256 400 18312
rect 119600 18256 120000 18312
rect 0 17920 400 17976
rect 119600 17920 120000 17976
rect 0 17584 400 17640
rect 119600 17584 120000 17640
rect 0 17248 400 17304
rect 119600 17248 120000 17304
rect 0 16912 400 16968
rect 119600 16912 120000 16968
rect 0 16576 400 16632
rect 119600 16576 120000 16632
rect 0 16240 400 16296
rect 119600 16240 120000 16296
rect 0 15904 400 15960
rect 119600 15904 120000 15960
rect 0 15568 400 15624
rect 119600 15568 120000 15624
rect 0 15232 400 15288
rect 119600 15232 120000 15288
rect 0 14896 400 14952
rect 119600 14896 120000 14952
rect 0 14560 400 14616
rect 119600 14560 120000 14616
rect 0 14224 400 14280
rect 119600 14224 120000 14280
rect 0 13888 400 13944
rect 119600 13888 120000 13944
rect 0 13552 400 13608
rect 119600 13552 120000 13608
rect 0 13216 400 13272
rect 119600 13216 120000 13272
rect 0 12880 400 12936
rect 119600 12880 120000 12936
rect 0 12544 400 12600
rect 119600 12544 120000 12600
rect 0 12208 400 12264
rect 119600 12208 120000 12264
rect 0 11872 400 11928
rect 119600 11872 120000 11928
rect 0 11536 400 11592
rect 119600 11536 120000 11592
rect 0 11200 400 11256
rect 119600 11200 120000 11256
rect 0 10864 400 10920
rect 119600 10864 120000 10920
rect 0 10528 400 10584
rect 119600 10528 120000 10584
rect 0 10192 400 10248
rect 119600 10192 120000 10248
rect 0 9856 400 9912
rect 119600 9856 120000 9912
rect 0 9520 400 9576
rect 119600 9520 120000 9576
rect 0 9184 400 9240
rect 119600 9184 120000 9240
rect 0 8848 400 8904
rect 119600 8848 120000 8904
rect 0 8512 400 8568
rect 119600 8512 120000 8568
rect 0 8176 400 8232
rect 119600 8176 120000 8232
rect 0 7840 400 7896
rect 119600 7840 120000 7896
rect 0 7504 400 7560
rect 119600 7504 120000 7560
rect 0 7168 400 7224
rect 119600 7168 120000 7224
rect 0 6832 400 6888
rect 119600 6832 120000 6888
rect 0 6496 400 6552
rect 119600 6496 120000 6552
rect 0 6160 400 6216
rect 119600 6160 120000 6216
rect 0 5824 400 5880
rect 119600 5824 120000 5880
rect 0 5488 400 5544
rect 119600 5488 120000 5544
rect 0 5152 400 5208
rect 119600 5152 120000 5208
rect 0 4816 400 4872
rect 119600 4816 120000 4872
rect 0 4480 400 4536
rect 119600 4480 120000 4536
rect 0 4144 400 4200
rect 119600 4144 120000 4200
rect 0 3808 400 3864
rect 119600 3808 120000 3864
rect 0 3472 400 3528
rect 119600 3472 120000 3528
rect 0 3136 400 3192
rect 119600 3136 120000 3192
rect 0 2800 400 2856
rect 119600 2800 120000 2856
rect 0 2464 400 2520
rect 119600 2464 120000 2520
rect 0 2128 400 2184
rect 119600 2128 120000 2184
<< obsm3 >>
rect 400 32790 119600 34034
rect 430 32674 119570 32790
rect 400 32454 119600 32674
rect 430 32338 119570 32454
rect 400 32118 119600 32338
rect 430 32002 119570 32118
rect 400 31782 119600 32002
rect 430 31666 119570 31782
rect 400 31446 119600 31666
rect 430 31330 119570 31446
rect 400 31110 119600 31330
rect 430 30994 119570 31110
rect 400 30774 119600 30994
rect 430 30658 119570 30774
rect 400 30438 119600 30658
rect 430 30322 119570 30438
rect 400 30102 119600 30322
rect 430 29986 119570 30102
rect 400 29766 119600 29986
rect 430 29650 119570 29766
rect 400 29430 119600 29650
rect 430 29314 119570 29430
rect 400 29094 119600 29314
rect 430 28978 119570 29094
rect 400 28758 119600 28978
rect 430 28642 119570 28758
rect 400 28422 119600 28642
rect 430 28306 119570 28422
rect 400 28086 119600 28306
rect 430 27970 119570 28086
rect 400 27750 119600 27970
rect 430 27634 119570 27750
rect 400 27414 119600 27634
rect 430 27298 119570 27414
rect 400 27078 119600 27298
rect 430 26962 119570 27078
rect 400 26742 119600 26962
rect 430 26626 119570 26742
rect 400 26406 119600 26626
rect 430 26290 119570 26406
rect 400 26070 119600 26290
rect 430 25954 119570 26070
rect 400 25734 119600 25954
rect 430 25618 119570 25734
rect 400 25398 119600 25618
rect 430 25282 119570 25398
rect 400 25062 119600 25282
rect 430 24946 119570 25062
rect 400 24726 119600 24946
rect 430 24610 119570 24726
rect 400 24390 119600 24610
rect 430 24274 119570 24390
rect 400 24054 119600 24274
rect 430 23938 119570 24054
rect 400 23718 119600 23938
rect 430 23602 119570 23718
rect 400 23382 119600 23602
rect 430 23266 119570 23382
rect 400 23046 119600 23266
rect 430 22930 119570 23046
rect 400 22710 119600 22930
rect 430 22594 119570 22710
rect 400 22374 119600 22594
rect 430 22258 119570 22374
rect 400 22038 119600 22258
rect 430 21922 119570 22038
rect 400 21702 119600 21922
rect 430 21586 119570 21702
rect 400 21366 119600 21586
rect 430 21250 119570 21366
rect 400 21030 119600 21250
rect 430 20914 119570 21030
rect 400 20694 119600 20914
rect 430 20578 119570 20694
rect 400 20358 119600 20578
rect 430 20242 119570 20358
rect 400 20022 119600 20242
rect 430 19906 119570 20022
rect 400 19686 119600 19906
rect 430 19570 119570 19686
rect 400 19350 119600 19570
rect 430 19234 119570 19350
rect 400 19014 119600 19234
rect 430 18898 119570 19014
rect 400 18678 119600 18898
rect 430 18562 119570 18678
rect 400 18342 119600 18562
rect 430 18226 119570 18342
rect 400 18006 119600 18226
rect 430 17890 119570 18006
rect 400 17670 119600 17890
rect 430 17554 119570 17670
rect 400 17334 119600 17554
rect 430 17218 119570 17334
rect 400 16998 119600 17218
rect 430 16882 119570 16998
rect 400 16662 119600 16882
rect 430 16546 119570 16662
rect 400 16326 119600 16546
rect 430 16210 119570 16326
rect 400 15990 119600 16210
rect 430 15874 119570 15990
rect 400 15654 119600 15874
rect 430 15538 119570 15654
rect 400 15318 119600 15538
rect 430 15202 119570 15318
rect 400 14982 119600 15202
rect 430 14866 119570 14982
rect 400 14646 119600 14866
rect 430 14530 119570 14646
rect 400 14310 119600 14530
rect 430 14194 119570 14310
rect 400 13974 119600 14194
rect 430 13858 119570 13974
rect 400 13638 119600 13858
rect 430 13522 119570 13638
rect 400 13302 119600 13522
rect 430 13186 119570 13302
rect 400 12966 119600 13186
rect 430 12850 119570 12966
rect 400 12630 119600 12850
rect 430 12514 119570 12630
rect 400 12294 119600 12514
rect 430 12178 119570 12294
rect 400 11958 119600 12178
rect 430 11842 119570 11958
rect 400 11622 119600 11842
rect 430 11506 119570 11622
rect 400 11286 119600 11506
rect 430 11170 119570 11286
rect 400 10950 119600 11170
rect 430 10834 119570 10950
rect 400 10614 119600 10834
rect 430 10498 119570 10614
rect 400 10278 119600 10498
rect 430 10162 119570 10278
rect 400 9942 119600 10162
rect 430 9826 119570 9942
rect 400 9606 119600 9826
rect 430 9490 119570 9606
rect 400 9270 119600 9490
rect 430 9154 119570 9270
rect 400 8934 119600 9154
rect 430 8818 119570 8934
rect 400 8598 119600 8818
rect 430 8482 119570 8598
rect 400 8262 119600 8482
rect 430 8146 119570 8262
rect 400 7926 119600 8146
rect 430 7810 119570 7926
rect 400 7590 119600 7810
rect 430 7474 119570 7590
rect 400 7254 119600 7474
rect 430 7138 119570 7254
rect 400 6918 119600 7138
rect 430 6802 119570 6918
rect 400 6582 119600 6802
rect 430 6466 119570 6582
rect 400 6246 119600 6466
rect 430 6130 119570 6246
rect 400 5910 119600 6130
rect 430 5794 119570 5910
rect 400 5574 119600 5794
rect 430 5458 119570 5574
rect 400 5238 119600 5458
rect 430 5122 119570 5238
rect 400 4902 119600 5122
rect 430 4786 119570 4902
rect 400 4566 119600 4786
rect 430 4450 119570 4566
rect 400 4230 119600 4450
rect 430 4114 119570 4230
rect 400 3894 119600 4114
rect 430 3778 119570 3894
rect 400 3558 119600 3778
rect 430 3442 119570 3558
rect 400 3222 119600 3442
rect 430 3106 119570 3222
rect 400 2886 119600 3106
rect 430 2770 119570 2886
rect 400 2550 119600 2770
rect 430 2434 119570 2550
rect 400 2214 119600 2434
rect 430 2098 119570 2214
rect 400 182 119600 2098
<< metal4 >>
rect 2224 1538 2384 33350
rect 9904 1538 10064 33350
rect 17584 1538 17744 33350
rect 25264 1538 25424 33350
rect 32944 1538 33104 33350
rect 40624 1538 40784 33350
rect 48304 1538 48464 33350
rect 55984 1538 56144 33350
rect 63664 1538 63824 33350
rect 71344 1538 71504 33350
rect 79024 1538 79184 33350
rect 86704 1538 86864 33350
rect 94384 1538 94544 33350
rect 102064 1538 102224 33350
rect 109744 1538 109904 33350
rect 117424 1538 117584 33350
<< obsm4 >>
rect 910 33380 118202 33759
rect 910 1508 2194 33380
rect 2414 1508 9874 33380
rect 10094 1508 17554 33380
rect 17774 1508 25234 33380
rect 25454 1508 32914 33380
rect 33134 1508 40594 33380
rect 40814 1508 48274 33380
rect 48494 1508 55954 33380
rect 56174 1508 63634 33380
rect 63854 1508 71314 33380
rect 71534 1508 78994 33380
rect 79214 1508 86674 33380
rect 86894 1508 94354 33380
rect 94574 1508 102034 33380
rect 102254 1508 109714 33380
rect 109934 1508 117394 33380
rect 117614 1508 118202 33380
rect 910 457 118202 1508
<< labels >>
rlabel metal2 s 8736 0 8792 400 6 c0_dbg_pc[0]
port 1 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 c0_dbg_pc[10]
port 2 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 c0_dbg_pc[11]
port 3 nsew signal input
rlabel metal2 s 39648 0 39704 400 6 c0_dbg_pc[12]
port 4 nsew signal input
rlabel metal2 s 41888 0 41944 400 6 c0_dbg_pc[13]
port 5 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 c0_dbg_pc[14]
port 6 nsew signal input
rlabel metal2 s 46368 0 46424 400 6 c0_dbg_pc[15]
port 7 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 c0_dbg_pc[1]
port 8 nsew signal input
rlabel metal2 s 14560 0 14616 400 6 c0_dbg_pc[2]
port 9 nsew signal input
rlabel metal2 s 17248 0 17304 400 6 c0_dbg_pc[3]
port 10 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 c0_dbg_pc[4]
port 11 nsew signal input
rlabel metal2 s 22624 0 22680 400 6 c0_dbg_pc[5]
port 12 nsew signal input
rlabel metal2 s 25312 0 25368 400 6 c0_dbg_pc[6]
port 13 nsew signal input
rlabel metal2 s 28000 0 28056 400 6 c0_dbg_pc[7]
port 14 nsew signal input
rlabel metal2 s 30688 0 30744 400 6 c0_dbg_pc[8]
port 15 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 c0_dbg_pc[9]
port 16 nsew signal input
rlabel metal2 s 8960 0 9016 400 6 c0_dbg_r0[0]
port 17 nsew signal input
rlabel metal2 s 35392 0 35448 400 6 c0_dbg_r0[10]
port 18 nsew signal input
rlabel metal2 s 37632 0 37688 400 6 c0_dbg_r0[11]
port 19 nsew signal input
rlabel metal2 s 39872 0 39928 400 6 c0_dbg_r0[12]
port 20 nsew signal input
rlabel metal2 s 42112 0 42168 400 6 c0_dbg_r0[13]
port 21 nsew signal input
rlabel metal2 s 44352 0 44408 400 6 c0_dbg_r0[14]
port 22 nsew signal input
rlabel metal2 s 46592 0 46648 400 6 c0_dbg_r0[15]
port 23 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 c0_dbg_r0[1]
port 24 nsew signal input
rlabel metal2 s 14784 0 14840 400 6 c0_dbg_r0[2]
port 25 nsew signal input
rlabel metal2 s 17472 0 17528 400 6 c0_dbg_r0[3]
port 26 nsew signal input
rlabel metal2 s 20160 0 20216 400 6 c0_dbg_r0[4]
port 27 nsew signal input
rlabel metal2 s 22848 0 22904 400 6 c0_dbg_r0[5]
port 28 nsew signal input
rlabel metal2 s 25536 0 25592 400 6 c0_dbg_r0[6]
port 29 nsew signal input
rlabel metal2 s 28224 0 28280 400 6 c0_dbg_r0[7]
port 30 nsew signal input
rlabel metal2 s 30912 0 30968 400 6 c0_dbg_r0[8]
port 31 nsew signal input
rlabel metal2 s 33152 0 33208 400 6 c0_dbg_r0[9]
port 32 nsew signal input
rlabel metal2 s 4928 0 4984 400 6 c0_disable
port 33 nsew signal output
rlabel metal2 s 9184 0 9240 400 6 c0_i_core_int_sreg[0]
port 34 nsew signal output
rlabel metal2 s 35616 0 35672 400 6 c0_i_core_int_sreg[10]
port 35 nsew signal output
rlabel metal2 s 37856 0 37912 400 6 c0_i_core_int_sreg[11]
port 36 nsew signal output
rlabel metal2 s 40096 0 40152 400 6 c0_i_core_int_sreg[12]
port 37 nsew signal output
rlabel metal2 s 42336 0 42392 400 6 c0_i_core_int_sreg[13]
port 38 nsew signal output
rlabel metal2 s 44576 0 44632 400 6 c0_i_core_int_sreg[14]
port 39 nsew signal output
rlabel metal2 s 46816 0 46872 400 6 c0_i_core_int_sreg[15]
port 40 nsew signal output
rlabel metal2 s 12096 0 12152 400 6 c0_i_core_int_sreg[1]
port 41 nsew signal output
rlabel metal2 s 15008 0 15064 400 6 c0_i_core_int_sreg[2]
port 42 nsew signal output
rlabel metal2 s 17696 0 17752 400 6 c0_i_core_int_sreg[3]
port 43 nsew signal output
rlabel metal2 s 20384 0 20440 400 6 c0_i_core_int_sreg[4]
port 44 nsew signal output
rlabel metal2 s 23072 0 23128 400 6 c0_i_core_int_sreg[5]
port 45 nsew signal output
rlabel metal2 s 25760 0 25816 400 6 c0_i_core_int_sreg[6]
port 46 nsew signal output
rlabel metal2 s 28448 0 28504 400 6 c0_i_core_int_sreg[7]
port 47 nsew signal output
rlabel metal2 s 31136 0 31192 400 6 c0_i_core_int_sreg[8]
port 48 nsew signal output
rlabel metal2 s 33376 0 33432 400 6 c0_i_core_int_sreg[9]
port 49 nsew signal output
rlabel metal2 s 5152 0 5208 400 6 c0_i_irq
port 50 nsew signal output
rlabel metal2 s 5376 0 5432 400 6 c0_i_mc_core_int
port 51 nsew signal output
rlabel metal2 s 5600 0 5656 400 6 c0_i_mem_ack
port 52 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 c0_i_mem_data[0]
port 53 nsew signal output
rlabel metal2 s 35840 0 35896 400 6 c0_i_mem_data[10]
port 54 nsew signal output
rlabel metal2 s 38080 0 38136 400 6 c0_i_mem_data[11]
port 55 nsew signal output
rlabel metal2 s 40320 0 40376 400 6 c0_i_mem_data[12]
port 56 nsew signal output
rlabel metal2 s 42560 0 42616 400 6 c0_i_mem_data[13]
port 57 nsew signal output
rlabel metal2 s 44800 0 44856 400 6 c0_i_mem_data[14]
port 58 nsew signal output
rlabel metal2 s 47040 0 47096 400 6 c0_i_mem_data[15]
port 59 nsew signal output
rlabel metal2 s 12320 0 12376 400 6 c0_i_mem_data[1]
port 60 nsew signal output
rlabel metal2 s 15232 0 15288 400 6 c0_i_mem_data[2]
port 61 nsew signal output
rlabel metal2 s 17920 0 17976 400 6 c0_i_mem_data[3]
port 62 nsew signal output
rlabel metal2 s 20608 0 20664 400 6 c0_i_mem_data[4]
port 63 nsew signal output
rlabel metal2 s 23296 0 23352 400 6 c0_i_mem_data[5]
port 64 nsew signal output
rlabel metal2 s 25984 0 26040 400 6 c0_i_mem_data[6]
port 65 nsew signal output
rlabel metal2 s 28672 0 28728 400 6 c0_i_mem_data[7]
port 66 nsew signal output
rlabel metal2 s 31360 0 31416 400 6 c0_i_mem_data[8]
port 67 nsew signal output
rlabel metal2 s 33600 0 33656 400 6 c0_i_mem_data[9]
port 68 nsew signal output
rlabel metal2 s 5824 0 5880 400 6 c0_i_mem_exception
port 69 nsew signal output
rlabel metal2 s 9632 0 9688 400 6 c0_i_req_data[0]
port 70 nsew signal output
rlabel metal2 s 36064 0 36120 400 6 c0_i_req_data[10]
port 71 nsew signal output
rlabel metal2 s 38304 0 38360 400 6 c0_i_req_data[11]
port 72 nsew signal output
rlabel metal2 s 40544 0 40600 400 6 c0_i_req_data[12]
port 73 nsew signal output
rlabel metal2 s 42784 0 42840 400 6 c0_i_req_data[13]
port 74 nsew signal output
rlabel metal2 s 45024 0 45080 400 6 c0_i_req_data[14]
port 75 nsew signal output
rlabel metal2 s 47264 0 47320 400 6 c0_i_req_data[15]
port 76 nsew signal output
rlabel metal2 s 48608 0 48664 400 6 c0_i_req_data[16]
port 77 nsew signal output
rlabel metal2 s 48832 0 48888 400 6 c0_i_req_data[17]
port 78 nsew signal output
rlabel metal2 s 49056 0 49112 400 6 c0_i_req_data[18]
port 79 nsew signal output
rlabel metal2 s 49280 0 49336 400 6 c0_i_req_data[19]
port 80 nsew signal output
rlabel metal2 s 12544 0 12600 400 6 c0_i_req_data[1]
port 81 nsew signal output
rlabel metal2 s 49504 0 49560 400 6 c0_i_req_data[20]
port 82 nsew signal output
rlabel metal2 s 49728 0 49784 400 6 c0_i_req_data[21]
port 83 nsew signal output
rlabel metal2 s 49952 0 50008 400 6 c0_i_req_data[22]
port 84 nsew signal output
rlabel metal2 s 50176 0 50232 400 6 c0_i_req_data[23]
port 85 nsew signal output
rlabel metal2 s 50400 0 50456 400 6 c0_i_req_data[24]
port 86 nsew signal output
rlabel metal2 s 50624 0 50680 400 6 c0_i_req_data[25]
port 87 nsew signal output
rlabel metal2 s 50848 0 50904 400 6 c0_i_req_data[26]
port 88 nsew signal output
rlabel metal2 s 51072 0 51128 400 6 c0_i_req_data[27]
port 89 nsew signal output
rlabel metal2 s 51296 0 51352 400 6 c0_i_req_data[28]
port 90 nsew signal output
rlabel metal2 s 51520 0 51576 400 6 c0_i_req_data[29]
port 91 nsew signal output
rlabel metal2 s 15456 0 15512 400 6 c0_i_req_data[2]
port 92 nsew signal output
rlabel metal2 s 51744 0 51800 400 6 c0_i_req_data[30]
port 93 nsew signal output
rlabel metal2 s 51968 0 52024 400 6 c0_i_req_data[31]
port 94 nsew signal output
rlabel metal2 s 18144 0 18200 400 6 c0_i_req_data[3]
port 95 nsew signal output
rlabel metal2 s 20832 0 20888 400 6 c0_i_req_data[4]
port 96 nsew signal output
rlabel metal2 s 23520 0 23576 400 6 c0_i_req_data[5]
port 97 nsew signal output
rlabel metal2 s 26208 0 26264 400 6 c0_i_req_data[6]
port 98 nsew signal output
rlabel metal2 s 28896 0 28952 400 6 c0_i_req_data[7]
port 99 nsew signal output
rlabel metal2 s 31584 0 31640 400 6 c0_i_req_data[8]
port 100 nsew signal output
rlabel metal2 s 33824 0 33880 400 6 c0_i_req_data[9]
port 101 nsew signal output
rlabel metal2 s 6048 0 6104 400 6 c0_i_req_data_valid
port 102 nsew signal output
rlabel metal2 s 6272 0 6328 400 6 c0_o_c_data_page
port 103 nsew signal input
rlabel metal2 s 6496 0 6552 400 6 c0_o_c_instr_long
port 104 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 c0_o_c_instr_page
port 105 nsew signal input
rlabel metal2 s 6944 0 7000 400 6 c0_o_icache_flush
port 106 nsew signal input
rlabel metal2 s 9856 0 9912 400 6 c0_o_instr_long_addr[0]
port 107 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 c0_o_instr_long_addr[1]
port 108 nsew signal input
rlabel metal2 s 15680 0 15736 400 6 c0_o_instr_long_addr[2]
port 109 nsew signal input
rlabel metal2 s 18368 0 18424 400 6 c0_o_instr_long_addr[3]
port 110 nsew signal input
rlabel metal2 s 21056 0 21112 400 6 c0_o_instr_long_addr[4]
port 111 nsew signal input
rlabel metal2 s 23744 0 23800 400 6 c0_o_instr_long_addr[5]
port 112 nsew signal input
rlabel metal2 s 26432 0 26488 400 6 c0_o_instr_long_addr[6]
port 113 nsew signal input
rlabel metal2 s 29120 0 29176 400 6 c0_o_instr_long_addr[7]
port 114 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 c0_o_mem_addr[0]
port 115 nsew signal input
rlabel metal2 s 36288 0 36344 400 6 c0_o_mem_addr[10]
port 116 nsew signal input
rlabel metal2 s 38528 0 38584 400 6 c0_o_mem_addr[11]
port 117 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 c0_o_mem_addr[12]
port 118 nsew signal input
rlabel metal2 s 43008 0 43064 400 6 c0_o_mem_addr[13]
port 119 nsew signal input
rlabel metal2 s 45248 0 45304 400 6 c0_o_mem_addr[14]
port 120 nsew signal input
rlabel metal2 s 47488 0 47544 400 6 c0_o_mem_addr[15]
port 121 nsew signal input
rlabel metal2 s 12992 0 13048 400 6 c0_o_mem_addr[1]
port 122 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 c0_o_mem_addr[2]
port 123 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 c0_o_mem_addr[3]
port 124 nsew signal input
rlabel metal2 s 21280 0 21336 400 6 c0_o_mem_addr[4]
port 125 nsew signal input
rlabel metal2 s 23968 0 24024 400 6 c0_o_mem_addr[5]
port 126 nsew signal input
rlabel metal2 s 26656 0 26712 400 6 c0_o_mem_addr[6]
port 127 nsew signal input
rlabel metal2 s 29344 0 29400 400 6 c0_o_mem_addr[7]
port 128 nsew signal input
rlabel metal2 s 31808 0 31864 400 6 c0_o_mem_addr[8]
port 129 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 c0_o_mem_addr[9]
port 130 nsew signal input
rlabel metal2 s 10304 0 10360 400 6 c0_o_mem_data[0]
port 131 nsew signal input
rlabel metal2 s 36512 0 36568 400 6 c0_o_mem_data[10]
port 132 nsew signal input
rlabel metal2 s 38752 0 38808 400 6 c0_o_mem_data[11]
port 133 nsew signal input
rlabel metal2 s 40992 0 41048 400 6 c0_o_mem_data[12]
port 134 nsew signal input
rlabel metal2 s 43232 0 43288 400 6 c0_o_mem_data[13]
port 135 nsew signal input
rlabel metal2 s 45472 0 45528 400 6 c0_o_mem_data[14]
port 136 nsew signal input
rlabel metal2 s 47712 0 47768 400 6 c0_o_mem_data[15]
port 137 nsew signal input
rlabel metal2 s 13216 0 13272 400 6 c0_o_mem_data[1]
port 138 nsew signal input
rlabel metal2 s 16128 0 16184 400 6 c0_o_mem_data[2]
port 139 nsew signal input
rlabel metal2 s 18816 0 18872 400 6 c0_o_mem_data[3]
port 140 nsew signal input
rlabel metal2 s 21504 0 21560 400 6 c0_o_mem_data[4]
port 141 nsew signal input
rlabel metal2 s 24192 0 24248 400 6 c0_o_mem_data[5]
port 142 nsew signal input
rlabel metal2 s 26880 0 26936 400 6 c0_o_mem_data[6]
port 143 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 c0_o_mem_data[7]
port 144 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 c0_o_mem_data[8]
port 145 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 c0_o_mem_data[9]
port 146 nsew signal input
rlabel metal2 s 10528 0 10584 400 6 c0_o_mem_high_addr[0]
port 147 nsew signal input
rlabel metal2 s 13440 0 13496 400 6 c0_o_mem_high_addr[1]
port 148 nsew signal input
rlabel metal2 s 16352 0 16408 400 6 c0_o_mem_high_addr[2]
port 149 nsew signal input
rlabel metal2 s 19040 0 19096 400 6 c0_o_mem_high_addr[3]
port 150 nsew signal input
rlabel metal2 s 21728 0 21784 400 6 c0_o_mem_high_addr[4]
port 151 nsew signal input
rlabel metal2 s 24416 0 24472 400 6 c0_o_mem_high_addr[5]
port 152 nsew signal input
rlabel metal2 s 27104 0 27160 400 6 c0_o_mem_high_addr[6]
port 153 nsew signal input
rlabel metal2 s 29792 0 29848 400 6 c0_o_mem_high_addr[7]
port 154 nsew signal input
rlabel metal2 s 7168 0 7224 400 6 c0_o_mem_long_mode
port 155 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 c0_o_mem_req
port 156 nsew signal input
rlabel metal2 s 10752 0 10808 400 6 c0_o_mem_sel[0]
port 157 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 c0_o_mem_sel[1]
port 158 nsew signal input
rlabel metal2 s 7616 0 7672 400 6 c0_o_mem_we
port 159 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 c0_o_req_active
port 160 nsew signal input
rlabel metal2 s 10976 0 11032 400 6 c0_o_req_addr[0]
port 161 nsew signal input
rlabel metal2 s 36736 0 36792 400 6 c0_o_req_addr[10]
port 162 nsew signal input
rlabel metal2 s 38976 0 39032 400 6 c0_o_req_addr[11]
port 163 nsew signal input
rlabel metal2 s 41216 0 41272 400 6 c0_o_req_addr[12]
port 164 nsew signal input
rlabel metal2 s 43456 0 43512 400 6 c0_o_req_addr[13]
port 165 nsew signal input
rlabel metal2 s 45696 0 45752 400 6 c0_o_req_addr[14]
port 166 nsew signal input
rlabel metal2 s 47936 0 47992 400 6 c0_o_req_addr[15]
port 167 nsew signal input
rlabel metal2 s 13888 0 13944 400 6 c0_o_req_addr[1]
port 168 nsew signal input
rlabel metal2 s 16576 0 16632 400 6 c0_o_req_addr[2]
port 169 nsew signal input
rlabel metal2 s 19264 0 19320 400 6 c0_o_req_addr[3]
port 170 nsew signal input
rlabel metal2 s 21952 0 22008 400 6 c0_o_req_addr[4]
port 171 nsew signal input
rlabel metal2 s 24640 0 24696 400 6 c0_o_req_addr[5]
port 172 nsew signal input
rlabel metal2 s 27328 0 27384 400 6 c0_o_req_addr[6]
port 173 nsew signal input
rlabel metal2 s 30016 0 30072 400 6 c0_o_req_addr[7]
port 174 nsew signal input
rlabel metal2 s 32256 0 32312 400 6 c0_o_req_addr[8]
port 175 nsew signal input
rlabel metal2 s 34496 0 34552 400 6 c0_o_req_addr[9]
port 176 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 c0_o_req_ppl_submit
port 177 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 c0_rst
port 178 nsew signal output
rlabel metal2 s 11200 0 11256 400 6 c0_sr_bus_addr[0]
port 179 nsew signal input
rlabel metal2 s 36960 0 37016 400 6 c0_sr_bus_addr[10]
port 180 nsew signal input
rlabel metal2 s 39200 0 39256 400 6 c0_sr_bus_addr[11]
port 181 nsew signal input
rlabel metal2 s 41440 0 41496 400 6 c0_sr_bus_addr[12]
port 182 nsew signal input
rlabel metal2 s 43680 0 43736 400 6 c0_sr_bus_addr[13]
port 183 nsew signal input
rlabel metal2 s 45920 0 45976 400 6 c0_sr_bus_addr[14]
port 184 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 c0_sr_bus_addr[15]
port 185 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 c0_sr_bus_addr[1]
port 186 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 c0_sr_bus_addr[2]
port 187 nsew signal input
rlabel metal2 s 19488 0 19544 400 6 c0_sr_bus_addr[3]
port 188 nsew signal input
rlabel metal2 s 22176 0 22232 400 6 c0_sr_bus_addr[4]
port 189 nsew signal input
rlabel metal2 s 24864 0 24920 400 6 c0_sr_bus_addr[5]
port 190 nsew signal input
rlabel metal2 s 27552 0 27608 400 6 c0_sr_bus_addr[6]
port 191 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 c0_sr_bus_addr[7]
port 192 nsew signal input
rlabel metal2 s 32480 0 32536 400 6 c0_sr_bus_addr[8]
port 193 nsew signal input
rlabel metal2 s 34720 0 34776 400 6 c0_sr_bus_addr[9]
port 194 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 c0_sr_bus_data_o[0]
port 195 nsew signal input
rlabel metal2 s 37184 0 37240 400 6 c0_sr_bus_data_o[10]
port 196 nsew signal input
rlabel metal2 s 39424 0 39480 400 6 c0_sr_bus_data_o[11]
port 197 nsew signal input
rlabel metal2 s 41664 0 41720 400 6 c0_sr_bus_data_o[12]
port 198 nsew signal input
rlabel metal2 s 43904 0 43960 400 6 c0_sr_bus_data_o[13]
port 199 nsew signal input
rlabel metal2 s 46144 0 46200 400 6 c0_sr_bus_data_o[14]
port 200 nsew signal input
rlabel metal2 s 48384 0 48440 400 6 c0_sr_bus_data_o[15]
port 201 nsew signal input
rlabel metal2 s 14336 0 14392 400 6 c0_sr_bus_data_o[1]
port 202 nsew signal input
rlabel metal2 s 17024 0 17080 400 6 c0_sr_bus_data_o[2]
port 203 nsew signal input
rlabel metal2 s 19712 0 19768 400 6 c0_sr_bus_data_o[3]
port 204 nsew signal input
rlabel metal2 s 22400 0 22456 400 6 c0_sr_bus_data_o[4]
port 205 nsew signal input
rlabel metal2 s 25088 0 25144 400 6 c0_sr_bus_data_o[5]
port 206 nsew signal input
rlabel metal2 s 27776 0 27832 400 6 c0_sr_bus_data_o[6]
port 207 nsew signal input
rlabel metal2 s 30464 0 30520 400 6 c0_sr_bus_data_o[7]
port 208 nsew signal input
rlabel metal2 s 32704 0 32760 400 6 c0_sr_bus_data_o[8]
port 209 nsew signal input
rlabel metal2 s 34944 0 35000 400 6 c0_sr_bus_data_o[9]
port 210 nsew signal input
rlabel metal2 s 8512 0 8568 400 6 c0_sr_bus_we
port 211 nsew signal input
rlabel metal2 s 71680 0 71736 400 6 c1_dbg_pc[0]
port 212 nsew signal input
rlabel metal2 s 98112 0 98168 400 6 c1_dbg_pc[10]
port 213 nsew signal input
rlabel metal2 s 100352 0 100408 400 6 c1_dbg_pc[11]
port 214 nsew signal input
rlabel metal2 s 102592 0 102648 400 6 c1_dbg_pc[12]
port 215 nsew signal input
rlabel metal2 s 104832 0 104888 400 6 c1_dbg_pc[13]
port 216 nsew signal input
rlabel metal2 s 107072 0 107128 400 6 c1_dbg_pc[14]
port 217 nsew signal input
rlabel metal2 s 109312 0 109368 400 6 c1_dbg_pc[15]
port 218 nsew signal input
rlabel metal2 s 74592 0 74648 400 6 c1_dbg_pc[1]
port 219 nsew signal input
rlabel metal2 s 77504 0 77560 400 6 c1_dbg_pc[2]
port 220 nsew signal input
rlabel metal2 s 80192 0 80248 400 6 c1_dbg_pc[3]
port 221 nsew signal input
rlabel metal2 s 82880 0 82936 400 6 c1_dbg_pc[4]
port 222 nsew signal input
rlabel metal2 s 85568 0 85624 400 6 c1_dbg_pc[5]
port 223 nsew signal input
rlabel metal2 s 88256 0 88312 400 6 c1_dbg_pc[6]
port 224 nsew signal input
rlabel metal2 s 90944 0 91000 400 6 c1_dbg_pc[7]
port 225 nsew signal input
rlabel metal2 s 93632 0 93688 400 6 c1_dbg_pc[8]
port 226 nsew signal input
rlabel metal2 s 95872 0 95928 400 6 c1_dbg_pc[9]
port 227 nsew signal input
rlabel metal2 s 71904 0 71960 400 6 c1_dbg_r0[0]
port 228 nsew signal input
rlabel metal2 s 98336 0 98392 400 6 c1_dbg_r0[10]
port 229 nsew signal input
rlabel metal2 s 100576 0 100632 400 6 c1_dbg_r0[11]
port 230 nsew signal input
rlabel metal2 s 102816 0 102872 400 6 c1_dbg_r0[12]
port 231 nsew signal input
rlabel metal2 s 105056 0 105112 400 6 c1_dbg_r0[13]
port 232 nsew signal input
rlabel metal2 s 107296 0 107352 400 6 c1_dbg_r0[14]
port 233 nsew signal input
rlabel metal2 s 109536 0 109592 400 6 c1_dbg_r0[15]
port 234 nsew signal input
rlabel metal2 s 74816 0 74872 400 6 c1_dbg_r0[1]
port 235 nsew signal input
rlabel metal2 s 77728 0 77784 400 6 c1_dbg_r0[2]
port 236 nsew signal input
rlabel metal2 s 80416 0 80472 400 6 c1_dbg_r0[3]
port 237 nsew signal input
rlabel metal2 s 83104 0 83160 400 6 c1_dbg_r0[4]
port 238 nsew signal input
rlabel metal2 s 85792 0 85848 400 6 c1_dbg_r0[5]
port 239 nsew signal input
rlabel metal2 s 88480 0 88536 400 6 c1_dbg_r0[6]
port 240 nsew signal input
rlabel metal2 s 91168 0 91224 400 6 c1_dbg_r0[7]
port 241 nsew signal input
rlabel metal2 s 93856 0 93912 400 6 c1_dbg_r0[8]
port 242 nsew signal input
rlabel metal2 s 96096 0 96152 400 6 c1_dbg_r0[9]
port 243 nsew signal input
rlabel metal2 s 67872 0 67928 400 6 c1_disable
port 244 nsew signal output
rlabel metal2 s 72128 0 72184 400 6 c1_i_core_int_sreg[0]
port 245 nsew signal output
rlabel metal2 s 98560 0 98616 400 6 c1_i_core_int_sreg[10]
port 246 nsew signal output
rlabel metal2 s 100800 0 100856 400 6 c1_i_core_int_sreg[11]
port 247 nsew signal output
rlabel metal2 s 103040 0 103096 400 6 c1_i_core_int_sreg[12]
port 248 nsew signal output
rlabel metal2 s 105280 0 105336 400 6 c1_i_core_int_sreg[13]
port 249 nsew signal output
rlabel metal2 s 107520 0 107576 400 6 c1_i_core_int_sreg[14]
port 250 nsew signal output
rlabel metal2 s 109760 0 109816 400 6 c1_i_core_int_sreg[15]
port 251 nsew signal output
rlabel metal2 s 75040 0 75096 400 6 c1_i_core_int_sreg[1]
port 252 nsew signal output
rlabel metal2 s 77952 0 78008 400 6 c1_i_core_int_sreg[2]
port 253 nsew signal output
rlabel metal2 s 80640 0 80696 400 6 c1_i_core_int_sreg[3]
port 254 nsew signal output
rlabel metal2 s 83328 0 83384 400 6 c1_i_core_int_sreg[4]
port 255 nsew signal output
rlabel metal2 s 86016 0 86072 400 6 c1_i_core_int_sreg[5]
port 256 nsew signal output
rlabel metal2 s 88704 0 88760 400 6 c1_i_core_int_sreg[6]
port 257 nsew signal output
rlabel metal2 s 91392 0 91448 400 6 c1_i_core_int_sreg[7]
port 258 nsew signal output
rlabel metal2 s 94080 0 94136 400 6 c1_i_core_int_sreg[8]
port 259 nsew signal output
rlabel metal2 s 96320 0 96376 400 6 c1_i_core_int_sreg[9]
port 260 nsew signal output
rlabel metal2 s 68096 0 68152 400 6 c1_i_irq
port 261 nsew signal output
rlabel metal2 s 68320 0 68376 400 6 c1_i_mc_core_int
port 262 nsew signal output
rlabel metal2 s 68544 0 68600 400 6 c1_i_mem_ack
port 263 nsew signal output
rlabel metal2 s 72352 0 72408 400 6 c1_i_mem_data[0]
port 264 nsew signal output
rlabel metal2 s 98784 0 98840 400 6 c1_i_mem_data[10]
port 265 nsew signal output
rlabel metal2 s 101024 0 101080 400 6 c1_i_mem_data[11]
port 266 nsew signal output
rlabel metal2 s 103264 0 103320 400 6 c1_i_mem_data[12]
port 267 nsew signal output
rlabel metal2 s 105504 0 105560 400 6 c1_i_mem_data[13]
port 268 nsew signal output
rlabel metal2 s 107744 0 107800 400 6 c1_i_mem_data[14]
port 269 nsew signal output
rlabel metal2 s 109984 0 110040 400 6 c1_i_mem_data[15]
port 270 nsew signal output
rlabel metal2 s 75264 0 75320 400 6 c1_i_mem_data[1]
port 271 nsew signal output
rlabel metal2 s 78176 0 78232 400 6 c1_i_mem_data[2]
port 272 nsew signal output
rlabel metal2 s 80864 0 80920 400 6 c1_i_mem_data[3]
port 273 nsew signal output
rlabel metal2 s 83552 0 83608 400 6 c1_i_mem_data[4]
port 274 nsew signal output
rlabel metal2 s 86240 0 86296 400 6 c1_i_mem_data[5]
port 275 nsew signal output
rlabel metal2 s 88928 0 88984 400 6 c1_i_mem_data[6]
port 276 nsew signal output
rlabel metal2 s 91616 0 91672 400 6 c1_i_mem_data[7]
port 277 nsew signal output
rlabel metal2 s 94304 0 94360 400 6 c1_i_mem_data[8]
port 278 nsew signal output
rlabel metal2 s 96544 0 96600 400 6 c1_i_mem_data[9]
port 279 nsew signal output
rlabel metal2 s 68768 0 68824 400 6 c1_i_mem_exception
port 280 nsew signal output
rlabel metal2 s 72576 0 72632 400 6 c1_i_req_data[0]
port 281 nsew signal output
rlabel metal2 s 99008 0 99064 400 6 c1_i_req_data[10]
port 282 nsew signal output
rlabel metal2 s 101248 0 101304 400 6 c1_i_req_data[11]
port 283 nsew signal output
rlabel metal2 s 103488 0 103544 400 6 c1_i_req_data[12]
port 284 nsew signal output
rlabel metal2 s 105728 0 105784 400 6 c1_i_req_data[13]
port 285 nsew signal output
rlabel metal2 s 107968 0 108024 400 6 c1_i_req_data[14]
port 286 nsew signal output
rlabel metal2 s 110208 0 110264 400 6 c1_i_req_data[15]
port 287 nsew signal output
rlabel metal2 s 111552 0 111608 400 6 c1_i_req_data[16]
port 288 nsew signal output
rlabel metal2 s 111776 0 111832 400 6 c1_i_req_data[17]
port 289 nsew signal output
rlabel metal2 s 112000 0 112056 400 6 c1_i_req_data[18]
port 290 nsew signal output
rlabel metal2 s 112224 0 112280 400 6 c1_i_req_data[19]
port 291 nsew signal output
rlabel metal2 s 75488 0 75544 400 6 c1_i_req_data[1]
port 292 nsew signal output
rlabel metal2 s 112448 0 112504 400 6 c1_i_req_data[20]
port 293 nsew signal output
rlabel metal2 s 112672 0 112728 400 6 c1_i_req_data[21]
port 294 nsew signal output
rlabel metal2 s 112896 0 112952 400 6 c1_i_req_data[22]
port 295 nsew signal output
rlabel metal2 s 113120 0 113176 400 6 c1_i_req_data[23]
port 296 nsew signal output
rlabel metal2 s 113344 0 113400 400 6 c1_i_req_data[24]
port 297 nsew signal output
rlabel metal2 s 113568 0 113624 400 6 c1_i_req_data[25]
port 298 nsew signal output
rlabel metal2 s 113792 0 113848 400 6 c1_i_req_data[26]
port 299 nsew signal output
rlabel metal2 s 114016 0 114072 400 6 c1_i_req_data[27]
port 300 nsew signal output
rlabel metal2 s 114240 0 114296 400 6 c1_i_req_data[28]
port 301 nsew signal output
rlabel metal2 s 114464 0 114520 400 6 c1_i_req_data[29]
port 302 nsew signal output
rlabel metal2 s 78400 0 78456 400 6 c1_i_req_data[2]
port 303 nsew signal output
rlabel metal2 s 114688 0 114744 400 6 c1_i_req_data[30]
port 304 nsew signal output
rlabel metal2 s 114912 0 114968 400 6 c1_i_req_data[31]
port 305 nsew signal output
rlabel metal2 s 81088 0 81144 400 6 c1_i_req_data[3]
port 306 nsew signal output
rlabel metal2 s 83776 0 83832 400 6 c1_i_req_data[4]
port 307 nsew signal output
rlabel metal2 s 86464 0 86520 400 6 c1_i_req_data[5]
port 308 nsew signal output
rlabel metal2 s 89152 0 89208 400 6 c1_i_req_data[6]
port 309 nsew signal output
rlabel metal2 s 91840 0 91896 400 6 c1_i_req_data[7]
port 310 nsew signal output
rlabel metal2 s 94528 0 94584 400 6 c1_i_req_data[8]
port 311 nsew signal output
rlabel metal2 s 96768 0 96824 400 6 c1_i_req_data[9]
port 312 nsew signal output
rlabel metal2 s 68992 0 69048 400 6 c1_i_req_data_valid
port 313 nsew signal output
rlabel metal2 s 69216 0 69272 400 6 c1_o_c_data_page
port 314 nsew signal input
rlabel metal2 s 69440 0 69496 400 6 c1_o_c_instr_long
port 315 nsew signal input
rlabel metal2 s 69664 0 69720 400 6 c1_o_c_instr_page
port 316 nsew signal input
rlabel metal2 s 69888 0 69944 400 6 c1_o_icache_flush
port 317 nsew signal input
rlabel metal2 s 72800 0 72856 400 6 c1_o_instr_long_addr[0]
port 318 nsew signal input
rlabel metal2 s 75712 0 75768 400 6 c1_o_instr_long_addr[1]
port 319 nsew signal input
rlabel metal2 s 78624 0 78680 400 6 c1_o_instr_long_addr[2]
port 320 nsew signal input
rlabel metal2 s 81312 0 81368 400 6 c1_o_instr_long_addr[3]
port 321 nsew signal input
rlabel metal2 s 84000 0 84056 400 6 c1_o_instr_long_addr[4]
port 322 nsew signal input
rlabel metal2 s 86688 0 86744 400 6 c1_o_instr_long_addr[5]
port 323 nsew signal input
rlabel metal2 s 89376 0 89432 400 6 c1_o_instr_long_addr[6]
port 324 nsew signal input
rlabel metal2 s 92064 0 92120 400 6 c1_o_instr_long_addr[7]
port 325 nsew signal input
rlabel metal2 s 73024 0 73080 400 6 c1_o_mem_addr[0]
port 326 nsew signal input
rlabel metal2 s 99232 0 99288 400 6 c1_o_mem_addr[10]
port 327 nsew signal input
rlabel metal2 s 101472 0 101528 400 6 c1_o_mem_addr[11]
port 328 nsew signal input
rlabel metal2 s 103712 0 103768 400 6 c1_o_mem_addr[12]
port 329 nsew signal input
rlabel metal2 s 105952 0 106008 400 6 c1_o_mem_addr[13]
port 330 nsew signal input
rlabel metal2 s 108192 0 108248 400 6 c1_o_mem_addr[14]
port 331 nsew signal input
rlabel metal2 s 110432 0 110488 400 6 c1_o_mem_addr[15]
port 332 nsew signal input
rlabel metal2 s 75936 0 75992 400 6 c1_o_mem_addr[1]
port 333 nsew signal input
rlabel metal2 s 78848 0 78904 400 6 c1_o_mem_addr[2]
port 334 nsew signal input
rlabel metal2 s 81536 0 81592 400 6 c1_o_mem_addr[3]
port 335 nsew signal input
rlabel metal2 s 84224 0 84280 400 6 c1_o_mem_addr[4]
port 336 nsew signal input
rlabel metal2 s 86912 0 86968 400 6 c1_o_mem_addr[5]
port 337 nsew signal input
rlabel metal2 s 89600 0 89656 400 6 c1_o_mem_addr[6]
port 338 nsew signal input
rlabel metal2 s 92288 0 92344 400 6 c1_o_mem_addr[7]
port 339 nsew signal input
rlabel metal2 s 94752 0 94808 400 6 c1_o_mem_addr[8]
port 340 nsew signal input
rlabel metal2 s 96992 0 97048 400 6 c1_o_mem_addr[9]
port 341 nsew signal input
rlabel metal2 s 73248 0 73304 400 6 c1_o_mem_data[0]
port 342 nsew signal input
rlabel metal2 s 99456 0 99512 400 6 c1_o_mem_data[10]
port 343 nsew signal input
rlabel metal2 s 101696 0 101752 400 6 c1_o_mem_data[11]
port 344 nsew signal input
rlabel metal2 s 103936 0 103992 400 6 c1_o_mem_data[12]
port 345 nsew signal input
rlabel metal2 s 106176 0 106232 400 6 c1_o_mem_data[13]
port 346 nsew signal input
rlabel metal2 s 108416 0 108472 400 6 c1_o_mem_data[14]
port 347 nsew signal input
rlabel metal2 s 110656 0 110712 400 6 c1_o_mem_data[15]
port 348 nsew signal input
rlabel metal2 s 76160 0 76216 400 6 c1_o_mem_data[1]
port 349 nsew signal input
rlabel metal2 s 79072 0 79128 400 6 c1_o_mem_data[2]
port 350 nsew signal input
rlabel metal2 s 81760 0 81816 400 6 c1_o_mem_data[3]
port 351 nsew signal input
rlabel metal2 s 84448 0 84504 400 6 c1_o_mem_data[4]
port 352 nsew signal input
rlabel metal2 s 87136 0 87192 400 6 c1_o_mem_data[5]
port 353 nsew signal input
rlabel metal2 s 89824 0 89880 400 6 c1_o_mem_data[6]
port 354 nsew signal input
rlabel metal2 s 92512 0 92568 400 6 c1_o_mem_data[7]
port 355 nsew signal input
rlabel metal2 s 94976 0 95032 400 6 c1_o_mem_data[8]
port 356 nsew signal input
rlabel metal2 s 97216 0 97272 400 6 c1_o_mem_data[9]
port 357 nsew signal input
rlabel metal2 s 73472 0 73528 400 6 c1_o_mem_high_addr[0]
port 358 nsew signal input
rlabel metal2 s 76384 0 76440 400 6 c1_o_mem_high_addr[1]
port 359 nsew signal input
rlabel metal2 s 79296 0 79352 400 6 c1_o_mem_high_addr[2]
port 360 nsew signal input
rlabel metal2 s 81984 0 82040 400 6 c1_o_mem_high_addr[3]
port 361 nsew signal input
rlabel metal2 s 84672 0 84728 400 6 c1_o_mem_high_addr[4]
port 362 nsew signal input
rlabel metal2 s 87360 0 87416 400 6 c1_o_mem_high_addr[5]
port 363 nsew signal input
rlabel metal2 s 90048 0 90104 400 6 c1_o_mem_high_addr[6]
port 364 nsew signal input
rlabel metal2 s 92736 0 92792 400 6 c1_o_mem_high_addr[7]
port 365 nsew signal input
rlabel metal2 s 70112 0 70168 400 6 c1_o_mem_long_mode
port 366 nsew signal input
rlabel metal2 s 70336 0 70392 400 6 c1_o_mem_req
port 367 nsew signal input
rlabel metal2 s 73696 0 73752 400 6 c1_o_mem_sel[0]
port 368 nsew signal input
rlabel metal2 s 76608 0 76664 400 6 c1_o_mem_sel[1]
port 369 nsew signal input
rlabel metal2 s 70560 0 70616 400 6 c1_o_mem_we
port 370 nsew signal input
rlabel metal2 s 70784 0 70840 400 6 c1_o_req_active
port 371 nsew signal input
rlabel metal2 s 73920 0 73976 400 6 c1_o_req_addr[0]
port 372 nsew signal input
rlabel metal2 s 99680 0 99736 400 6 c1_o_req_addr[10]
port 373 nsew signal input
rlabel metal2 s 101920 0 101976 400 6 c1_o_req_addr[11]
port 374 nsew signal input
rlabel metal2 s 104160 0 104216 400 6 c1_o_req_addr[12]
port 375 nsew signal input
rlabel metal2 s 106400 0 106456 400 6 c1_o_req_addr[13]
port 376 nsew signal input
rlabel metal2 s 108640 0 108696 400 6 c1_o_req_addr[14]
port 377 nsew signal input
rlabel metal2 s 110880 0 110936 400 6 c1_o_req_addr[15]
port 378 nsew signal input
rlabel metal2 s 76832 0 76888 400 6 c1_o_req_addr[1]
port 379 nsew signal input
rlabel metal2 s 79520 0 79576 400 6 c1_o_req_addr[2]
port 380 nsew signal input
rlabel metal2 s 82208 0 82264 400 6 c1_o_req_addr[3]
port 381 nsew signal input
rlabel metal2 s 84896 0 84952 400 6 c1_o_req_addr[4]
port 382 nsew signal input
rlabel metal2 s 87584 0 87640 400 6 c1_o_req_addr[5]
port 383 nsew signal input
rlabel metal2 s 90272 0 90328 400 6 c1_o_req_addr[6]
port 384 nsew signal input
rlabel metal2 s 92960 0 93016 400 6 c1_o_req_addr[7]
port 385 nsew signal input
rlabel metal2 s 95200 0 95256 400 6 c1_o_req_addr[8]
port 386 nsew signal input
rlabel metal2 s 97440 0 97496 400 6 c1_o_req_addr[9]
port 387 nsew signal input
rlabel metal2 s 71008 0 71064 400 6 c1_o_req_ppl_submit
port 388 nsew signal input
rlabel metal2 s 71232 0 71288 400 6 c1_rst
port 389 nsew signal output
rlabel metal2 s 74144 0 74200 400 6 c1_sr_bus_addr[0]
port 390 nsew signal input
rlabel metal2 s 99904 0 99960 400 6 c1_sr_bus_addr[10]
port 391 nsew signal input
rlabel metal2 s 102144 0 102200 400 6 c1_sr_bus_addr[11]
port 392 nsew signal input
rlabel metal2 s 104384 0 104440 400 6 c1_sr_bus_addr[12]
port 393 nsew signal input
rlabel metal2 s 106624 0 106680 400 6 c1_sr_bus_addr[13]
port 394 nsew signal input
rlabel metal2 s 108864 0 108920 400 6 c1_sr_bus_addr[14]
port 395 nsew signal input
rlabel metal2 s 111104 0 111160 400 6 c1_sr_bus_addr[15]
port 396 nsew signal input
rlabel metal2 s 77056 0 77112 400 6 c1_sr_bus_addr[1]
port 397 nsew signal input
rlabel metal2 s 79744 0 79800 400 6 c1_sr_bus_addr[2]
port 398 nsew signal input
rlabel metal2 s 82432 0 82488 400 6 c1_sr_bus_addr[3]
port 399 nsew signal input
rlabel metal2 s 85120 0 85176 400 6 c1_sr_bus_addr[4]
port 400 nsew signal input
rlabel metal2 s 87808 0 87864 400 6 c1_sr_bus_addr[5]
port 401 nsew signal input
rlabel metal2 s 90496 0 90552 400 6 c1_sr_bus_addr[6]
port 402 nsew signal input
rlabel metal2 s 93184 0 93240 400 6 c1_sr_bus_addr[7]
port 403 nsew signal input
rlabel metal2 s 95424 0 95480 400 6 c1_sr_bus_addr[8]
port 404 nsew signal input
rlabel metal2 s 97664 0 97720 400 6 c1_sr_bus_addr[9]
port 405 nsew signal input
rlabel metal2 s 74368 0 74424 400 6 c1_sr_bus_data_o[0]
port 406 nsew signal input
rlabel metal2 s 100128 0 100184 400 6 c1_sr_bus_data_o[10]
port 407 nsew signal input
rlabel metal2 s 102368 0 102424 400 6 c1_sr_bus_data_o[11]
port 408 nsew signal input
rlabel metal2 s 104608 0 104664 400 6 c1_sr_bus_data_o[12]
port 409 nsew signal input
rlabel metal2 s 106848 0 106904 400 6 c1_sr_bus_data_o[13]
port 410 nsew signal input
rlabel metal2 s 109088 0 109144 400 6 c1_sr_bus_data_o[14]
port 411 nsew signal input
rlabel metal2 s 111328 0 111384 400 6 c1_sr_bus_data_o[15]
port 412 nsew signal input
rlabel metal2 s 77280 0 77336 400 6 c1_sr_bus_data_o[1]
port 413 nsew signal input
rlabel metal2 s 79968 0 80024 400 6 c1_sr_bus_data_o[2]
port 414 nsew signal input
rlabel metal2 s 82656 0 82712 400 6 c1_sr_bus_data_o[3]
port 415 nsew signal input
rlabel metal2 s 85344 0 85400 400 6 c1_sr_bus_data_o[4]
port 416 nsew signal input
rlabel metal2 s 88032 0 88088 400 6 c1_sr_bus_data_o[5]
port 417 nsew signal input
rlabel metal2 s 90720 0 90776 400 6 c1_sr_bus_data_o[6]
port 418 nsew signal input
rlabel metal2 s 93408 0 93464 400 6 c1_sr_bus_data_o[7]
port 419 nsew signal input
rlabel metal2 s 95648 0 95704 400 6 c1_sr_bus_data_o[8]
port 420 nsew signal input
rlabel metal2 s 97888 0 97944 400 6 c1_sr_bus_data_o[9]
port 421 nsew signal input
rlabel metal2 s 71456 0 71512 400 6 c1_sr_bus_we
port 422 nsew signal input
rlabel metal2 s 52192 0 52248 400 6 core_clock
port 423 nsew signal input
rlabel metal2 s 52416 0 52472 400 6 core_reset
port 424 nsew signal input
rlabel metal2 s 3024 34600 3080 35000 6 dcache_mem_ack
port 425 nsew signal input
rlabel metal2 s 13776 34600 13832 35000 6 dcache_mem_addr[0]
port 426 nsew signal output
rlabel metal2 s 71120 34600 71176 35000 6 dcache_mem_addr[10]
port 427 nsew signal output
rlabel metal2 s 76496 34600 76552 35000 6 dcache_mem_addr[11]
port 428 nsew signal output
rlabel metal2 s 81872 34600 81928 35000 6 dcache_mem_addr[12]
port 429 nsew signal output
rlabel metal2 s 87248 34600 87304 35000 6 dcache_mem_addr[13]
port 430 nsew signal output
rlabel metal2 s 92624 34600 92680 35000 6 dcache_mem_addr[14]
port 431 nsew signal output
rlabel metal2 s 98000 34600 98056 35000 6 dcache_mem_addr[15]
port 432 nsew signal output
rlabel metal2 s 103376 34600 103432 35000 6 dcache_mem_addr[16]
port 433 nsew signal output
rlabel metal2 s 105168 34600 105224 35000 6 dcache_mem_addr[17]
port 434 nsew signal output
rlabel metal2 s 106960 34600 107016 35000 6 dcache_mem_addr[18]
port 435 nsew signal output
rlabel metal2 s 108752 34600 108808 35000 6 dcache_mem_addr[19]
port 436 nsew signal output
rlabel metal2 s 20944 34600 21000 35000 6 dcache_mem_addr[1]
port 437 nsew signal output
rlabel metal2 s 110544 34600 110600 35000 6 dcache_mem_addr[20]
port 438 nsew signal output
rlabel metal2 s 112336 34600 112392 35000 6 dcache_mem_addr[21]
port 439 nsew signal output
rlabel metal2 s 114128 34600 114184 35000 6 dcache_mem_addr[22]
port 440 nsew signal output
rlabel metal2 s 115920 34600 115976 35000 6 dcache_mem_addr[23]
port 441 nsew signal output
rlabel metal2 s 28112 34600 28168 35000 6 dcache_mem_addr[2]
port 442 nsew signal output
rlabel metal2 s 33488 34600 33544 35000 6 dcache_mem_addr[3]
port 443 nsew signal output
rlabel metal2 s 38864 34600 38920 35000 6 dcache_mem_addr[4]
port 444 nsew signal output
rlabel metal2 s 44240 34600 44296 35000 6 dcache_mem_addr[5]
port 445 nsew signal output
rlabel metal2 s 49616 34600 49672 35000 6 dcache_mem_addr[6]
port 446 nsew signal output
rlabel metal2 s 54992 34600 55048 35000 6 dcache_mem_addr[7]
port 447 nsew signal output
rlabel metal2 s 60368 34600 60424 35000 6 dcache_mem_addr[8]
port 448 nsew signal output
rlabel metal2 s 65744 34600 65800 35000 6 dcache_mem_addr[9]
port 449 nsew signal output
rlabel metal2 s 3920 34600 3976 35000 6 dcache_mem_cache_enable
port 450 nsew signal output
rlabel metal2 s 4816 34600 4872 35000 6 dcache_mem_exception
port 451 nsew signal input
rlabel metal2 s 14672 34600 14728 35000 6 dcache_mem_i_data[0]
port 452 nsew signal output
rlabel metal2 s 72016 34600 72072 35000 6 dcache_mem_i_data[10]
port 453 nsew signal output
rlabel metal2 s 77392 34600 77448 35000 6 dcache_mem_i_data[11]
port 454 nsew signal output
rlabel metal2 s 82768 34600 82824 35000 6 dcache_mem_i_data[12]
port 455 nsew signal output
rlabel metal2 s 88144 34600 88200 35000 6 dcache_mem_i_data[13]
port 456 nsew signal output
rlabel metal2 s 93520 34600 93576 35000 6 dcache_mem_i_data[14]
port 457 nsew signal output
rlabel metal2 s 98896 34600 98952 35000 6 dcache_mem_i_data[15]
port 458 nsew signal output
rlabel metal2 s 21840 34600 21896 35000 6 dcache_mem_i_data[1]
port 459 nsew signal output
rlabel metal2 s 29008 34600 29064 35000 6 dcache_mem_i_data[2]
port 460 nsew signal output
rlabel metal2 s 34384 34600 34440 35000 6 dcache_mem_i_data[3]
port 461 nsew signal output
rlabel metal2 s 39760 34600 39816 35000 6 dcache_mem_i_data[4]
port 462 nsew signal output
rlabel metal2 s 45136 34600 45192 35000 6 dcache_mem_i_data[5]
port 463 nsew signal output
rlabel metal2 s 50512 34600 50568 35000 6 dcache_mem_i_data[6]
port 464 nsew signal output
rlabel metal2 s 55888 34600 55944 35000 6 dcache_mem_i_data[7]
port 465 nsew signal output
rlabel metal2 s 61264 34600 61320 35000 6 dcache_mem_i_data[8]
port 466 nsew signal output
rlabel metal2 s 66640 34600 66696 35000 6 dcache_mem_i_data[9]
port 467 nsew signal output
rlabel metal2 s 15568 34600 15624 35000 6 dcache_mem_o_data[0]
port 468 nsew signal input
rlabel metal2 s 72912 34600 72968 35000 6 dcache_mem_o_data[10]
port 469 nsew signal input
rlabel metal2 s 78288 34600 78344 35000 6 dcache_mem_o_data[11]
port 470 nsew signal input
rlabel metal2 s 83664 34600 83720 35000 6 dcache_mem_o_data[12]
port 471 nsew signal input
rlabel metal2 s 89040 34600 89096 35000 6 dcache_mem_o_data[13]
port 472 nsew signal input
rlabel metal2 s 94416 34600 94472 35000 6 dcache_mem_o_data[14]
port 473 nsew signal input
rlabel metal2 s 99792 34600 99848 35000 6 dcache_mem_o_data[15]
port 474 nsew signal input
rlabel metal2 s 22736 34600 22792 35000 6 dcache_mem_o_data[1]
port 475 nsew signal input
rlabel metal2 s 29904 34600 29960 35000 6 dcache_mem_o_data[2]
port 476 nsew signal input
rlabel metal2 s 35280 34600 35336 35000 6 dcache_mem_o_data[3]
port 477 nsew signal input
rlabel metal2 s 40656 34600 40712 35000 6 dcache_mem_o_data[4]
port 478 nsew signal input
rlabel metal2 s 46032 34600 46088 35000 6 dcache_mem_o_data[5]
port 479 nsew signal input
rlabel metal2 s 51408 34600 51464 35000 6 dcache_mem_o_data[6]
port 480 nsew signal input
rlabel metal2 s 56784 34600 56840 35000 6 dcache_mem_o_data[7]
port 481 nsew signal input
rlabel metal2 s 62160 34600 62216 35000 6 dcache_mem_o_data[8]
port 482 nsew signal input
rlabel metal2 s 67536 34600 67592 35000 6 dcache_mem_o_data[9]
port 483 nsew signal input
rlabel metal2 s 5712 34600 5768 35000 6 dcache_mem_req
port 484 nsew signal output
rlabel metal2 s 16464 34600 16520 35000 6 dcache_mem_sel[0]
port 485 nsew signal output
rlabel metal2 s 23632 34600 23688 35000 6 dcache_mem_sel[1]
port 486 nsew signal output
rlabel metal2 s 6608 34600 6664 35000 6 dcache_mem_we
port 487 nsew signal output
rlabel metal2 s 7504 34600 7560 35000 6 dcache_rst
port 488 nsew signal output
rlabel metal2 s 8400 34600 8456 35000 6 dcache_wb_4_burst
port 489 nsew signal input
rlabel metal2 s 9296 34600 9352 35000 6 dcache_wb_ack
port 490 nsew signal output
rlabel metal2 s 17360 34600 17416 35000 6 dcache_wb_adr[0]
port 491 nsew signal input
rlabel metal2 s 73808 34600 73864 35000 6 dcache_wb_adr[10]
port 492 nsew signal input
rlabel metal2 s 79184 34600 79240 35000 6 dcache_wb_adr[11]
port 493 nsew signal input
rlabel metal2 s 84560 34600 84616 35000 6 dcache_wb_adr[12]
port 494 nsew signal input
rlabel metal2 s 89936 34600 89992 35000 6 dcache_wb_adr[13]
port 495 nsew signal input
rlabel metal2 s 95312 34600 95368 35000 6 dcache_wb_adr[14]
port 496 nsew signal input
rlabel metal2 s 100688 34600 100744 35000 6 dcache_wb_adr[15]
port 497 nsew signal input
rlabel metal2 s 104272 34600 104328 35000 6 dcache_wb_adr[16]
port 498 nsew signal input
rlabel metal2 s 106064 34600 106120 35000 6 dcache_wb_adr[17]
port 499 nsew signal input
rlabel metal2 s 107856 34600 107912 35000 6 dcache_wb_adr[18]
port 500 nsew signal input
rlabel metal2 s 109648 34600 109704 35000 6 dcache_wb_adr[19]
port 501 nsew signal input
rlabel metal2 s 24528 34600 24584 35000 6 dcache_wb_adr[1]
port 502 nsew signal input
rlabel metal2 s 111440 34600 111496 35000 6 dcache_wb_adr[20]
port 503 nsew signal input
rlabel metal2 s 113232 34600 113288 35000 6 dcache_wb_adr[21]
port 504 nsew signal input
rlabel metal2 s 115024 34600 115080 35000 6 dcache_wb_adr[22]
port 505 nsew signal input
rlabel metal2 s 116816 34600 116872 35000 6 dcache_wb_adr[23]
port 506 nsew signal input
rlabel metal2 s 30800 34600 30856 35000 6 dcache_wb_adr[2]
port 507 nsew signal input
rlabel metal2 s 36176 34600 36232 35000 6 dcache_wb_adr[3]
port 508 nsew signal input
rlabel metal2 s 41552 34600 41608 35000 6 dcache_wb_adr[4]
port 509 nsew signal input
rlabel metal2 s 46928 34600 46984 35000 6 dcache_wb_adr[5]
port 510 nsew signal input
rlabel metal2 s 52304 34600 52360 35000 6 dcache_wb_adr[6]
port 511 nsew signal input
rlabel metal2 s 57680 34600 57736 35000 6 dcache_wb_adr[7]
port 512 nsew signal input
rlabel metal2 s 63056 34600 63112 35000 6 dcache_wb_adr[8]
port 513 nsew signal input
rlabel metal2 s 68432 34600 68488 35000 6 dcache_wb_adr[9]
port 514 nsew signal input
rlabel metal2 s 10192 34600 10248 35000 6 dcache_wb_cyc
port 515 nsew signal input
rlabel metal2 s 11088 34600 11144 35000 6 dcache_wb_err
port 516 nsew signal output
rlabel metal2 s 18256 34600 18312 35000 6 dcache_wb_i_dat[0]
port 517 nsew signal output
rlabel metal2 s 74704 34600 74760 35000 6 dcache_wb_i_dat[10]
port 518 nsew signal output
rlabel metal2 s 80080 34600 80136 35000 6 dcache_wb_i_dat[11]
port 519 nsew signal output
rlabel metal2 s 85456 34600 85512 35000 6 dcache_wb_i_dat[12]
port 520 nsew signal output
rlabel metal2 s 90832 34600 90888 35000 6 dcache_wb_i_dat[13]
port 521 nsew signal output
rlabel metal2 s 96208 34600 96264 35000 6 dcache_wb_i_dat[14]
port 522 nsew signal output
rlabel metal2 s 101584 34600 101640 35000 6 dcache_wb_i_dat[15]
port 523 nsew signal output
rlabel metal2 s 25424 34600 25480 35000 6 dcache_wb_i_dat[1]
port 524 nsew signal output
rlabel metal2 s 31696 34600 31752 35000 6 dcache_wb_i_dat[2]
port 525 nsew signal output
rlabel metal2 s 37072 34600 37128 35000 6 dcache_wb_i_dat[3]
port 526 nsew signal output
rlabel metal2 s 42448 34600 42504 35000 6 dcache_wb_i_dat[4]
port 527 nsew signal output
rlabel metal2 s 47824 34600 47880 35000 6 dcache_wb_i_dat[5]
port 528 nsew signal output
rlabel metal2 s 53200 34600 53256 35000 6 dcache_wb_i_dat[6]
port 529 nsew signal output
rlabel metal2 s 58576 34600 58632 35000 6 dcache_wb_i_dat[7]
port 530 nsew signal output
rlabel metal2 s 63952 34600 64008 35000 6 dcache_wb_i_dat[8]
port 531 nsew signal output
rlabel metal2 s 69328 34600 69384 35000 6 dcache_wb_i_dat[9]
port 532 nsew signal output
rlabel metal2 s 19152 34600 19208 35000 6 dcache_wb_o_dat[0]
port 533 nsew signal input
rlabel metal2 s 75600 34600 75656 35000 6 dcache_wb_o_dat[10]
port 534 nsew signal input
rlabel metal2 s 80976 34600 81032 35000 6 dcache_wb_o_dat[11]
port 535 nsew signal input
rlabel metal2 s 86352 34600 86408 35000 6 dcache_wb_o_dat[12]
port 536 nsew signal input
rlabel metal2 s 91728 34600 91784 35000 6 dcache_wb_o_dat[13]
port 537 nsew signal input
rlabel metal2 s 97104 34600 97160 35000 6 dcache_wb_o_dat[14]
port 538 nsew signal input
rlabel metal2 s 102480 34600 102536 35000 6 dcache_wb_o_dat[15]
port 539 nsew signal input
rlabel metal2 s 26320 34600 26376 35000 6 dcache_wb_o_dat[1]
port 540 nsew signal input
rlabel metal2 s 32592 34600 32648 35000 6 dcache_wb_o_dat[2]
port 541 nsew signal input
rlabel metal2 s 37968 34600 38024 35000 6 dcache_wb_o_dat[3]
port 542 nsew signal input
rlabel metal2 s 43344 34600 43400 35000 6 dcache_wb_o_dat[4]
port 543 nsew signal input
rlabel metal2 s 48720 34600 48776 35000 6 dcache_wb_o_dat[5]
port 544 nsew signal input
rlabel metal2 s 54096 34600 54152 35000 6 dcache_wb_o_dat[6]
port 545 nsew signal input
rlabel metal2 s 59472 34600 59528 35000 6 dcache_wb_o_dat[7]
port 546 nsew signal input
rlabel metal2 s 64848 34600 64904 35000 6 dcache_wb_o_dat[8]
port 547 nsew signal input
rlabel metal2 s 70224 34600 70280 35000 6 dcache_wb_o_dat[9]
port 548 nsew signal input
rlabel metal2 s 20048 34600 20104 35000 6 dcache_wb_sel[0]
port 549 nsew signal input
rlabel metal2 s 27216 34600 27272 35000 6 dcache_wb_sel[1]
port 550 nsew signal input
rlabel metal2 s 11984 34600 12040 35000 6 dcache_wb_stb
port 551 nsew signal input
rlabel metal2 s 12880 34600 12936 35000 6 dcache_wb_we
port 552 nsew signal input
rlabel metal3 s 0 2128 400 2184 6 ic0_mem_ack
port 553 nsew signal input
rlabel metal3 s 0 5488 400 5544 6 ic0_mem_addr[0]
port 554 nsew signal output
rlabel metal3 s 0 19600 400 19656 6 ic0_mem_addr[10]
port 555 nsew signal output
rlabel metal3 s 0 20944 400 21000 6 ic0_mem_addr[11]
port 556 nsew signal output
rlabel metal3 s 0 22288 400 22344 6 ic0_mem_addr[12]
port 557 nsew signal output
rlabel metal3 s 0 23632 400 23688 6 ic0_mem_addr[13]
port 558 nsew signal output
rlabel metal3 s 0 24976 400 25032 6 ic0_mem_addr[14]
port 559 nsew signal output
rlabel metal3 s 0 26320 400 26376 6 ic0_mem_addr[15]
port 560 nsew signal output
rlabel metal3 s 0 7168 400 7224 6 ic0_mem_addr[1]
port 561 nsew signal output
rlabel metal3 s 0 8848 400 8904 6 ic0_mem_addr[2]
port 562 nsew signal output
rlabel metal3 s 0 10192 400 10248 6 ic0_mem_addr[3]
port 563 nsew signal output
rlabel metal3 s 0 11536 400 11592 6 ic0_mem_addr[4]
port 564 nsew signal output
rlabel metal3 s 0 12880 400 12936 6 ic0_mem_addr[5]
port 565 nsew signal output
rlabel metal3 s 0 14224 400 14280 6 ic0_mem_addr[6]
port 566 nsew signal output
rlabel metal3 s 0 15568 400 15624 6 ic0_mem_addr[7]
port 567 nsew signal output
rlabel metal3 s 0 16912 400 16968 6 ic0_mem_addr[8]
port 568 nsew signal output
rlabel metal3 s 0 18256 400 18312 6 ic0_mem_addr[9]
port 569 nsew signal output
rlabel metal3 s 0 2464 400 2520 6 ic0_mem_cache_flush
port 570 nsew signal output
rlabel metal3 s 0 5824 400 5880 6 ic0_mem_data[0]
port 571 nsew signal input
rlabel metal3 s 0 19936 400 19992 6 ic0_mem_data[10]
port 572 nsew signal input
rlabel metal3 s 0 21280 400 21336 6 ic0_mem_data[11]
port 573 nsew signal input
rlabel metal3 s 0 22624 400 22680 6 ic0_mem_data[12]
port 574 nsew signal input
rlabel metal3 s 0 23968 400 24024 6 ic0_mem_data[13]
port 575 nsew signal input
rlabel metal3 s 0 25312 400 25368 6 ic0_mem_data[14]
port 576 nsew signal input
rlabel metal3 s 0 26656 400 26712 6 ic0_mem_data[15]
port 577 nsew signal input
rlabel metal3 s 0 27664 400 27720 6 ic0_mem_data[16]
port 578 nsew signal input
rlabel metal3 s 0 28000 400 28056 6 ic0_mem_data[17]
port 579 nsew signal input
rlabel metal3 s 0 28336 400 28392 6 ic0_mem_data[18]
port 580 nsew signal input
rlabel metal3 s 0 28672 400 28728 6 ic0_mem_data[19]
port 581 nsew signal input
rlabel metal3 s 0 7504 400 7560 6 ic0_mem_data[1]
port 582 nsew signal input
rlabel metal3 s 0 29008 400 29064 6 ic0_mem_data[20]
port 583 nsew signal input
rlabel metal3 s 0 29344 400 29400 6 ic0_mem_data[21]
port 584 nsew signal input
rlabel metal3 s 0 29680 400 29736 6 ic0_mem_data[22]
port 585 nsew signal input
rlabel metal3 s 0 30016 400 30072 6 ic0_mem_data[23]
port 586 nsew signal input
rlabel metal3 s 0 30352 400 30408 6 ic0_mem_data[24]
port 587 nsew signal input
rlabel metal3 s 0 30688 400 30744 6 ic0_mem_data[25]
port 588 nsew signal input
rlabel metal3 s 0 31024 400 31080 6 ic0_mem_data[26]
port 589 nsew signal input
rlabel metal3 s 0 31360 400 31416 6 ic0_mem_data[27]
port 590 nsew signal input
rlabel metal3 s 0 31696 400 31752 6 ic0_mem_data[28]
port 591 nsew signal input
rlabel metal3 s 0 32032 400 32088 6 ic0_mem_data[29]
port 592 nsew signal input
rlabel metal3 s 0 9184 400 9240 6 ic0_mem_data[2]
port 593 nsew signal input
rlabel metal3 s 0 32368 400 32424 6 ic0_mem_data[30]
port 594 nsew signal input
rlabel metal3 s 0 32704 400 32760 6 ic0_mem_data[31]
port 595 nsew signal input
rlabel metal3 s 0 10528 400 10584 6 ic0_mem_data[3]
port 596 nsew signal input
rlabel metal3 s 0 11872 400 11928 6 ic0_mem_data[4]
port 597 nsew signal input
rlabel metal3 s 0 13216 400 13272 6 ic0_mem_data[5]
port 598 nsew signal input
rlabel metal3 s 0 14560 400 14616 6 ic0_mem_data[6]
port 599 nsew signal input
rlabel metal3 s 0 15904 400 15960 6 ic0_mem_data[7]
port 600 nsew signal input
rlabel metal3 s 0 17248 400 17304 6 ic0_mem_data[8]
port 601 nsew signal input
rlabel metal3 s 0 18592 400 18648 6 ic0_mem_data[9]
port 602 nsew signal input
rlabel metal3 s 0 2800 400 2856 6 ic0_mem_ppl_submit
port 603 nsew signal output
rlabel metal3 s 0 3136 400 3192 6 ic0_mem_req
port 604 nsew signal output
rlabel metal3 s 0 3472 400 3528 6 ic0_rst
port 605 nsew signal output
rlabel metal3 s 0 3808 400 3864 6 ic0_wb_ack
port 606 nsew signal output
rlabel metal3 s 0 6160 400 6216 6 ic0_wb_adr[0]
port 607 nsew signal input
rlabel metal3 s 0 20272 400 20328 6 ic0_wb_adr[10]
port 608 nsew signal input
rlabel metal3 s 0 21616 400 21672 6 ic0_wb_adr[11]
port 609 nsew signal input
rlabel metal3 s 0 22960 400 23016 6 ic0_wb_adr[12]
port 610 nsew signal input
rlabel metal3 s 0 24304 400 24360 6 ic0_wb_adr[13]
port 611 nsew signal input
rlabel metal3 s 0 25648 400 25704 6 ic0_wb_adr[14]
port 612 nsew signal input
rlabel metal3 s 0 26992 400 27048 6 ic0_wb_adr[15]
port 613 nsew signal input
rlabel metal3 s 0 7840 400 7896 6 ic0_wb_adr[1]
port 614 nsew signal input
rlabel metal3 s 0 9520 400 9576 6 ic0_wb_adr[2]
port 615 nsew signal input
rlabel metal3 s 0 10864 400 10920 6 ic0_wb_adr[3]
port 616 nsew signal input
rlabel metal3 s 0 12208 400 12264 6 ic0_wb_adr[4]
port 617 nsew signal input
rlabel metal3 s 0 13552 400 13608 6 ic0_wb_adr[5]
port 618 nsew signal input
rlabel metal3 s 0 14896 400 14952 6 ic0_wb_adr[6]
port 619 nsew signal input
rlabel metal3 s 0 16240 400 16296 6 ic0_wb_adr[7]
port 620 nsew signal input
rlabel metal3 s 0 17584 400 17640 6 ic0_wb_adr[8]
port 621 nsew signal input
rlabel metal3 s 0 18928 400 18984 6 ic0_wb_adr[9]
port 622 nsew signal input
rlabel metal3 s 0 4144 400 4200 6 ic0_wb_cyc
port 623 nsew signal input
rlabel metal3 s 0 4480 400 4536 6 ic0_wb_err
port 624 nsew signal output
rlabel metal3 s 0 6496 400 6552 6 ic0_wb_i_dat[0]
port 625 nsew signal output
rlabel metal3 s 0 20608 400 20664 6 ic0_wb_i_dat[10]
port 626 nsew signal output
rlabel metal3 s 0 21952 400 22008 6 ic0_wb_i_dat[11]
port 627 nsew signal output
rlabel metal3 s 0 23296 400 23352 6 ic0_wb_i_dat[12]
port 628 nsew signal output
rlabel metal3 s 0 24640 400 24696 6 ic0_wb_i_dat[13]
port 629 nsew signal output
rlabel metal3 s 0 25984 400 26040 6 ic0_wb_i_dat[14]
port 630 nsew signal output
rlabel metal3 s 0 27328 400 27384 6 ic0_wb_i_dat[15]
port 631 nsew signal output
rlabel metal3 s 0 8176 400 8232 6 ic0_wb_i_dat[1]
port 632 nsew signal output
rlabel metal3 s 0 9856 400 9912 6 ic0_wb_i_dat[2]
port 633 nsew signal output
rlabel metal3 s 0 11200 400 11256 6 ic0_wb_i_dat[3]
port 634 nsew signal output
rlabel metal3 s 0 12544 400 12600 6 ic0_wb_i_dat[4]
port 635 nsew signal output
rlabel metal3 s 0 13888 400 13944 6 ic0_wb_i_dat[5]
port 636 nsew signal output
rlabel metal3 s 0 15232 400 15288 6 ic0_wb_i_dat[6]
port 637 nsew signal output
rlabel metal3 s 0 16576 400 16632 6 ic0_wb_i_dat[7]
port 638 nsew signal output
rlabel metal3 s 0 17920 400 17976 6 ic0_wb_i_dat[8]
port 639 nsew signal output
rlabel metal3 s 0 19264 400 19320 6 ic0_wb_i_dat[9]
port 640 nsew signal output
rlabel metal3 s 0 6832 400 6888 6 ic0_wb_sel[0]
port 641 nsew signal input
rlabel metal3 s 0 8512 400 8568 6 ic0_wb_sel[1]
port 642 nsew signal input
rlabel metal3 s 0 4816 400 4872 6 ic0_wb_stb
port 643 nsew signal input
rlabel metal3 s 0 5152 400 5208 6 ic0_wb_we
port 644 nsew signal input
rlabel metal3 s 119600 2128 120000 2184 6 ic1_mem_ack
port 645 nsew signal input
rlabel metal3 s 119600 5488 120000 5544 6 ic1_mem_addr[0]
port 646 nsew signal output
rlabel metal3 s 119600 19600 120000 19656 6 ic1_mem_addr[10]
port 647 nsew signal output
rlabel metal3 s 119600 20944 120000 21000 6 ic1_mem_addr[11]
port 648 nsew signal output
rlabel metal3 s 119600 22288 120000 22344 6 ic1_mem_addr[12]
port 649 nsew signal output
rlabel metal3 s 119600 23632 120000 23688 6 ic1_mem_addr[13]
port 650 nsew signal output
rlabel metal3 s 119600 24976 120000 25032 6 ic1_mem_addr[14]
port 651 nsew signal output
rlabel metal3 s 119600 26320 120000 26376 6 ic1_mem_addr[15]
port 652 nsew signal output
rlabel metal3 s 119600 7168 120000 7224 6 ic1_mem_addr[1]
port 653 nsew signal output
rlabel metal3 s 119600 8848 120000 8904 6 ic1_mem_addr[2]
port 654 nsew signal output
rlabel metal3 s 119600 10192 120000 10248 6 ic1_mem_addr[3]
port 655 nsew signal output
rlabel metal3 s 119600 11536 120000 11592 6 ic1_mem_addr[4]
port 656 nsew signal output
rlabel metal3 s 119600 12880 120000 12936 6 ic1_mem_addr[5]
port 657 nsew signal output
rlabel metal3 s 119600 14224 120000 14280 6 ic1_mem_addr[6]
port 658 nsew signal output
rlabel metal3 s 119600 15568 120000 15624 6 ic1_mem_addr[7]
port 659 nsew signal output
rlabel metal3 s 119600 16912 120000 16968 6 ic1_mem_addr[8]
port 660 nsew signal output
rlabel metal3 s 119600 18256 120000 18312 6 ic1_mem_addr[9]
port 661 nsew signal output
rlabel metal3 s 119600 2464 120000 2520 6 ic1_mem_cache_flush
port 662 nsew signal output
rlabel metal3 s 119600 5824 120000 5880 6 ic1_mem_data[0]
port 663 nsew signal input
rlabel metal3 s 119600 19936 120000 19992 6 ic1_mem_data[10]
port 664 nsew signal input
rlabel metal3 s 119600 21280 120000 21336 6 ic1_mem_data[11]
port 665 nsew signal input
rlabel metal3 s 119600 22624 120000 22680 6 ic1_mem_data[12]
port 666 nsew signal input
rlabel metal3 s 119600 23968 120000 24024 6 ic1_mem_data[13]
port 667 nsew signal input
rlabel metal3 s 119600 25312 120000 25368 6 ic1_mem_data[14]
port 668 nsew signal input
rlabel metal3 s 119600 26656 120000 26712 6 ic1_mem_data[15]
port 669 nsew signal input
rlabel metal3 s 119600 27664 120000 27720 6 ic1_mem_data[16]
port 670 nsew signal input
rlabel metal3 s 119600 28000 120000 28056 6 ic1_mem_data[17]
port 671 nsew signal input
rlabel metal3 s 119600 28336 120000 28392 6 ic1_mem_data[18]
port 672 nsew signal input
rlabel metal3 s 119600 28672 120000 28728 6 ic1_mem_data[19]
port 673 nsew signal input
rlabel metal3 s 119600 7504 120000 7560 6 ic1_mem_data[1]
port 674 nsew signal input
rlabel metal3 s 119600 29008 120000 29064 6 ic1_mem_data[20]
port 675 nsew signal input
rlabel metal3 s 119600 29344 120000 29400 6 ic1_mem_data[21]
port 676 nsew signal input
rlabel metal3 s 119600 29680 120000 29736 6 ic1_mem_data[22]
port 677 nsew signal input
rlabel metal3 s 119600 30016 120000 30072 6 ic1_mem_data[23]
port 678 nsew signal input
rlabel metal3 s 119600 30352 120000 30408 6 ic1_mem_data[24]
port 679 nsew signal input
rlabel metal3 s 119600 30688 120000 30744 6 ic1_mem_data[25]
port 680 nsew signal input
rlabel metal3 s 119600 31024 120000 31080 6 ic1_mem_data[26]
port 681 nsew signal input
rlabel metal3 s 119600 31360 120000 31416 6 ic1_mem_data[27]
port 682 nsew signal input
rlabel metal3 s 119600 31696 120000 31752 6 ic1_mem_data[28]
port 683 nsew signal input
rlabel metal3 s 119600 32032 120000 32088 6 ic1_mem_data[29]
port 684 nsew signal input
rlabel metal3 s 119600 9184 120000 9240 6 ic1_mem_data[2]
port 685 nsew signal input
rlabel metal3 s 119600 32368 120000 32424 6 ic1_mem_data[30]
port 686 nsew signal input
rlabel metal3 s 119600 32704 120000 32760 6 ic1_mem_data[31]
port 687 nsew signal input
rlabel metal3 s 119600 10528 120000 10584 6 ic1_mem_data[3]
port 688 nsew signal input
rlabel metal3 s 119600 11872 120000 11928 6 ic1_mem_data[4]
port 689 nsew signal input
rlabel metal3 s 119600 13216 120000 13272 6 ic1_mem_data[5]
port 690 nsew signal input
rlabel metal3 s 119600 14560 120000 14616 6 ic1_mem_data[6]
port 691 nsew signal input
rlabel metal3 s 119600 15904 120000 15960 6 ic1_mem_data[7]
port 692 nsew signal input
rlabel metal3 s 119600 17248 120000 17304 6 ic1_mem_data[8]
port 693 nsew signal input
rlabel metal3 s 119600 18592 120000 18648 6 ic1_mem_data[9]
port 694 nsew signal input
rlabel metal3 s 119600 2800 120000 2856 6 ic1_mem_ppl_submit
port 695 nsew signal output
rlabel metal3 s 119600 3136 120000 3192 6 ic1_mem_req
port 696 nsew signal output
rlabel metal3 s 119600 3472 120000 3528 6 ic1_rst
port 697 nsew signal output
rlabel metal3 s 119600 3808 120000 3864 6 ic1_wb_ack
port 698 nsew signal output
rlabel metal3 s 119600 6160 120000 6216 6 ic1_wb_adr[0]
port 699 nsew signal input
rlabel metal3 s 119600 20272 120000 20328 6 ic1_wb_adr[10]
port 700 nsew signal input
rlabel metal3 s 119600 21616 120000 21672 6 ic1_wb_adr[11]
port 701 nsew signal input
rlabel metal3 s 119600 22960 120000 23016 6 ic1_wb_adr[12]
port 702 nsew signal input
rlabel metal3 s 119600 24304 120000 24360 6 ic1_wb_adr[13]
port 703 nsew signal input
rlabel metal3 s 119600 25648 120000 25704 6 ic1_wb_adr[14]
port 704 nsew signal input
rlabel metal3 s 119600 26992 120000 27048 6 ic1_wb_adr[15]
port 705 nsew signal input
rlabel metal3 s 119600 7840 120000 7896 6 ic1_wb_adr[1]
port 706 nsew signal input
rlabel metal3 s 119600 9520 120000 9576 6 ic1_wb_adr[2]
port 707 nsew signal input
rlabel metal3 s 119600 10864 120000 10920 6 ic1_wb_adr[3]
port 708 nsew signal input
rlabel metal3 s 119600 12208 120000 12264 6 ic1_wb_adr[4]
port 709 nsew signal input
rlabel metal3 s 119600 13552 120000 13608 6 ic1_wb_adr[5]
port 710 nsew signal input
rlabel metal3 s 119600 14896 120000 14952 6 ic1_wb_adr[6]
port 711 nsew signal input
rlabel metal3 s 119600 16240 120000 16296 6 ic1_wb_adr[7]
port 712 nsew signal input
rlabel metal3 s 119600 17584 120000 17640 6 ic1_wb_adr[8]
port 713 nsew signal input
rlabel metal3 s 119600 18928 120000 18984 6 ic1_wb_adr[9]
port 714 nsew signal input
rlabel metal3 s 119600 4144 120000 4200 6 ic1_wb_cyc
port 715 nsew signal input
rlabel metal3 s 119600 4480 120000 4536 6 ic1_wb_err
port 716 nsew signal output
rlabel metal3 s 119600 6496 120000 6552 6 ic1_wb_i_dat[0]
port 717 nsew signal output
rlabel metal3 s 119600 20608 120000 20664 6 ic1_wb_i_dat[10]
port 718 nsew signal output
rlabel metal3 s 119600 21952 120000 22008 6 ic1_wb_i_dat[11]
port 719 nsew signal output
rlabel metal3 s 119600 23296 120000 23352 6 ic1_wb_i_dat[12]
port 720 nsew signal output
rlabel metal3 s 119600 24640 120000 24696 6 ic1_wb_i_dat[13]
port 721 nsew signal output
rlabel metal3 s 119600 25984 120000 26040 6 ic1_wb_i_dat[14]
port 722 nsew signal output
rlabel metal3 s 119600 27328 120000 27384 6 ic1_wb_i_dat[15]
port 723 nsew signal output
rlabel metal3 s 119600 8176 120000 8232 6 ic1_wb_i_dat[1]
port 724 nsew signal output
rlabel metal3 s 119600 9856 120000 9912 6 ic1_wb_i_dat[2]
port 725 nsew signal output
rlabel metal3 s 119600 11200 120000 11256 6 ic1_wb_i_dat[3]
port 726 nsew signal output
rlabel metal3 s 119600 12544 120000 12600 6 ic1_wb_i_dat[4]
port 727 nsew signal output
rlabel metal3 s 119600 13888 120000 13944 6 ic1_wb_i_dat[5]
port 728 nsew signal output
rlabel metal3 s 119600 15232 120000 15288 6 ic1_wb_i_dat[6]
port 729 nsew signal output
rlabel metal3 s 119600 16576 120000 16632 6 ic1_wb_i_dat[7]
port 730 nsew signal output
rlabel metal3 s 119600 17920 120000 17976 6 ic1_wb_i_dat[8]
port 731 nsew signal output
rlabel metal3 s 119600 19264 120000 19320 6 ic1_wb_i_dat[9]
port 732 nsew signal output
rlabel metal3 s 119600 6832 120000 6888 6 ic1_wb_sel[0]
port 733 nsew signal input
rlabel metal3 s 119600 8512 120000 8568 6 ic1_wb_sel[1]
port 734 nsew signal input
rlabel metal3 s 119600 4816 120000 4872 6 ic1_wb_stb
port 735 nsew signal input
rlabel metal3 s 119600 5152 120000 5208 6 ic1_wb_we
port 736 nsew signal input
rlabel metal2 s 52640 0 52696 400 6 inner_disable
port 737 nsew signal input
rlabel metal2 s 52864 0 52920 400 6 inner_embed_mode
port 738 nsew signal input
rlabel metal2 s 53088 0 53144 400 6 inner_ext_irq
port 739 nsew signal input
rlabel metal2 s 53312 0 53368 400 6 inner_wb_4_burst
port 740 nsew signal output
rlabel metal2 s 53536 0 53592 400 6 inner_wb_8_burst
port 741 nsew signal output
rlabel metal2 s 53760 0 53816 400 6 inner_wb_ack
port 742 nsew signal input
rlabel metal2 s 54880 0 54936 400 6 inner_wb_adr[0]
port 743 nsew signal output
rlabel metal2 s 62048 0 62104 400 6 inner_wb_adr[10]
port 744 nsew signal output
rlabel metal2 s 62720 0 62776 400 6 inner_wb_adr[11]
port 745 nsew signal output
rlabel metal2 s 63392 0 63448 400 6 inner_wb_adr[12]
port 746 nsew signal output
rlabel metal2 s 64064 0 64120 400 6 inner_wb_adr[13]
port 747 nsew signal output
rlabel metal2 s 64736 0 64792 400 6 inner_wb_adr[14]
port 748 nsew signal output
rlabel metal2 s 65408 0 65464 400 6 inner_wb_adr[15]
port 749 nsew signal output
rlabel metal2 s 66080 0 66136 400 6 inner_wb_adr[16]
port 750 nsew signal output
rlabel metal2 s 66304 0 66360 400 6 inner_wb_adr[17]
port 751 nsew signal output
rlabel metal2 s 66528 0 66584 400 6 inner_wb_adr[18]
port 752 nsew signal output
rlabel metal2 s 66752 0 66808 400 6 inner_wb_adr[19]
port 753 nsew signal output
rlabel metal2 s 55776 0 55832 400 6 inner_wb_adr[1]
port 754 nsew signal output
rlabel metal2 s 66976 0 67032 400 6 inner_wb_adr[20]
port 755 nsew signal output
rlabel metal2 s 67200 0 67256 400 6 inner_wb_adr[21]
port 756 nsew signal output
rlabel metal2 s 67424 0 67480 400 6 inner_wb_adr[22]
port 757 nsew signal output
rlabel metal2 s 67648 0 67704 400 6 inner_wb_adr[23]
port 758 nsew signal output
rlabel metal2 s 56672 0 56728 400 6 inner_wb_adr[2]
port 759 nsew signal output
rlabel metal2 s 57344 0 57400 400 6 inner_wb_adr[3]
port 760 nsew signal output
rlabel metal2 s 58016 0 58072 400 6 inner_wb_adr[4]
port 761 nsew signal output
rlabel metal2 s 58688 0 58744 400 6 inner_wb_adr[5]
port 762 nsew signal output
rlabel metal2 s 59360 0 59416 400 6 inner_wb_adr[6]
port 763 nsew signal output
rlabel metal2 s 60032 0 60088 400 6 inner_wb_adr[7]
port 764 nsew signal output
rlabel metal2 s 60704 0 60760 400 6 inner_wb_adr[8]
port 765 nsew signal output
rlabel metal2 s 61376 0 61432 400 6 inner_wb_adr[9]
port 766 nsew signal output
rlabel metal2 s 53984 0 54040 400 6 inner_wb_cyc
port 767 nsew signal output
rlabel metal2 s 54208 0 54264 400 6 inner_wb_err
port 768 nsew signal input
rlabel metal2 s 55104 0 55160 400 6 inner_wb_i_dat[0]
port 769 nsew signal input
rlabel metal2 s 62272 0 62328 400 6 inner_wb_i_dat[10]
port 770 nsew signal input
rlabel metal2 s 62944 0 63000 400 6 inner_wb_i_dat[11]
port 771 nsew signal input
rlabel metal2 s 63616 0 63672 400 6 inner_wb_i_dat[12]
port 772 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 inner_wb_i_dat[13]
port 773 nsew signal input
rlabel metal2 s 64960 0 65016 400 6 inner_wb_i_dat[14]
port 774 nsew signal input
rlabel metal2 s 65632 0 65688 400 6 inner_wb_i_dat[15]
port 775 nsew signal input
rlabel metal2 s 56000 0 56056 400 6 inner_wb_i_dat[1]
port 776 nsew signal input
rlabel metal2 s 56896 0 56952 400 6 inner_wb_i_dat[2]
port 777 nsew signal input
rlabel metal2 s 57568 0 57624 400 6 inner_wb_i_dat[3]
port 778 nsew signal input
rlabel metal2 s 58240 0 58296 400 6 inner_wb_i_dat[4]
port 779 nsew signal input
rlabel metal2 s 58912 0 58968 400 6 inner_wb_i_dat[5]
port 780 nsew signal input
rlabel metal2 s 59584 0 59640 400 6 inner_wb_i_dat[6]
port 781 nsew signal input
rlabel metal2 s 60256 0 60312 400 6 inner_wb_i_dat[7]
port 782 nsew signal input
rlabel metal2 s 60928 0 60984 400 6 inner_wb_i_dat[8]
port 783 nsew signal input
rlabel metal2 s 61600 0 61656 400 6 inner_wb_i_dat[9]
port 784 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 inner_wb_o_dat[0]
port 785 nsew signal output
rlabel metal2 s 62496 0 62552 400 6 inner_wb_o_dat[10]
port 786 nsew signal output
rlabel metal2 s 63168 0 63224 400 6 inner_wb_o_dat[11]
port 787 nsew signal output
rlabel metal2 s 63840 0 63896 400 6 inner_wb_o_dat[12]
port 788 nsew signal output
rlabel metal2 s 64512 0 64568 400 6 inner_wb_o_dat[13]
port 789 nsew signal output
rlabel metal2 s 65184 0 65240 400 6 inner_wb_o_dat[14]
port 790 nsew signal output
rlabel metal2 s 65856 0 65912 400 6 inner_wb_o_dat[15]
port 791 nsew signal output
rlabel metal2 s 56224 0 56280 400 6 inner_wb_o_dat[1]
port 792 nsew signal output
rlabel metal2 s 57120 0 57176 400 6 inner_wb_o_dat[2]
port 793 nsew signal output
rlabel metal2 s 57792 0 57848 400 6 inner_wb_o_dat[3]
port 794 nsew signal output
rlabel metal2 s 58464 0 58520 400 6 inner_wb_o_dat[4]
port 795 nsew signal output
rlabel metal2 s 59136 0 59192 400 6 inner_wb_o_dat[5]
port 796 nsew signal output
rlabel metal2 s 59808 0 59864 400 6 inner_wb_o_dat[6]
port 797 nsew signal output
rlabel metal2 s 60480 0 60536 400 6 inner_wb_o_dat[7]
port 798 nsew signal output
rlabel metal2 s 61152 0 61208 400 6 inner_wb_o_dat[8]
port 799 nsew signal output
rlabel metal2 s 61824 0 61880 400 6 inner_wb_o_dat[9]
port 800 nsew signal output
rlabel metal2 s 55552 0 55608 400 6 inner_wb_sel[0]
port 801 nsew signal output
rlabel metal2 s 56448 0 56504 400 6 inner_wb_sel[1]
port 802 nsew signal output
rlabel metal2 s 54432 0 54488 400 6 inner_wb_stb
port 803 nsew signal output
rlabel metal2 s 54656 0 54712 400 6 inner_wb_we
port 804 nsew signal output
rlabel metal4 s 2224 1538 2384 33350 6 vccd1
port 805 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 33350 6 vccd1
port 805 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 33350 6 vccd1
port 805 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 33350 6 vccd1
port 805 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 33350 6 vccd1
port 805 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 33350 6 vccd1
port 805 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 33350 6 vccd1
port 805 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 33350 6 vccd1
port 805 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 33350 6 vssd1
port 806 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 33350 6 vssd1
port 806 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 33350 6 vssd1
port 806 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 33350 6 vssd1
port 806 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 33350 6 vssd1
port 806 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 33350 6 vssd1
port 806 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 33350 6 vssd1
port 806 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 33350 6 vssd1
port 806 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 120000 35000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12442090
string GDS_FILE /home/piotro/caravel_user_project/openlane/inner_interconnect/runs/23_11_07_19_07/results/signoff/interconnect_inner.magic.gds
string GDS_START 486390
<< end >>

